VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ycell
  CLASS BLOCK ;
  FOREIGN ycell ;
  ORIGIN 0.000 0.000 ;
  SIZE 65.480 BY 76.200 ;
  PIN cbitin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 72.200 17.850 76.200 ;
    END
  END cbitin
  PIN cbitout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END cbitout
  PIN confclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 72.200 10.490 76.200 ;
    END
  END confclk
  PIN confclko
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END confclko
  PIN dempty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END dempty
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END din[1]
  PIN dout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END dout[1]
  PIN hempty
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END hempty
  PIN hempty2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.480 44.240 65.480 44.840 ;
    END
  END hempty2
  PIN lempty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END lempty
  PIN lin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END lin[0]
  PIN lin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END lin[1]
  PIN lout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END lout[0]
  PIN lout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END lout[1]
  PIN rempty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.480 31.320 65.480 31.920 ;
    END
  END rempty
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 72.200 3.590 76.200 ;
    END
  END reset
  PIN reseto
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END reseto
  PIN rin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.480 18.400 65.480 19.000 ;
    END
  END rin[0]
  PIN rin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.480 6.160 65.480 6.760 ;
    END
  END rin[1]
  PIN rout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.480 69.400 65.480 70.000 ;
    END
  END rout[0]
  PIN rout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.480 56.480 65.480 57.080 ;
    END
  END rout[1]
  PIN uempty
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 72.200 39.470 76.200 ;
    END
  END uempty
  PIN uin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 72.200 32.570 76.200 ;
    END
  END uin[0]
  PIN uin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 72.200 25.210 76.200 ;
    END
  END uin[1]
  PIN uout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 72.200 61.550 76.200 ;
    END
  END uout[0]
  PIN uout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 72.200 54.190 76.200 ;
    END
  END uout[1]
  PIN vempty
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 72.200 46.830 76.200 ;
    END
  END vempty
  PIN vempty2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END vempty2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 49.955 10.640 51.555 65.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.860 10.640 33.460 65.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 13.765 10.640 15.365 65.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 40.905 10.640 42.505 65.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 22.815 10.640 24.415 65.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 59.800 65.365 ;
      LAYER met1 ;
        RECT 3.290 10.640 61.570 65.520 ;
      LAYER met2 ;
        RECT 3.870 71.920 9.930 72.200 ;
        RECT 10.770 71.920 17.290 72.200 ;
        RECT 18.130 71.920 24.650 72.200 ;
        RECT 25.490 71.920 32.010 72.200 ;
        RECT 32.850 71.920 38.910 72.200 ;
        RECT 39.750 71.920 46.270 72.200 ;
        RECT 47.110 71.920 53.630 72.200 ;
        RECT 54.470 71.920 60.990 72.200 ;
        RECT 3.320 4.280 61.540 71.920 ;
        RECT 3.870 4.000 9.930 4.280 ;
        RECT 10.770 4.000 17.290 4.280 ;
        RECT 18.130 4.000 24.650 4.280 ;
        RECT 25.490 4.000 32.010 4.280 ;
        RECT 32.850 4.000 38.910 4.280 ;
        RECT 39.750 4.000 46.270 4.280 ;
        RECT 47.110 4.000 53.630 4.280 ;
        RECT 54.470 4.000 60.990 4.280 ;
      LAYER met3 ;
        RECT 4.400 69.000 61.080 69.865 ;
        RECT 4.000 57.480 61.480 69.000 ;
        RECT 4.400 56.080 61.080 57.480 ;
        RECT 4.000 45.240 61.480 56.080 ;
        RECT 4.400 43.840 61.080 45.240 ;
        RECT 4.000 32.320 61.480 43.840 ;
        RECT 4.400 30.920 61.080 32.320 ;
        RECT 4.000 19.400 61.480 30.920 ;
        RECT 4.400 18.000 61.080 19.400 ;
        RECT 4.000 7.160 61.480 18.000 ;
        RECT 4.400 6.295 61.080 7.160 ;
      LAYER met4 ;
        RECT 24.815 10.640 31.460 65.520 ;
        RECT 33.860 10.640 40.505 65.520 ;
        RECT 42.905 10.640 49.555 65.520 ;
  END
END ycell
END LIBRARY

