*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 D Q RESET_B CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A Y VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE Z VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 D Q SET_B CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt gpio_control_block mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out pad_gpio_ana_en
+ pad_gpio_ana_pol pad_gpio_ana_sel pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover
+ pad_gpio_ib_mode_sel pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel
+ pad_gpio_vtrip_sel resetn serial_clock serial_data_in serial_data_out user_gpio_in
+ user_gpio_oeb user_gpio_out VPWR VGND
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_062_ _062_/A _062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_045_ _042_/A _045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_044_ _042_/A _044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_061_ _062_/A _061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ _062_/A _060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_043_ _042_/A _043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_042_ _042_/A _042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_041_ _081_/A _042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_040_ _064_/A _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _086_/D _087_/D _049_/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ _083_/D _086_/D _050_/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_097_ _088_/D _083_/D _051_/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_096_ _095_/Q _088_/D _053_/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_079_ _039_/A _079_/B _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__and2_4
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_095_ serial_data_in _095_/Q _054_/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_078_ resetn _079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__inv_2
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_094_ _103_/D pad_gpio_ana_pol _055_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_077_ _077_/A pad_gpio_in _077_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__nand2_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_093_ _093_/D pad_gpio_ana_sel _056_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_076_ _082_/Q _074_/X _075_/Y _077_/A user_gpio_out pad_gpio_out VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_059_ _062_/A _059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgpio_in_buf _077_/Y gpio_in_buf/TE user_gpio_in VGND VGND VPWR VPWR sky130_fd_sc_hd__einvp_8
X_092_ _100_/Q pad_gpio_ana_en _057_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ _081_/A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_075_ pad_gpio_dm[0] _073_/X _075_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__nand2_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_091_ serial_data_out pad_gpio_dm[2] _059_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_074_ mgmt_gpio_out _073_/X _074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_4
X_057_ _053_/A _057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ _106_/Q pad_gpio_dm[1] _060_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_073_ mgmt_gpio_oeb _072_/Y pad_gpio_dm[1] _073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__and3_4
X_056_ _053_/A _056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_039_ _039_/A resetn _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_072_ pad_gpio_dm[2] _072_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_1
X_055_ _053_/A _055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_107_ _106_/Q serial_data_out _081_/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_071_ _088_/Q mgmt_gpio_oeb _082_/Q user_gpio_oeb _077_/A pad_gpio_outenb VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__a32o_4
X_106_ _105_/Q _106_/Q _042_/A _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
X_054_ _053_/A _054_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_070_ _082_/Q _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__inv_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_053_ _053_/A _053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ _105_/D _105_/Q _042_/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_104_ _103_/Q _105_/D _043_/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
X_052_ _081_/A _053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_051_ _051_/A _051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_103_ _103_/D _103_/Q _044_/X _039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_050_ _051_/A _050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_102_ _093_/D _103_/D _045_/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgpio_logic_high gpio_in_buf/TE gpio_logic_high/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_101_ _100_/Q _093_/D _047_/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ _087_/D _100_/Q _048_/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ _105_/Q pad_gpio_dm[0] _061_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfstp_4
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X _097_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_serial_clock serial_clock clkbuf_0_serial_clock/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_088_ _088_/D _088_/Q _062_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_087_ _087_/D pad_gpio_ib_mode_sel _063_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_086_ _086_/D pad_gpio_inenb _065_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ _069_/A _069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_085_ _105_/D pad_gpio_vtrip_sel _066_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_068_ _069_/A _068_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_067_ _069_/A _067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_084_ _103_/Q pad_gpio_slow_sel _067_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 serial_data_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ _083_/D pad_gpio_holdover _068_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfrtp_4
X_066_ _069_/A _066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_049_ _051_/A _049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_065_ _069_/A _065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_082_ _095_/Q _082_/Q _069_/X _079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_048_ _051_/A _048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_081_ _081_/A _081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_064_ _064_/A _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_047_ _051_/A _047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_080_ _082_/Q pad_gpio_in mgmt_gpio_in VGND VGND VPWR VPWR sky130_fd_sc_hd__and2_4
X_063_ _062_/A _063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_046_ _081_/A _051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

