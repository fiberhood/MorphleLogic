// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module mgmt_protect_hv(mprj2_vdd_logic1, mprj_vdd_logic1, vccd, vssd, vdda1, vssa1, vdda2, vssa2);
  output mprj2_vdd_logic1;
  wire mprj2_vdd_logic1_h;
  output mprj_vdd_logic1;
  wire mprj_vdd_logic1_h;
  input vccd;
  input vdda1;
  input vdda2;
  input vssa1;
  input vssa2;
  input vssd;
  sky130_fd_sc_hvl__decap_8 FILLER_0_0 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_136 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_152 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_16 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_168 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_176 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_216 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_232 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_24 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_240 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_248 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_256 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_264 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_272 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_4 FILLER_0_296 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_0_300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_64 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_72 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_8 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_88 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_96 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_0 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_4 FILLER_1_131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_148 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_156 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_16 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_164 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_172 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_188 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_220 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_24 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_244 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_252 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_260 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_268 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_4 FILLER_1_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_1_280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_1_282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_1_300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_1_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_4 FILLER_1_78 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_8 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_99 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_0 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_139 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_155 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_16 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_163 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_179 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_187 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_195 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_203 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_211 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_219 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_235 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_24 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_251 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_259 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_2_300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_64 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_72 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_8 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_2_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_99 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hvl__conb_1 mprj2_logic_high_hvl (
    .HI(mprj2_vdd_logic1_h),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__lsbufhv2lv_1 mprj2_logic_high_lv (
    .A(mprj2_vdd_logic1_h),
    .LVPWR(vccd),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(mprj2_vdd_logic1)
  );
  sky130_fd_sc_hvl__conb_1 mprj_logic_high_hvl (
    .HI(mprj_vdd_logic1_h),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1)
  );
  sky130_fd_sc_hvl__lsbufhv2lv_1 mprj_logic_high_lv (
    .A(mprj_vdd_logic1_h),
    .LVPWR(vccd),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vdda1),
    .VPWR(vdda1),
    .X(mprj_vdd_logic1)
  );
endmodule
