VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1691.030 84.220 1691.350 84.280 ;
        RECT 1713.110 84.220 1713.430 84.280 ;
        RECT 1691.030 84.080 1713.430 84.220 ;
        RECT 1691.030 84.020 1691.350 84.080 ;
        RECT 1713.110 84.020 1713.430 84.080 ;
        RECT 1799.590 84.220 1799.910 84.280 ;
        RECT 1811.090 84.220 1811.410 84.280 ;
        RECT 1799.590 84.080 1811.410 84.220 ;
        RECT 1799.590 84.020 1799.910 84.080 ;
        RECT 1811.090 84.020 1811.410 84.080 ;
        RECT 1896.190 84.220 1896.510 84.280 ;
        RECT 1898.030 84.220 1898.350 84.280 ;
        RECT 1896.190 84.080 1898.350 84.220 ;
        RECT 1896.190 84.020 1896.510 84.080 ;
        RECT 1898.030 84.020 1898.350 84.080 ;
        RECT 1593.970 83.880 1594.290 83.940 ;
        RECT 1607.770 83.880 1608.090 83.940 ;
        RECT 1593.970 83.740 1608.090 83.880 ;
        RECT 1593.970 83.680 1594.290 83.740 ;
        RECT 1607.770 83.680 1608.090 83.740 ;
        RECT 1993.250 83.880 1993.570 83.940 ;
        RECT 2004.290 83.880 2004.610 83.940 ;
        RECT 1993.250 83.740 2004.610 83.880 ;
        RECT 1993.250 83.680 1993.570 83.740 ;
        RECT 2004.290 83.680 2004.610 83.740 ;
        RECT 2089.850 83.880 2090.170 83.940 ;
        RECT 2091.230 83.880 2091.550 83.940 ;
        RECT 2089.850 83.740 2091.550 83.880 ;
        RECT 2089.850 83.680 2090.170 83.740 ;
        RECT 2091.230 83.680 2091.550 83.740 ;
        RECT 869.470 83.540 869.790 83.600 ;
        RECT 917.310 83.540 917.630 83.600 ;
        RECT 869.470 83.400 917.630 83.540 ;
        RECT 869.470 83.340 869.790 83.400 ;
        RECT 917.310 83.340 917.630 83.400 ;
        RECT 2221.870 83.540 2222.190 83.600 ;
        RECT 2236.130 83.540 2236.450 83.600 ;
        RECT 2221.870 83.400 2236.450 83.540 ;
        RECT 2221.870 83.340 2222.190 83.400 ;
        RECT 2236.130 83.340 2236.450 83.400 ;
        RECT 2380.110 83.540 2380.430 83.600 ;
        RECT 2414.610 83.540 2414.930 83.600 ;
        RECT 2380.110 83.400 2414.930 83.540 ;
        RECT 2380.110 83.340 2380.430 83.400 ;
        RECT 2414.610 83.340 2414.930 83.400 ;
      LAYER via ;
        RECT 1691.060 84.020 1691.320 84.280 ;
        RECT 1713.140 84.020 1713.400 84.280 ;
        RECT 1799.620 84.020 1799.880 84.280 ;
        RECT 1811.120 84.020 1811.380 84.280 ;
        RECT 1896.220 84.020 1896.480 84.280 ;
        RECT 1898.060 84.020 1898.320 84.280 ;
        RECT 1594.000 83.680 1594.260 83.940 ;
        RECT 1607.800 83.680 1608.060 83.940 ;
        RECT 1993.280 83.680 1993.540 83.940 ;
        RECT 2004.320 83.680 2004.580 83.940 ;
        RECT 2089.880 83.680 2090.140 83.940 ;
        RECT 2091.260 83.680 2091.520 83.940 ;
        RECT 869.500 83.340 869.760 83.600 ;
        RECT 917.340 83.340 917.600 83.600 ;
        RECT 2221.900 83.340 2222.160 83.600 ;
        RECT 2236.160 83.340 2236.420 83.600 ;
        RECT 2380.140 83.340 2380.400 83.600 ;
        RECT 2414.640 83.340 2414.900 83.600 ;
      LAYER met2 ;
        RECT 756.350 2723.130 756.910 2731.680 ;
        RECT 757.710 2723.130 757.990 2723.245 ;
        RECT 756.350 2722.990 757.990 2723.130 ;
        RECT 756.350 2722.680 756.910 2722.990 ;
        RECT 757.710 2722.875 757.990 2722.990 ;
        RECT 758.630 1185.395 758.910 1185.765 ;
        RECT 758.700 1105.525 758.840 1185.395 ;
        RECT 758.630 1105.155 758.910 1105.525 ;
        RECT 758.170 1031.035 758.450 1031.405 ;
        RECT 758.240 966.125 758.380 1031.035 ;
        RECT 758.170 965.755 758.450 966.125 ;
        RECT 757.250 886.195 757.530 886.565 ;
        RECT 757.320 827.405 757.460 886.195 ;
        RECT 757.250 827.035 757.530 827.405 ;
        RECT 757.710 564.555 757.990 564.925 ;
        RECT 757.780 521.405 757.920 564.555 ;
        RECT 757.710 521.035 757.990 521.405 ;
        RECT 755.410 463.915 755.690 464.285 ;
        RECT 755.480 456.805 755.620 463.915 ;
        RECT 755.410 456.435 755.690 456.805 ;
        RECT 756.790 406.795 757.070 407.165 ;
        RECT 756.860 359.565 757.000 406.795 ;
        RECT 756.790 359.195 757.070 359.565 ;
        RECT 2359.430 85.155 2359.710 85.525 ;
        RECT 2236.150 84.475 2236.430 84.845 ;
        RECT 1691.060 84.165 1691.320 84.310 ;
        RECT 1713.140 84.165 1713.400 84.310 ;
        RECT 1799.620 84.165 1799.880 84.310 ;
        RECT 1811.120 84.165 1811.380 84.310 ;
        RECT 1896.220 84.165 1896.480 84.310 ;
        RECT 1898.060 84.165 1898.320 84.310 ;
        RECT 1510.730 84.050 1511.010 84.165 ;
        RECT 1511.650 84.050 1511.930 84.165 ;
        RECT 1510.730 83.910 1511.930 84.050 ;
        RECT 1510.730 83.795 1511.010 83.910 ;
        RECT 1511.650 83.795 1511.930 83.910 ;
        RECT 1593.990 83.795 1594.270 84.165 ;
        RECT 1607.790 83.795 1608.070 84.165 ;
        RECT 1691.050 83.795 1691.330 84.165 ;
        RECT 1713.130 83.795 1713.410 84.165 ;
        RECT 1799.610 83.795 1799.890 84.165 ;
        RECT 1811.110 83.795 1811.390 84.165 ;
        RECT 1896.210 83.795 1896.490 84.165 ;
        RECT 1898.050 83.795 1898.330 84.165 ;
        RECT 1993.270 83.795 1993.550 84.165 ;
        RECT 2004.310 83.795 2004.590 84.165 ;
        RECT 2089.870 83.795 2090.150 84.165 ;
        RECT 2091.250 83.795 2091.530 84.165 ;
        RECT 2186.010 83.795 2186.290 84.165 ;
        RECT 1594.000 83.650 1594.260 83.795 ;
        RECT 1607.800 83.650 1608.060 83.795 ;
        RECT 1993.280 83.650 1993.540 83.795 ;
        RECT 2004.320 83.650 2004.580 83.795 ;
        RECT 2089.880 83.650 2090.140 83.795 ;
        RECT 2091.260 83.650 2091.520 83.795 ;
        RECT 869.500 83.485 869.760 83.630 ;
        RECT 917.340 83.485 917.600 83.630 ;
        RECT 869.490 83.115 869.770 83.485 ;
        RECT 917.330 83.115 917.610 83.485 ;
        RECT 2186.080 82.125 2186.220 83.795 ;
        RECT 2236.220 83.630 2236.360 84.475 ;
        RECT 2221.900 83.485 2222.160 83.630 ;
        RECT 2221.890 83.115 2222.170 83.485 ;
        RECT 2236.160 83.310 2236.420 83.630 ;
        RECT 2359.500 83.485 2359.640 85.155 ;
        RECT 2414.630 84.475 2414.910 84.845 ;
        RECT 2414.700 83.630 2414.840 84.475 ;
        RECT 2380.140 83.485 2380.400 83.630 ;
        RECT 2359.430 83.115 2359.710 83.485 ;
        RECT 2380.130 83.115 2380.410 83.485 ;
        RECT 2414.640 83.310 2414.900 83.630 ;
        RECT 2186.010 81.755 2186.290 82.125 ;
      LAYER via2 ;
        RECT 757.710 2722.920 757.990 2723.200 ;
        RECT 758.630 1185.440 758.910 1185.720 ;
        RECT 758.630 1105.200 758.910 1105.480 ;
        RECT 758.170 1031.080 758.450 1031.360 ;
        RECT 758.170 965.800 758.450 966.080 ;
        RECT 757.250 886.240 757.530 886.520 ;
        RECT 757.250 827.080 757.530 827.360 ;
        RECT 757.710 564.600 757.990 564.880 ;
        RECT 757.710 521.080 757.990 521.360 ;
        RECT 755.410 463.960 755.690 464.240 ;
        RECT 755.410 456.480 755.690 456.760 ;
        RECT 756.790 406.840 757.070 407.120 ;
        RECT 756.790 359.240 757.070 359.520 ;
        RECT 2359.430 85.200 2359.710 85.480 ;
        RECT 2236.150 84.520 2236.430 84.800 ;
        RECT 1510.730 83.840 1511.010 84.120 ;
        RECT 1511.650 83.840 1511.930 84.120 ;
        RECT 1593.990 83.840 1594.270 84.120 ;
        RECT 1607.790 83.840 1608.070 84.120 ;
        RECT 1691.050 83.840 1691.330 84.120 ;
        RECT 1713.130 83.840 1713.410 84.120 ;
        RECT 1799.610 83.840 1799.890 84.120 ;
        RECT 1811.110 83.840 1811.390 84.120 ;
        RECT 1896.210 83.840 1896.490 84.120 ;
        RECT 1898.050 83.840 1898.330 84.120 ;
        RECT 1993.270 83.840 1993.550 84.120 ;
        RECT 2004.310 83.840 2004.590 84.120 ;
        RECT 2089.870 83.840 2090.150 84.120 ;
        RECT 2091.250 83.840 2091.530 84.120 ;
        RECT 2186.010 83.840 2186.290 84.120 ;
        RECT 869.490 83.160 869.770 83.440 ;
        RECT 917.330 83.160 917.610 83.440 ;
        RECT 2221.890 83.160 2222.170 83.440 ;
        RECT 2414.630 84.520 2414.910 84.800 ;
        RECT 2359.430 83.160 2359.710 83.440 ;
        RECT 2380.130 83.160 2380.410 83.440 ;
        RECT 2186.010 81.800 2186.290 82.080 ;
      LAYER met3 ;
        RECT 757.685 2723.210 758.015 2723.225 ;
        RECT 758.350 2723.210 758.730 2723.220 ;
        RECT 757.685 2722.910 758.730 2723.210 ;
        RECT 757.685 2722.895 758.015 2722.910 ;
        RECT 758.350 2722.900 758.730 2722.910 ;
        RECT 753.750 2560.010 754.130 2560.020 ;
        RECT 757.430 2560.010 757.810 2560.020 ;
        RECT 753.750 2559.710 757.810 2560.010 ;
        RECT 753.750 2559.700 754.130 2559.710 ;
        RECT 757.430 2559.700 757.810 2559.710 ;
        RECT 753.750 2513.090 754.130 2513.100 ;
        RECT 753.750 2512.790 755.930 2513.090 ;
        RECT 753.750 2512.780 754.130 2512.790 ;
        RECT 755.630 2512.420 755.930 2512.790 ;
        RECT 755.590 2512.100 755.970 2512.420 ;
        RECT 757.430 2284.610 757.810 2284.620 ;
        RECT 756.550 2284.310 757.810 2284.610 ;
        RECT 756.550 2283.260 756.850 2284.310 ;
        RECT 757.430 2284.300 757.810 2284.310 ;
        RECT 756.510 2282.940 756.890 2283.260 ;
        RECT 756.510 2236.020 756.890 2236.340 ;
        RECT 756.550 2234.970 756.850 2236.020 ;
        RECT 757.430 2234.970 757.810 2234.980 ;
        RECT 756.550 2234.670 757.810 2234.970 ;
        RECT 757.430 2234.660 757.810 2234.670 ;
        RECT 757.430 2207.460 757.810 2207.780 ;
        RECT 754.670 2207.090 755.050 2207.100 ;
        RECT 757.470 2207.090 757.770 2207.460 ;
        RECT 754.670 2206.790 757.770 2207.090 ;
        RECT 754.670 2206.780 755.050 2206.790 ;
        RECT 754.670 2160.170 755.050 2160.180 ;
        RECT 758.350 2160.170 758.730 2160.180 ;
        RECT 754.670 2159.870 758.730 2160.170 ;
        RECT 754.670 2159.860 755.050 2159.870 ;
        RECT 758.350 2159.860 758.730 2159.870 ;
        RECT 758.350 2139.460 758.730 2139.780 ;
        RECT 758.390 2139.100 758.690 2139.460 ;
        RECT 758.350 2138.780 758.730 2139.100 ;
        RECT 758.350 2118.380 758.730 2118.700 ;
        RECT 758.390 2118.020 758.690 2118.380 ;
        RECT 758.350 2117.700 758.730 2118.020 ;
        RECT 756.510 2062.620 756.890 2062.940 ;
        RECT 756.550 2062.250 756.850 2062.620 ;
        RECT 757.430 2062.250 757.810 2062.260 ;
        RECT 756.550 2061.950 757.810 2062.250 ;
        RECT 757.430 2061.940 757.810 2061.950 ;
        RECT 757.430 2014.340 757.810 2014.660 ;
        RECT 755.590 2013.970 755.970 2013.980 ;
        RECT 757.470 2013.970 757.770 2014.340 ;
        RECT 755.590 2013.670 757.770 2013.970 ;
        RECT 755.590 2013.660 755.970 2013.670 ;
        RECT 755.590 1967.050 755.970 1967.060 ;
        RECT 758.350 1967.050 758.730 1967.060 ;
        RECT 755.590 1966.750 758.730 1967.050 ;
        RECT 755.590 1966.740 755.970 1966.750 ;
        RECT 758.350 1966.740 758.730 1966.750 ;
        RECT 758.350 1946.650 758.730 1946.660 ;
        RECT 757.470 1946.350 758.730 1946.650 ;
        RECT 757.470 1945.300 757.770 1946.350 ;
        RECT 758.350 1946.340 758.730 1946.350 ;
        RECT 757.430 1944.980 757.810 1945.300 ;
        RECT 757.430 1822.210 757.810 1822.220 ;
        RECT 758.350 1822.210 758.730 1822.220 ;
        RECT 757.430 1821.910 758.730 1822.210 ;
        RECT 757.430 1821.900 757.810 1821.910 ;
        RECT 758.350 1821.900 758.730 1821.910 ;
        RECT 758.350 1781.410 758.730 1781.420 ;
        RECT 757.470 1781.110 758.730 1781.410 ;
        RECT 757.470 1780.740 757.770 1781.110 ;
        RECT 758.350 1781.100 758.730 1781.110 ;
        RECT 757.430 1780.420 757.810 1780.740 ;
        RECT 757.430 1742.650 757.810 1742.660 ;
        RECT 761.110 1742.650 761.490 1742.660 ;
        RECT 757.430 1742.350 761.490 1742.650 ;
        RECT 757.430 1742.340 757.810 1742.350 ;
        RECT 761.110 1742.340 761.490 1742.350 ;
        RECT 760.190 1677.370 760.570 1677.380 ;
        RECT 761.110 1677.370 761.490 1677.380 ;
        RECT 760.190 1677.070 761.490 1677.370 ;
        RECT 760.190 1677.060 760.570 1677.070 ;
        RECT 761.110 1677.060 761.490 1677.070 ;
        RECT 760.190 1675.700 760.570 1676.020 ;
        RECT 759.270 1670.570 759.650 1670.580 ;
        RECT 760.230 1670.570 760.530 1675.700 ;
        RECT 759.270 1670.270 760.530 1670.570 ;
        RECT 759.270 1670.260 759.650 1670.270 ;
        RECT 759.270 1637.250 759.650 1637.260 ;
        RECT 757.470 1636.950 759.650 1637.250 ;
        RECT 757.470 1635.900 757.770 1636.950 ;
        RECT 759.270 1636.940 759.650 1636.950 ;
        RECT 757.430 1635.580 757.810 1635.900 ;
        RECT 753.750 1628.410 754.130 1628.420 ;
        RECT 757.430 1628.410 757.810 1628.420 ;
        RECT 753.750 1628.110 757.810 1628.410 ;
        RECT 753.750 1628.100 754.130 1628.110 ;
        RECT 757.430 1628.100 757.810 1628.110 ;
        RECT 753.750 1581.490 754.130 1581.500 ;
        RECT 756.510 1581.490 756.890 1581.500 ;
        RECT 753.750 1581.190 756.890 1581.490 ;
        RECT 753.750 1581.180 754.130 1581.190 ;
        RECT 756.510 1581.180 756.890 1581.190 ;
        RECT 756.510 1580.130 756.890 1580.140 ;
        RECT 757.430 1580.130 757.810 1580.140 ;
        RECT 756.510 1579.830 757.810 1580.130 ;
        RECT 756.510 1579.820 756.890 1579.830 ;
        RECT 757.430 1579.820 757.810 1579.830 ;
        RECT 756.510 1573.330 756.890 1573.340 ;
        RECT 757.430 1573.330 757.810 1573.340 ;
        RECT 756.510 1573.030 757.810 1573.330 ;
        RECT 756.510 1573.020 756.890 1573.030 ;
        RECT 757.430 1573.020 757.810 1573.030 ;
        RECT 755.590 1525.050 755.970 1525.060 ;
        RECT 756.510 1525.050 756.890 1525.060 ;
        RECT 755.590 1524.750 756.890 1525.050 ;
        RECT 755.590 1524.740 755.970 1524.750 ;
        RECT 756.510 1524.740 756.890 1524.750 ;
        RECT 755.590 1484.250 755.970 1484.260 ;
        RECT 758.350 1484.250 758.730 1484.260 ;
        RECT 755.590 1483.950 758.730 1484.250 ;
        RECT 755.590 1483.940 755.970 1483.950 ;
        RECT 758.350 1483.940 758.730 1483.950 ;
        RECT 758.350 1463.850 758.730 1463.860 ;
        RECT 757.470 1463.550 758.730 1463.850 ;
        RECT 757.470 1462.500 757.770 1463.550 ;
        RECT 758.350 1463.540 758.730 1463.550 ;
        RECT 757.430 1462.180 757.810 1462.500 ;
        RECT 755.590 1404.010 755.970 1404.020 ;
        RECT 757.430 1404.010 757.810 1404.020 ;
        RECT 755.590 1403.710 757.810 1404.010 ;
        RECT 755.590 1403.700 755.970 1403.710 ;
        RECT 757.430 1403.700 757.810 1403.710 ;
        RECT 755.590 1380.210 755.970 1380.220 ;
        RECT 757.430 1380.210 757.810 1380.220 ;
        RECT 755.590 1379.910 757.810 1380.210 ;
        RECT 755.590 1379.900 755.970 1379.910 ;
        RECT 757.430 1379.900 757.810 1379.910 ;
        RECT 755.590 1331.250 755.970 1331.260 ;
        RECT 757.430 1331.250 757.810 1331.260 ;
        RECT 755.590 1330.950 757.810 1331.250 ;
        RECT 755.590 1330.940 755.970 1330.950 ;
        RECT 757.430 1330.940 757.810 1330.950 ;
        RECT 755.590 1283.650 755.970 1283.660 ;
        RECT 757.430 1283.650 757.810 1283.660 ;
        RECT 755.590 1283.350 757.810 1283.650 ;
        RECT 755.590 1283.340 755.970 1283.350 ;
        RECT 757.430 1283.340 757.810 1283.350 ;
        RECT 755.590 1234.690 755.970 1234.700 ;
        RECT 757.430 1234.690 757.810 1234.700 ;
        RECT 755.590 1234.390 757.810 1234.690 ;
        RECT 755.590 1234.380 755.970 1234.390 ;
        RECT 757.430 1234.380 757.810 1234.390 ;
        RECT 755.590 1187.090 755.970 1187.100 ;
        RECT 757.430 1187.090 757.810 1187.100 ;
        RECT 755.590 1186.790 757.810 1187.090 ;
        RECT 755.590 1186.780 755.970 1186.790 ;
        RECT 757.430 1186.780 757.810 1186.790 ;
        RECT 757.430 1186.100 757.810 1186.420 ;
        RECT 757.470 1185.730 757.770 1186.100 ;
        RECT 758.605 1185.730 758.935 1185.745 ;
        RECT 757.470 1185.430 758.935 1185.730 ;
        RECT 758.605 1185.415 758.935 1185.430 ;
        RECT 758.605 1105.490 758.935 1105.505 ;
        RECT 757.470 1105.190 758.935 1105.490 ;
        RECT 757.470 1104.820 757.770 1105.190 ;
        RECT 758.605 1105.175 758.935 1105.190 ;
        RECT 757.430 1104.500 757.810 1104.820 ;
        RECT 757.430 1062.340 757.810 1062.660 ;
        RECT 756.510 1061.970 756.890 1061.980 ;
        RECT 757.470 1061.970 757.770 1062.340 ;
        RECT 756.510 1061.670 757.770 1061.970 ;
        RECT 756.510 1061.660 756.890 1061.670 ;
        RECT 756.510 1031.370 756.890 1031.380 ;
        RECT 758.145 1031.370 758.475 1031.385 ;
        RECT 756.510 1031.070 758.475 1031.370 ;
        RECT 756.510 1031.060 756.890 1031.070 ;
        RECT 758.145 1031.055 758.475 1031.070 ;
        RECT 758.145 966.100 758.475 966.105 ;
        RECT 758.145 966.090 758.730 966.100 ;
        RECT 757.920 965.790 758.730 966.090 ;
        RECT 758.145 965.780 758.730 965.790 ;
        RECT 758.145 965.775 758.475 965.780 ;
        RECT 756.510 886.530 756.890 886.540 ;
        RECT 757.225 886.530 757.555 886.545 ;
        RECT 756.510 886.230 757.555 886.530 ;
        RECT 756.510 886.220 756.890 886.230 ;
        RECT 757.225 886.215 757.555 886.230 ;
        RECT 755.590 827.370 755.970 827.380 ;
        RECT 757.225 827.370 757.555 827.385 ;
        RECT 755.590 827.070 757.555 827.370 ;
        RECT 755.590 827.060 755.970 827.070 ;
        RECT 757.225 827.055 757.555 827.070 ;
        RECT 755.590 783.170 755.970 783.180 ;
        RECT 757.430 783.170 757.810 783.180 ;
        RECT 755.590 782.870 757.810 783.170 ;
        RECT 755.590 782.860 755.970 782.870 ;
        RECT 757.430 782.860 757.810 782.870 ;
        RECT 757.430 738.970 757.810 738.980 ;
        RECT 756.550 738.670 757.810 738.970 ;
        RECT 756.550 737.620 756.850 738.670 ;
        RECT 757.430 738.660 757.810 738.670 ;
        RECT 756.510 737.300 756.890 737.620 ;
        RECT 756.510 573.730 756.890 573.740 ;
        RECT 756.510 573.430 757.770 573.730 ;
        RECT 756.510 573.420 756.890 573.430 ;
        RECT 757.470 573.060 757.770 573.430 ;
        RECT 757.430 572.740 757.810 573.060 ;
        RECT 757.430 565.260 757.810 565.580 ;
        RECT 757.470 564.905 757.770 565.260 ;
        RECT 757.470 564.590 758.015 564.905 ;
        RECT 757.685 564.575 758.015 564.590 ;
        RECT 756.510 521.370 756.890 521.380 ;
        RECT 757.685 521.370 758.015 521.385 ;
        RECT 756.510 521.070 758.015 521.370 ;
        RECT 756.510 521.060 756.890 521.070 ;
        RECT 757.685 521.055 758.015 521.070 ;
        RECT 755.385 464.250 755.715 464.265 ;
        RECT 756.510 464.250 756.890 464.260 ;
        RECT 755.385 463.950 756.890 464.250 ;
        RECT 755.385 463.935 755.715 463.950 ;
        RECT 756.510 463.940 756.890 463.950 ;
        RECT 755.385 456.770 755.715 456.785 ;
        RECT 754.710 456.470 755.715 456.770 ;
        RECT 754.710 456.100 755.010 456.470 ;
        RECT 755.385 456.455 755.715 456.470 ;
        RECT 754.670 455.780 755.050 456.100 ;
        RECT 754.670 415.290 755.050 415.300 ;
        RECT 754.670 414.990 756.850 415.290 ;
        RECT 754.670 414.980 755.050 414.990 ;
        RECT 756.550 414.620 756.850 414.990 ;
        RECT 756.510 414.300 756.890 414.620 ;
        RECT 756.765 407.140 757.095 407.145 ;
        RECT 756.510 407.130 757.095 407.140 ;
        RECT 756.310 406.830 757.095 407.130 ;
        RECT 756.510 406.820 757.095 406.830 ;
        RECT 756.765 406.815 757.095 406.820 ;
        RECT 756.765 359.530 757.095 359.545 ;
        RECT 757.430 359.530 757.810 359.540 ;
        RECT 756.765 359.230 757.810 359.530 ;
        RECT 756.765 359.215 757.095 359.230 ;
        RECT 757.430 359.220 757.810 359.230 ;
        RECT 756.510 279.290 756.890 279.300 ;
        RECT 758.350 279.290 758.730 279.300 ;
        RECT 756.510 278.990 758.730 279.290 ;
        RECT 756.510 278.980 756.890 278.990 ;
        RECT 758.350 278.980 758.730 278.990 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 2311.310 85.490 2311.690 85.500 ;
        RECT 2359.405 85.490 2359.735 85.505 ;
        RECT 2311.310 85.190 2359.735 85.490 ;
        RECT 2311.310 85.180 2311.690 85.190 ;
        RECT 2359.405 85.175 2359.735 85.190 ;
        RECT 2236.125 84.810 2236.455 84.825 ;
        RECT 2414.605 84.810 2414.935 84.825 ;
        RECT 1365.590 84.510 1414.650 84.810 ;
        RECT 758.350 83.450 758.730 83.460 ;
        RECT 869.465 83.450 869.795 83.465 ;
        RECT 758.350 83.150 869.795 83.450 ;
        RECT 758.350 83.140 758.730 83.150 ;
        RECT 869.465 83.135 869.795 83.150 ;
        RECT 917.305 83.450 917.635 83.465 ;
        RECT 1365.590 83.450 1365.890 84.510 ;
        RECT 917.305 83.150 1365.890 83.450 ;
        RECT 1414.350 83.450 1414.650 84.510 ;
        RECT 2236.125 84.510 2294.170 84.810 ;
        RECT 2236.125 84.495 2236.455 84.510 ;
        RECT 1510.705 84.130 1511.035 84.145 ;
        RECT 1463.110 83.830 1511.035 84.130 ;
        RECT 1463.110 83.450 1463.410 83.830 ;
        RECT 1510.705 83.815 1511.035 83.830 ;
        RECT 1511.625 84.130 1511.955 84.145 ;
        RECT 1593.965 84.130 1594.295 84.145 ;
        RECT 1511.625 83.830 1559.090 84.130 ;
        RECT 1511.625 83.815 1511.955 83.830 ;
        RECT 1414.350 83.150 1463.410 83.450 ;
        RECT 1558.790 83.450 1559.090 83.830 ;
        RECT 1559.710 83.830 1594.295 84.130 ;
        RECT 1559.710 83.450 1560.010 83.830 ;
        RECT 1593.965 83.815 1594.295 83.830 ;
        RECT 1607.765 84.130 1608.095 84.145 ;
        RECT 1691.025 84.130 1691.355 84.145 ;
        RECT 1607.765 83.830 1641.890 84.130 ;
        RECT 1607.765 83.815 1608.095 83.830 ;
        RECT 1558.790 83.150 1560.010 83.450 ;
        RECT 1641.590 83.450 1641.890 83.830 ;
        RECT 1656.310 83.830 1691.355 84.130 ;
        RECT 1656.310 83.450 1656.610 83.830 ;
        RECT 1691.025 83.815 1691.355 83.830 ;
        RECT 1713.105 84.130 1713.435 84.145 ;
        RECT 1799.585 84.130 1799.915 84.145 ;
        RECT 1713.105 83.830 1752.290 84.130 ;
        RECT 1713.105 83.815 1713.435 83.830 ;
        RECT 1641.590 83.150 1656.610 83.450 ;
        RECT 1751.990 83.450 1752.290 83.830 ;
        RECT 1752.910 83.830 1799.915 84.130 ;
        RECT 1752.910 83.450 1753.210 83.830 ;
        RECT 1799.585 83.815 1799.915 83.830 ;
        RECT 1811.085 84.130 1811.415 84.145 ;
        RECT 1896.185 84.130 1896.515 84.145 ;
        RECT 1811.085 83.830 1835.090 84.130 ;
        RECT 1811.085 83.815 1811.415 83.830 ;
        RECT 1751.990 83.150 1753.210 83.450 ;
        RECT 1834.790 83.450 1835.090 83.830 ;
        RECT 1849.510 83.830 1896.515 84.130 ;
        RECT 1849.510 83.450 1849.810 83.830 ;
        RECT 1896.185 83.815 1896.515 83.830 ;
        RECT 1898.025 84.130 1898.355 84.145 ;
        RECT 1993.245 84.130 1993.575 84.145 ;
        RECT 1898.025 83.830 1945.490 84.130 ;
        RECT 1898.025 83.815 1898.355 83.830 ;
        RECT 1834.790 83.150 1849.810 83.450 ;
        RECT 1945.190 83.450 1945.490 83.830 ;
        RECT 1946.110 83.830 1993.575 84.130 ;
        RECT 1946.110 83.450 1946.410 83.830 ;
        RECT 1993.245 83.815 1993.575 83.830 ;
        RECT 2004.285 84.130 2004.615 84.145 ;
        RECT 2089.845 84.130 2090.175 84.145 ;
        RECT 2004.285 83.830 2028.290 84.130 ;
        RECT 2004.285 83.815 2004.615 83.830 ;
        RECT 1945.190 83.150 1946.410 83.450 ;
        RECT 2027.990 83.450 2028.290 83.830 ;
        RECT 2042.710 83.830 2090.175 84.130 ;
        RECT 2042.710 83.450 2043.010 83.830 ;
        RECT 2089.845 83.815 2090.175 83.830 ;
        RECT 2091.225 84.130 2091.555 84.145 ;
        RECT 2185.985 84.130 2186.315 84.145 ;
        RECT 2091.225 83.830 2124.890 84.130 ;
        RECT 2091.225 83.815 2091.555 83.830 ;
        RECT 2027.990 83.150 2043.010 83.450 ;
        RECT 2124.590 83.450 2124.890 83.830 ;
        RECT 2139.310 83.830 2186.315 84.130 ;
        RECT 2293.870 84.130 2294.170 84.510 ;
        RECT 2414.605 84.510 2449.650 84.810 ;
        RECT 2414.605 84.495 2414.935 84.510 ;
        RECT 2311.310 84.130 2311.690 84.140 ;
        RECT 2293.870 83.830 2311.690 84.130 ;
        RECT 2449.350 84.130 2449.650 84.510 ;
        RECT 2498.110 84.510 2546.250 84.810 ;
        RECT 2449.350 83.830 2497.490 84.130 ;
        RECT 2139.310 83.450 2139.610 83.830 ;
        RECT 2185.985 83.815 2186.315 83.830 ;
        RECT 2311.310 83.820 2311.690 83.830 ;
        RECT 2221.865 83.450 2222.195 83.465 ;
        RECT 2124.590 83.150 2139.610 83.450 ;
        RECT 2221.190 83.150 2222.195 83.450 ;
        RECT 917.305 83.135 917.635 83.150 ;
        RECT 2185.985 82.090 2186.315 82.105 ;
        RECT 2221.190 82.090 2221.490 83.150 ;
        RECT 2221.865 83.135 2222.195 83.150 ;
        RECT 2359.405 83.450 2359.735 83.465 ;
        RECT 2380.105 83.450 2380.435 83.465 ;
        RECT 2359.405 83.150 2380.435 83.450 ;
        RECT 2497.190 83.450 2497.490 83.830 ;
        RECT 2498.110 83.450 2498.410 84.510 ;
        RECT 2545.950 84.130 2546.250 84.510 ;
        RECT 2594.710 84.510 2642.850 84.810 ;
        RECT 2545.950 83.830 2594.090 84.130 ;
        RECT 2497.190 83.150 2498.410 83.450 ;
        RECT 2593.790 83.450 2594.090 83.830 ;
        RECT 2594.710 83.450 2595.010 84.510 ;
        RECT 2642.550 84.130 2642.850 84.510 ;
        RECT 2691.310 84.510 2739.450 84.810 ;
        RECT 2642.550 83.830 2690.690 84.130 ;
        RECT 2593.790 83.150 2595.010 83.450 ;
        RECT 2690.390 83.450 2690.690 83.830 ;
        RECT 2691.310 83.450 2691.610 84.510 ;
        RECT 2739.150 84.130 2739.450 84.510 ;
        RECT 2787.910 84.510 2836.050 84.810 ;
        RECT 2739.150 83.830 2787.290 84.130 ;
        RECT 2690.390 83.150 2691.610 83.450 ;
        RECT 2786.990 83.450 2787.290 83.830 ;
        RECT 2787.910 83.450 2788.210 84.510 ;
        RECT 2835.750 84.130 2836.050 84.510 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2835.750 83.830 2883.890 84.130 ;
        RECT 2786.990 83.150 2788.210 83.450 ;
        RECT 2883.590 83.450 2883.890 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2883.590 83.150 2884.810 83.450 ;
        RECT 2359.405 83.135 2359.735 83.150 ;
        RECT 2380.105 83.135 2380.435 83.150 ;
        RECT 2185.985 81.790 2221.490 82.090 ;
        RECT 2185.985 81.775 2186.315 81.790 ;
      LAYER via3 ;
        RECT 758.380 2722.900 758.700 2723.220 ;
        RECT 753.780 2559.700 754.100 2560.020 ;
        RECT 757.460 2559.700 757.780 2560.020 ;
        RECT 753.780 2512.780 754.100 2513.100 ;
        RECT 755.620 2512.100 755.940 2512.420 ;
        RECT 757.460 2284.300 757.780 2284.620 ;
        RECT 756.540 2282.940 756.860 2283.260 ;
        RECT 756.540 2236.020 756.860 2236.340 ;
        RECT 757.460 2234.660 757.780 2234.980 ;
        RECT 757.460 2207.460 757.780 2207.780 ;
        RECT 754.700 2206.780 755.020 2207.100 ;
        RECT 754.700 2159.860 755.020 2160.180 ;
        RECT 758.380 2159.860 758.700 2160.180 ;
        RECT 758.380 2139.460 758.700 2139.780 ;
        RECT 758.380 2138.780 758.700 2139.100 ;
        RECT 758.380 2118.380 758.700 2118.700 ;
        RECT 758.380 2117.700 758.700 2118.020 ;
        RECT 756.540 2062.620 756.860 2062.940 ;
        RECT 757.460 2061.940 757.780 2062.260 ;
        RECT 757.460 2014.340 757.780 2014.660 ;
        RECT 755.620 2013.660 755.940 2013.980 ;
        RECT 755.620 1966.740 755.940 1967.060 ;
        RECT 758.380 1966.740 758.700 1967.060 ;
        RECT 758.380 1946.340 758.700 1946.660 ;
        RECT 757.460 1944.980 757.780 1945.300 ;
        RECT 757.460 1821.900 757.780 1822.220 ;
        RECT 758.380 1821.900 758.700 1822.220 ;
        RECT 758.380 1781.100 758.700 1781.420 ;
        RECT 757.460 1780.420 757.780 1780.740 ;
        RECT 757.460 1742.340 757.780 1742.660 ;
        RECT 761.140 1742.340 761.460 1742.660 ;
        RECT 760.220 1677.060 760.540 1677.380 ;
        RECT 761.140 1677.060 761.460 1677.380 ;
        RECT 760.220 1675.700 760.540 1676.020 ;
        RECT 759.300 1670.260 759.620 1670.580 ;
        RECT 759.300 1636.940 759.620 1637.260 ;
        RECT 757.460 1635.580 757.780 1635.900 ;
        RECT 753.780 1628.100 754.100 1628.420 ;
        RECT 757.460 1628.100 757.780 1628.420 ;
        RECT 753.780 1581.180 754.100 1581.500 ;
        RECT 756.540 1581.180 756.860 1581.500 ;
        RECT 756.540 1579.820 756.860 1580.140 ;
        RECT 757.460 1579.820 757.780 1580.140 ;
        RECT 756.540 1573.020 756.860 1573.340 ;
        RECT 757.460 1573.020 757.780 1573.340 ;
        RECT 755.620 1524.740 755.940 1525.060 ;
        RECT 756.540 1524.740 756.860 1525.060 ;
        RECT 755.620 1483.940 755.940 1484.260 ;
        RECT 758.380 1483.940 758.700 1484.260 ;
        RECT 758.380 1463.540 758.700 1463.860 ;
        RECT 757.460 1462.180 757.780 1462.500 ;
        RECT 755.620 1403.700 755.940 1404.020 ;
        RECT 757.460 1403.700 757.780 1404.020 ;
        RECT 755.620 1379.900 755.940 1380.220 ;
        RECT 757.460 1379.900 757.780 1380.220 ;
        RECT 755.620 1330.940 755.940 1331.260 ;
        RECT 757.460 1330.940 757.780 1331.260 ;
        RECT 755.620 1283.340 755.940 1283.660 ;
        RECT 757.460 1283.340 757.780 1283.660 ;
        RECT 755.620 1234.380 755.940 1234.700 ;
        RECT 757.460 1234.380 757.780 1234.700 ;
        RECT 755.620 1186.780 755.940 1187.100 ;
        RECT 757.460 1186.780 757.780 1187.100 ;
        RECT 757.460 1186.100 757.780 1186.420 ;
        RECT 757.460 1104.500 757.780 1104.820 ;
        RECT 757.460 1062.340 757.780 1062.660 ;
        RECT 756.540 1061.660 756.860 1061.980 ;
        RECT 756.540 1031.060 756.860 1031.380 ;
        RECT 758.380 965.780 758.700 966.100 ;
        RECT 756.540 886.220 756.860 886.540 ;
        RECT 755.620 827.060 755.940 827.380 ;
        RECT 755.620 782.860 755.940 783.180 ;
        RECT 757.460 782.860 757.780 783.180 ;
        RECT 757.460 738.660 757.780 738.980 ;
        RECT 756.540 737.300 756.860 737.620 ;
        RECT 756.540 573.420 756.860 573.740 ;
        RECT 757.460 572.740 757.780 573.060 ;
        RECT 757.460 565.260 757.780 565.580 ;
        RECT 756.540 521.060 756.860 521.380 ;
        RECT 756.540 463.940 756.860 464.260 ;
        RECT 754.700 455.780 755.020 456.100 ;
        RECT 754.700 414.980 755.020 415.300 ;
        RECT 756.540 414.300 756.860 414.620 ;
        RECT 756.540 406.820 756.860 407.140 ;
        RECT 757.460 359.220 757.780 359.540 ;
        RECT 756.540 278.980 756.860 279.300 ;
        RECT 758.380 278.980 758.700 279.300 ;
        RECT 2311.340 85.180 2311.660 85.500 ;
        RECT 758.380 83.140 758.700 83.460 ;
        RECT 2311.340 83.820 2311.660 84.140 ;
      LAYER met4 ;
        RECT 758.375 2722.895 758.705 2723.225 ;
        RECT 758.390 2670.850 758.690 2722.895 ;
        RECT 757.470 2670.550 758.690 2670.850 ;
        RECT 757.470 2560.025 757.770 2670.550 ;
        RECT 753.775 2559.695 754.105 2560.025 ;
        RECT 757.455 2559.695 757.785 2560.025 ;
        RECT 753.790 2513.105 754.090 2559.695 ;
        RECT 753.775 2512.775 754.105 2513.105 ;
        RECT 755.615 2512.095 755.945 2512.425 ;
        RECT 755.630 2477.050 755.930 2512.095 ;
        RECT 755.630 2476.750 756.850 2477.050 ;
        RECT 756.550 2426.050 756.850 2476.750 ;
        RECT 756.550 2425.750 757.770 2426.050 ;
        RECT 757.470 2284.625 757.770 2425.750 ;
        RECT 757.455 2284.295 757.785 2284.625 ;
        RECT 756.535 2282.935 756.865 2283.265 ;
        RECT 756.550 2236.345 756.850 2282.935 ;
        RECT 756.535 2236.015 756.865 2236.345 ;
        RECT 757.455 2234.655 757.785 2234.985 ;
        RECT 757.470 2207.785 757.770 2234.655 ;
        RECT 757.455 2207.455 757.785 2207.785 ;
        RECT 754.695 2206.775 755.025 2207.105 ;
        RECT 754.710 2160.185 755.010 2206.775 ;
        RECT 754.695 2159.855 755.025 2160.185 ;
        RECT 758.375 2159.855 758.705 2160.185 ;
        RECT 758.390 2139.785 758.690 2159.855 ;
        RECT 758.375 2139.455 758.705 2139.785 ;
        RECT 758.375 2138.775 758.705 2139.105 ;
        RECT 758.390 2118.705 758.690 2138.775 ;
        RECT 758.375 2118.375 758.705 2118.705 ;
        RECT 758.375 2117.695 758.705 2118.025 ;
        RECT 758.390 2089.450 758.690 2117.695 ;
        RECT 756.550 2089.150 758.690 2089.450 ;
        RECT 756.550 2062.945 756.850 2089.150 ;
        RECT 756.535 2062.615 756.865 2062.945 ;
        RECT 757.455 2061.935 757.785 2062.265 ;
        RECT 757.470 2014.665 757.770 2061.935 ;
        RECT 757.455 2014.335 757.785 2014.665 ;
        RECT 755.615 2013.655 755.945 2013.985 ;
        RECT 755.630 1967.065 755.930 2013.655 ;
        RECT 755.615 1966.735 755.945 1967.065 ;
        RECT 758.375 1966.735 758.705 1967.065 ;
        RECT 758.390 1946.665 758.690 1966.735 ;
        RECT 758.375 1946.335 758.705 1946.665 ;
        RECT 757.455 1944.975 757.785 1945.305 ;
        RECT 757.470 1822.225 757.770 1944.975 ;
        RECT 757.455 1821.895 757.785 1822.225 ;
        RECT 758.375 1821.895 758.705 1822.225 ;
        RECT 758.390 1781.425 758.690 1821.895 ;
        RECT 758.375 1781.095 758.705 1781.425 ;
        RECT 757.455 1780.415 757.785 1780.745 ;
        RECT 757.470 1742.665 757.770 1780.415 ;
        RECT 757.455 1742.335 757.785 1742.665 ;
        RECT 761.135 1742.335 761.465 1742.665 ;
        RECT 761.150 1677.385 761.450 1742.335 ;
        RECT 760.215 1677.055 760.545 1677.385 ;
        RECT 761.135 1677.055 761.465 1677.385 ;
        RECT 760.230 1676.025 760.530 1677.055 ;
        RECT 760.215 1675.695 760.545 1676.025 ;
        RECT 759.295 1670.255 759.625 1670.585 ;
        RECT 759.310 1637.265 759.610 1670.255 ;
        RECT 759.295 1636.935 759.625 1637.265 ;
        RECT 757.455 1635.575 757.785 1635.905 ;
        RECT 757.470 1628.425 757.770 1635.575 ;
        RECT 753.775 1628.095 754.105 1628.425 ;
        RECT 757.455 1628.095 757.785 1628.425 ;
        RECT 753.790 1581.505 754.090 1628.095 ;
        RECT 753.775 1581.175 754.105 1581.505 ;
        RECT 756.535 1581.175 756.865 1581.505 ;
        RECT 756.550 1580.145 756.850 1581.175 ;
        RECT 756.535 1579.815 756.865 1580.145 ;
        RECT 757.455 1579.815 757.785 1580.145 ;
        RECT 757.470 1573.345 757.770 1579.815 ;
        RECT 756.535 1573.015 756.865 1573.345 ;
        RECT 757.455 1573.015 757.785 1573.345 ;
        RECT 756.550 1525.065 756.850 1573.015 ;
        RECT 755.615 1524.735 755.945 1525.065 ;
        RECT 756.535 1524.735 756.865 1525.065 ;
        RECT 755.630 1484.265 755.930 1524.735 ;
        RECT 755.615 1483.935 755.945 1484.265 ;
        RECT 758.375 1483.935 758.705 1484.265 ;
        RECT 758.390 1463.865 758.690 1483.935 ;
        RECT 758.375 1463.535 758.705 1463.865 ;
        RECT 757.455 1462.175 757.785 1462.505 ;
        RECT 757.470 1404.025 757.770 1462.175 ;
        RECT 755.615 1403.695 755.945 1404.025 ;
        RECT 757.455 1403.695 757.785 1404.025 ;
        RECT 755.630 1380.225 755.930 1403.695 ;
        RECT 755.615 1379.895 755.945 1380.225 ;
        RECT 757.455 1379.895 757.785 1380.225 ;
        RECT 757.470 1331.265 757.770 1379.895 ;
        RECT 755.615 1330.935 755.945 1331.265 ;
        RECT 757.455 1330.935 757.785 1331.265 ;
        RECT 755.630 1283.665 755.930 1330.935 ;
        RECT 755.615 1283.335 755.945 1283.665 ;
        RECT 757.455 1283.335 757.785 1283.665 ;
        RECT 757.470 1234.705 757.770 1283.335 ;
        RECT 755.615 1234.375 755.945 1234.705 ;
        RECT 757.455 1234.375 757.785 1234.705 ;
        RECT 755.630 1187.105 755.930 1234.375 ;
        RECT 755.615 1186.775 755.945 1187.105 ;
        RECT 757.455 1186.775 757.785 1187.105 ;
        RECT 757.470 1186.425 757.770 1186.775 ;
        RECT 757.455 1186.095 757.785 1186.425 ;
        RECT 757.455 1104.495 757.785 1104.825 ;
        RECT 757.470 1062.665 757.770 1104.495 ;
        RECT 757.455 1062.335 757.785 1062.665 ;
        RECT 756.535 1061.655 756.865 1061.985 ;
        RECT 756.550 1031.385 756.850 1061.655 ;
        RECT 756.535 1031.055 756.865 1031.385 ;
        RECT 758.375 965.775 758.705 966.105 ;
        RECT 758.390 940.250 758.690 965.775 ;
        RECT 756.550 939.950 758.690 940.250 ;
        RECT 756.550 886.545 756.850 939.950 ;
        RECT 756.535 886.215 756.865 886.545 ;
        RECT 755.615 827.055 755.945 827.385 ;
        RECT 755.630 783.185 755.930 827.055 ;
        RECT 755.615 782.855 755.945 783.185 ;
        RECT 757.455 782.855 757.785 783.185 ;
        RECT 757.470 738.985 757.770 782.855 ;
        RECT 757.455 738.655 757.785 738.985 ;
        RECT 756.535 737.295 756.865 737.625 ;
        RECT 756.550 573.745 756.850 737.295 ;
        RECT 756.535 573.415 756.865 573.745 ;
        RECT 757.455 572.735 757.785 573.065 ;
        RECT 757.470 565.585 757.770 572.735 ;
        RECT 757.455 565.255 757.785 565.585 ;
        RECT 756.535 521.055 756.865 521.385 ;
        RECT 756.550 464.265 756.850 521.055 ;
        RECT 756.535 463.935 756.865 464.265 ;
        RECT 754.695 455.775 755.025 456.105 ;
        RECT 754.710 415.305 755.010 455.775 ;
        RECT 754.695 414.975 755.025 415.305 ;
        RECT 756.535 414.295 756.865 414.625 ;
        RECT 756.550 407.145 756.850 414.295 ;
        RECT 756.535 406.815 756.865 407.145 ;
        RECT 757.455 359.215 757.785 359.545 ;
        RECT 757.470 348.650 757.770 359.215 ;
        RECT 756.550 348.350 757.770 348.650 ;
        RECT 756.550 279.305 756.850 348.350 ;
        RECT 756.535 278.975 756.865 279.305 ;
        RECT 758.375 278.975 758.705 279.305 ;
        RECT 758.390 165.050 758.690 278.975 ;
        RECT 758.390 164.750 759.610 165.050 ;
        RECT 759.310 117.450 759.610 164.750 ;
        RECT 758.390 117.150 759.610 117.450 ;
        RECT 758.390 83.465 758.690 117.150 ;
        RECT 2311.335 85.175 2311.665 85.505 ;
        RECT 2311.350 84.145 2311.650 85.175 ;
        RECT 2311.335 83.815 2311.665 84.145 ;
        RECT 758.375 83.135 758.705 83.465 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.010 2724.320 1145.330 2724.380 ;
        RECT 2248.550 2724.320 2248.870 2724.380 ;
        RECT 1145.010 2724.180 2248.870 2724.320 ;
        RECT 1145.010 2724.120 1145.330 2724.180 ;
        RECT 2248.550 2724.120 2248.870 2724.180 ;
        RECT 2248.550 2435.660 2248.870 2435.720 ;
        RECT 2900.370 2435.660 2900.690 2435.720 ;
        RECT 2248.550 2435.520 2900.690 2435.660 ;
        RECT 2248.550 2435.460 2248.870 2435.520 ;
        RECT 2900.370 2435.460 2900.690 2435.520 ;
      LAYER via ;
        RECT 1145.040 2724.120 1145.300 2724.380 ;
        RECT 2248.580 2724.120 2248.840 2724.380 ;
        RECT 2248.580 2435.460 2248.840 2435.720 ;
        RECT 2900.400 2435.460 2900.660 2435.720 ;
      LAYER met2 ;
        RECT 1144.130 2724.490 1144.690 2731.680 ;
        RECT 1144.130 2724.410 1145.240 2724.490 ;
        RECT 1144.130 2724.350 1145.300 2724.410 ;
        RECT 1144.130 2722.680 1144.690 2724.350 ;
        RECT 1145.040 2724.090 1145.300 2724.350 ;
        RECT 2248.580 2724.090 2248.840 2724.410 ;
        RECT 2248.640 2435.750 2248.780 2724.090 ;
        RECT 2248.580 2435.430 2248.840 2435.750 ;
        RECT 2900.400 2435.430 2900.660 2435.750 ;
        RECT 2900.460 2434.245 2900.600 2435.430 ;
        RECT 2900.390 2433.875 2900.670 2434.245 ;
      LAYER via2 ;
        RECT 2900.390 2433.920 2900.670 2434.200 ;
      LAYER met3 ;
        RECT 2900.365 2434.210 2900.695 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.365 2433.910 2924.800 2434.210 ;
        RECT 2900.365 2433.895 2900.695 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1184.570 2724.660 1184.890 2724.720 ;
        RECT 2245.330 2724.660 2245.650 2724.720 ;
        RECT 1184.570 2724.520 2245.650 2724.660 ;
        RECT 1184.570 2724.460 1184.890 2724.520 ;
        RECT 2245.330 2724.460 2245.650 2724.520 ;
        RECT 2245.330 2670.260 2245.650 2670.320 ;
        RECT 2899.450 2670.260 2899.770 2670.320 ;
        RECT 2245.330 2670.120 2899.770 2670.260 ;
        RECT 2245.330 2670.060 2245.650 2670.120 ;
        RECT 2899.450 2670.060 2899.770 2670.120 ;
      LAYER via ;
        RECT 1184.600 2724.460 1184.860 2724.720 ;
        RECT 2245.360 2724.460 2245.620 2724.720 ;
        RECT 2245.360 2670.060 2245.620 2670.320 ;
        RECT 2899.480 2670.060 2899.740 2670.320 ;
      LAYER met2 ;
        RECT 1182.770 2724.490 1183.330 2731.680 ;
        RECT 1184.600 2724.490 1184.860 2724.750 ;
        RECT 1182.770 2724.430 1184.860 2724.490 ;
        RECT 2245.360 2724.430 2245.620 2724.750 ;
        RECT 1182.770 2724.350 1184.800 2724.430 ;
        RECT 1182.770 2722.680 1183.330 2724.350 ;
        RECT 2245.420 2670.350 2245.560 2724.430 ;
        RECT 2245.360 2670.030 2245.620 2670.350 ;
        RECT 2899.480 2670.030 2899.740 2670.350 ;
        RECT 2899.540 2669.525 2899.680 2670.030 ;
        RECT 2899.470 2669.155 2899.750 2669.525 ;
      LAYER via2 ;
        RECT 2899.470 2669.200 2899.750 2669.480 ;
      LAYER met3 ;
        RECT 2899.445 2669.490 2899.775 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2899.445 2669.190 2924.800 2669.490 ;
        RECT 2899.445 2669.175 2899.775 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.810 2898.400 1228.130 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1227.810 2898.260 2901.150 2898.400 ;
        RECT 1227.810 2898.200 1228.130 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1227.840 2898.200 1228.100 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1227.840 2898.170 1228.100 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1227.900 2731.970 1228.040 2898.170 ;
        RECT 1224.680 2731.830 1228.040 2731.970 ;
        RECT 1221.870 2731.290 1222.430 2731.680 ;
        RECT 1224.680 2731.290 1224.820 2731.830 ;
        RECT 1221.870 2731.150 1224.820 2731.290 ;
        RECT 1221.870 2722.680 1222.430 2731.150 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 3133.000 1262.630 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1262.310 3132.860 2901.150 3133.000 ;
        RECT 1262.310 3132.800 1262.630 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1262.340 3132.800 1262.600 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1262.340 3132.770 1262.600 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1260.510 2731.290 1261.070 2731.680 ;
        RECT 1262.400 2731.290 1262.540 3132.770 ;
        RECT 1260.510 2731.150 1262.540 2731.290 ;
        RECT 1260.510 2722.680 1261.070 2731.150 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1303.710 3367.600 1304.030 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1303.710 3367.460 2901.150 3367.600 ;
        RECT 1303.710 3367.400 1304.030 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1303.740 3367.400 1304.000 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1303.740 3367.370 1304.000 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1303.800 2731.970 1303.940 3367.370 ;
        RECT 1301.500 2731.830 1303.940 2731.970 ;
        RECT 1299.150 2730.610 1299.710 2731.680 ;
        RECT 1301.500 2730.610 1301.640 2731.830 ;
        RECT 1299.150 2730.470 1301.640 2730.610 ;
        RECT 1299.150 2722.680 1299.710 2730.470 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2795.565 3008.405 2795.735 3042.915 ;
        RECT 2796.485 2946.525 2796.655 2994.635 ;
        RECT 2795.105 2753.065 2795.275 2801.175 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2795.565 3042.745 2795.735 3042.915 ;
        RECT 2796.485 2994.465 2796.655 2994.635 ;
        RECT 2795.105 2801.005 2795.275 2801.175 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.295 3042.760 2795.810 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.505 3008.560 2795.795 3008.605 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.505 3008.420 2796.730 3008.560 ;
        RECT 2795.505 3008.375 2795.795 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2796.215 2994.480 2796.730 2994.620 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2796.425 2946.680 2796.715 2946.725 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2796.425 2946.540 2797.190 2946.680 ;
        RECT 2796.425 2946.495 2796.715 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2815.580 2795.350 2815.840 ;
        RECT 2795.120 2815.160 2795.260 2815.580 ;
        RECT 2795.030 2814.900 2795.350 2815.160 ;
        RECT 2795.030 2801.160 2795.350 2801.220 ;
        RECT 2794.835 2801.020 2795.350 2801.160 ;
        RECT 2795.030 2800.960 2795.350 2801.020 ;
        RECT 2795.045 2753.220 2795.335 2753.265 ;
        RECT 2795.490 2753.220 2795.810 2753.280 ;
        RECT 2795.045 2753.080 2795.810 2753.220 ;
        RECT 2795.045 2753.035 2795.335 2753.080 ;
        RECT 2795.490 2753.020 2795.810 2753.080 ;
        RECT 1338.210 2749.480 1338.530 2749.540 ;
        RECT 2795.490 2749.480 2795.810 2749.540 ;
        RECT 1338.210 2749.340 2795.810 2749.480 ;
        RECT 1338.210 2749.280 1338.530 2749.340 ;
        RECT 2795.490 2749.280 2795.810 2749.340 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2815.580 2795.320 2815.840 ;
        RECT 2795.060 2814.900 2795.320 2815.160 ;
        RECT 2795.060 2800.960 2795.320 2801.220 ;
        RECT 2795.520 2753.020 2795.780 2753.280 ;
        RECT 1338.240 2749.280 1338.500 2749.540 ;
        RECT 2795.520 2749.280 2795.780 2749.540 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2849.610 2795.720 2863.070 ;
        RECT 2795.120 2849.470 2795.720 2849.610 ;
        RECT 2795.120 2815.870 2795.260 2849.470 ;
        RECT 2795.060 2815.550 2795.320 2815.870 ;
        RECT 2795.060 2814.870 2795.320 2815.190 ;
        RECT 2795.120 2801.250 2795.260 2814.870 ;
        RECT 2795.060 2800.930 2795.320 2801.250 ;
        RECT 2795.520 2752.990 2795.780 2753.310 ;
        RECT 2795.580 2749.570 2795.720 2752.990 ;
        RECT 1338.240 2749.250 1338.500 2749.570 ;
        RECT 2795.520 2749.250 2795.780 2749.570 ;
        RECT 1338.300 2731.680 1338.440 2749.250 ;
        RECT 1338.250 2722.680 1338.810 2731.680 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2469.350 2946.340 2469.670 2946.400 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2469.350 2946.200 2471.050 2946.340 ;
        RECT 2469.350 2946.140 2469.670 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 1376.850 2749.820 1377.170 2749.880 ;
        RECT 2470.270 2749.820 2470.590 2749.880 ;
        RECT 1376.850 2749.680 2470.590 2749.820 ;
        RECT 1376.850 2749.620 1377.170 2749.680 ;
        RECT 2470.270 2749.620 2470.590 2749.680 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2469.380 2946.140 2469.640 2946.400 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 1376.880 2749.620 1377.140 2749.880 ;
        RECT 2470.300 2749.620 2470.560 2749.880 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2469.380 2946.110 2469.640 2946.430 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2469.440 2898.685 2469.580 2946.110 ;
        RECT 2469.370 2898.315 2469.650 2898.685 ;
        RECT 2470.290 2898.315 2470.570 2898.685 ;
        RECT 2470.360 2863.210 2470.500 2898.315 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2815.610 2470.960 2863.070 ;
        RECT 2470.820 2815.470 2471.420 2815.610 ;
        RECT 2471.280 2787.730 2471.420 2815.470 ;
        RECT 2470.360 2787.590 2471.420 2787.730 ;
        RECT 2470.360 2749.910 2470.500 2787.590 ;
        RECT 1376.880 2749.590 1377.140 2749.910 ;
        RECT 2470.300 2749.590 2470.560 2749.910 ;
        RECT 1376.940 2731.680 1377.080 2749.590 ;
        RECT 1376.890 2722.680 1377.450 2731.680 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
        RECT 2469.370 2898.360 2469.650 2898.640 ;
        RECT 2470.290 2898.360 2470.570 2898.640 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
        RECT 2469.345 2898.650 2469.675 2898.665 ;
        RECT 2470.265 2898.650 2470.595 2898.665 ;
        RECT 2469.345 2898.350 2470.595 2898.650 ;
        RECT 2469.345 2898.335 2469.675 2898.350 ;
        RECT 2470.265 2898.335 2470.595 2898.350 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2146.965 3008.405 2147.135 3042.915 ;
        RECT 2147.885 2946.525 2148.055 2994.635 ;
        RECT 2146.045 2753.065 2146.215 2767.175 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2146.965 3042.745 2147.135 3042.915 ;
        RECT 2147.885 2994.465 2148.055 2994.635 ;
        RECT 2146.045 2767.005 2146.215 2767.175 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.695 3042.760 2147.210 3042.900 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.905 3008.560 2147.195 3008.605 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.905 3008.420 2148.130 3008.560 ;
        RECT 2146.905 3008.375 2147.195 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2147.615 2994.480 2148.130 2994.620 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 2146.430 2815.580 2146.750 2815.840 ;
        RECT 2146.520 2815.160 2146.660 2815.580 ;
        RECT 2146.430 2814.900 2146.750 2815.160 ;
        RECT 2145.970 2767.160 2146.290 2767.220 ;
        RECT 2145.775 2767.020 2146.290 2767.160 ;
        RECT 2145.970 2766.960 2146.290 2767.020 ;
        RECT 2145.970 2753.220 2146.290 2753.280 ;
        RECT 2145.775 2753.080 2146.290 2753.220 ;
        RECT 2145.970 2753.020 2146.290 2753.080 ;
        RECT 1415.490 2750.160 1415.810 2750.220 ;
        RECT 2145.970 2750.160 2146.290 2750.220 ;
        RECT 1415.490 2750.020 2146.290 2750.160 ;
        RECT 1415.490 2749.960 1415.810 2750.020 ;
        RECT 2145.970 2749.960 2146.290 2750.020 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 2146.460 2815.580 2146.720 2815.840 ;
        RECT 2146.460 2814.900 2146.720 2815.160 ;
        RECT 2146.000 2766.960 2146.260 2767.220 ;
        RECT 2146.000 2753.020 2146.260 2753.280 ;
        RECT 1415.520 2749.960 1415.780 2750.220 ;
        RECT 2146.000 2749.960 2146.260 2750.220 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2912.430 2148.500 2946.450 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2849.610 2147.120 2863.070 ;
        RECT 2146.520 2849.470 2147.120 2849.610 ;
        RECT 2146.520 2815.870 2146.660 2849.470 ;
        RECT 2146.460 2815.550 2146.720 2815.870 ;
        RECT 2146.460 2814.870 2146.720 2815.190 ;
        RECT 2146.520 2801.330 2146.660 2814.870 ;
        RECT 2146.060 2801.190 2146.660 2801.330 ;
        RECT 2146.060 2767.250 2146.200 2801.190 ;
        RECT 2146.000 2766.930 2146.260 2767.250 ;
        RECT 2146.000 2752.990 2146.260 2753.310 ;
        RECT 2146.060 2750.250 2146.200 2752.990 ;
        RECT 1415.520 2749.930 1415.780 2750.250 ;
        RECT 2146.000 2749.930 2146.260 2750.250 ;
        RECT 1415.580 2731.680 1415.720 2749.930 ;
        RECT 1415.530 2722.680 1416.090 2731.680 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1821.745 3332.765 1821.915 3380.875 ;
      LAYER mcon ;
        RECT 1821.745 3380.705 1821.915 3380.875 ;
      LAYER met1 ;
        RECT 1821.670 3380.860 1821.990 3380.920 ;
        RECT 1821.475 3380.720 1821.990 3380.860 ;
        RECT 1821.670 3380.660 1821.990 3380.720 ;
        RECT 1821.685 3332.920 1821.975 3332.965 ;
        RECT 1822.130 3332.920 1822.450 3332.980 ;
        RECT 1821.685 3332.780 1822.450 3332.920 ;
        RECT 1821.685 3332.735 1821.975 3332.780 ;
        RECT 1822.130 3332.720 1822.450 3332.780 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1821.670 2981.020 1821.990 2981.080 ;
        RECT 1822.590 2981.020 1822.910 2981.080 ;
        RECT 1821.670 2980.880 1822.910 2981.020 ;
        RECT 1821.670 2980.820 1821.990 2980.880 ;
        RECT 1822.590 2980.820 1822.910 2980.880 ;
        RECT 1820.750 2946.340 1821.070 2946.400 ;
        RECT 1822.130 2946.340 1822.450 2946.400 ;
        RECT 1820.750 2946.200 1822.450 2946.340 ;
        RECT 1820.750 2946.140 1821.070 2946.200 ;
        RECT 1822.130 2946.140 1822.450 2946.200 ;
        RECT 1454.590 2750.500 1454.910 2750.560 ;
        RECT 1821.670 2750.500 1821.990 2750.560 ;
        RECT 1454.590 2750.360 1821.990 2750.500 ;
        RECT 1454.590 2750.300 1454.910 2750.360 ;
        RECT 1821.670 2750.300 1821.990 2750.360 ;
      LAYER via ;
        RECT 1821.700 3380.660 1821.960 3380.920 ;
        RECT 1822.160 3332.720 1822.420 3332.980 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1821.700 2980.820 1821.960 2981.080 ;
        RECT 1822.620 2980.820 1822.880 2981.080 ;
        RECT 1820.780 2946.140 1821.040 2946.400 ;
        RECT 1822.160 2946.140 1822.420 2946.400 ;
        RECT 1454.620 2750.300 1454.880 2750.560 ;
        RECT 1821.700 2750.300 1821.960 2750.560 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3430.445 1825.580 3517.230 ;
        RECT 1825.370 3430.075 1825.650 3430.445 ;
        RECT 1822.610 3429.395 1822.890 3429.765 ;
        RECT 1822.680 3394.970 1822.820 3429.395 ;
        RECT 1821.760 3394.830 1822.820 3394.970 ;
        RECT 1821.760 3380.950 1821.900 3394.830 ;
        RECT 1821.700 3380.630 1821.960 3380.950 ;
        RECT 1822.160 3332.690 1822.420 3333.010 ;
        RECT 1822.220 3298.410 1822.360 3332.690 ;
        RECT 1822.220 3298.270 1822.820 3298.410 ;
        RECT 1822.680 3270.790 1822.820 3298.270 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 2981.110 1822.820 3028.990 ;
        RECT 1821.700 2980.850 1821.960 2981.110 ;
        RECT 1821.700 2980.790 1822.360 2980.850 ;
        RECT 1822.620 2980.790 1822.880 2981.110 ;
        RECT 1821.760 2980.710 1822.360 2980.790 ;
        RECT 1822.220 2980.170 1822.360 2980.710 ;
        RECT 1822.220 2980.030 1822.820 2980.170 ;
        RECT 1822.680 2959.770 1822.820 2980.030 ;
        RECT 1822.220 2959.630 1822.820 2959.770 ;
        RECT 1822.220 2946.430 1822.360 2959.630 ;
        RECT 1820.780 2946.110 1821.040 2946.430 ;
        RECT 1822.160 2946.110 1822.420 2946.430 ;
        RECT 1820.840 2898.685 1820.980 2946.110 ;
        RECT 1820.770 2898.315 1821.050 2898.685 ;
        RECT 1821.690 2898.315 1821.970 2898.685 ;
        RECT 1821.760 2863.210 1821.900 2898.315 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2815.610 1822.360 2863.070 ;
        RECT 1822.220 2815.470 1822.820 2815.610 ;
        RECT 1822.680 2787.730 1822.820 2815.470 ;
        RECT 1821.760 2787.590 1822.820 2787.730 ;
        RECT 1821.760 2750.590 1821.900 2787.590 ;
        RECT 1454.620 2750.270 1454.880 2750.590 ;
        RECT 1821.700 2750.270 1821.960 2750.590 ;
        RECT 1454.680 2731.680 1454.820 2750.270 ;
        RECT 1454.630 2722.680 1455.190 2731.680 ;
      LAYER via2 ;
        RECT 1825.370 3430.120 1825.650 3430.400 ;
        RECT 1822.610 3429.440 1822.890 3429.720 ;
        RECT 1820.770 2898.360 1821.050 2898.640 ;
        RECT 1821.690 2898.360 1821.970 2898.640 ;
      LAYER met3 ;
        RECT 1825.345 3430.410 1825.675 3430.425 ;
        RECT 1821.910 3430.110 1825.675 3430.410 ;
        RECT 1821.910 3429.730 1822.210 3430.110 ;
        RECT 1825.345 3430.095 1825.675 3430.110 ;
        RECT 1822.585 3429.730 1822.915 3429.745 ;
        RECT 1821.910 3429.430 1822.915 3429.730 ;
        RECT 1822.585 3429.415 1822.915 3429.430 ;
        RECT 1820.745 2898.650 1821.075 2898.665 ;
        RECT 1821.665 2898.650 1821.995 2898.665 ;
        RECT 1820.745 2898.350 1821.995 2898.650 ;
        RECT 1820.745 2898.335 1821.075 2898.350 ;
        RECT 1821.665 2898.335 1821.995 2898.350 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 3332.765 1499.455 3422.355 ;
        RECT 1498.365 3008.405 1498.535 3042.915 ;
        RECT 1499.285 2946.525 1499.455 2994.635 ;
        RECT 1497.905 2753.065 1498.075 2801.175 ;
      LAYER mcon ;
        RECT 1499.285 3422.185 1499.455 3422.355 ;
        RECT 1498.365 3042.745 1498.535 3042.915 ;
        RECT 1499.285 2994.465 1499.455 2994.635 ;
        RECT 1497.905 2801.005 1498.075 2801.175 ;
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1499.225 3422.340 1499.515 3422.385 ;
        RECT 1497.830 3422.200 1499.515 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1499.225 3422.155 1499.515 3422.200 ;
        RECT 1499.225 3332.920 1499.515 3332.965 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1499.225 3332.780 1499.990 3332.920 ;
        RECT 1499.225 3332.735 1499.515 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1498.095 3042.760 1498.610 3042.900 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1498.305 3008.560 1498.595 3008.605 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1498.305 3008.420 1499.530 3008.560 ;
        RECT 1498.305 3008.375 1498.595 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1499.015 2994.480 1499.530 2994.620 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1499.225 2946.680 1499.515 2946.725 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1499.225 2946.540 1499.990 2946.680 ;
        RECT 1499.225 2946.495 1499.515 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 1497.830 2815.580 1498.150 2815.840 ;
        RECT 1497.920 2815.160 1498.060 2815.580 ;
        RECT 1497.830 2814.900 1498.150 2815.160 ;
        RECT 1497.830 2801.160 1498.150 2801.220 ;
        RECT 1497.635 2801.020 1498.150 2801.160 ;
        RECT 1497.830 2800.960 1498.150 2801.020 ;
        RECT 1497.845 2753.220 1498.135 2753.265 ;
        RECT 1498.290 2753.220 1498.610 2753.280 ;
        RECT 1497.845 2753.080 1498.610 2753.220 ;
        RECT 1497.845 2753.035 1498.135 2753.080 ;
        RECT 1498.290 2753.020 1498.610 2753.080 ;
        RECT 1493.230 2746.420 1493.550 2746.480 ;
        RECT 1497.830 2746.420 1498.150 2746.480 ;
        RECT 1493.230 2746.280 1498.150 2746.420 ;
        RECT 1493.230 2746.220 1493.550 2746.280 ;
        RECT 1497.830 2746.220 1498.150 2746.280 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 1497.860 2815.580 1498.120 2815.840 ;
        RECT 1497.860 2814.900 1498.120 2815.160 ;
        RECT 1497.860 2800.960 1498.120 2801.220 ;
        RECT 1498.320 2753.020 1498.580 2753.280 ;
        RECT 1493.260 2746.220 1493.520 2746.480 ;
        RECT 1497.860 2746.220 1498.120 2746.480 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3443.170 1500.820 3517.600 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3236.450 1498.980 3298.270 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2849.610 1498.520 2863.070 ;
        RECT 1497.920 2849.470 1498.520 2849.610 ;
        RECT 1497.920 2815.870 1498.060 2849.470 ;
        RECT 1497.860 2815.550 1498.120 2815.870 ;
        RECT 1497.860 2814.870 1498.120 2815.190 ;
        RECT 1497.920 2802.805 1498.060 2814.870 ;
        RECT 1497.850 2802.435 1498.130 2802.805 ;
        RECT 1497.850 2801.755 1498.130 2802.125 ;
        RECT 1497.920 2801.250 1498.060 2801.755 ;
        RECT 1497.860 2800.930 1498.120 2801.250 ;
        RECT 1498.380 2753.310 1498.520 2753.465 ;
        RECT 1498.320 2753.050 1498.580 2753.310 ;
        RECT 1497.920 2752.990 1498.580 2753.050 ;
        RECT 1497.920 2752.910 1498.520 2752.990 ;
        RECT 1497.920 2746.510 1498.060 2752.910 ;
        RECT 1493.260 2746.190 1493.520 2746.510 ;
        RECT 1497.860 2746.190 1498.120 2746.510 ;
        RECT 1493.320 2731.680 1493.460 2746.190 ;
        RECT 1493.270 2722.680 1493.830 2731.680 ;
      LAYER via2 ;
        RECT 1497.850 2802.480 1498.130 2802.760 ;
        RECT 1497.850 2801.800 1498.130 2802.080 ;
      LAYER met3 ;
        RECT 1497.825 2802.770 1498.155 2802.785 ;
        RECT 1497.150 2802.470 1498.155 2802.770 ;
        RECT 1497.150 2802.090 1497.450 2802.470 ;
        RECT 1497.825 2802.455 1498.155 2802.470 ;
        RECT 1497.825 2802.090 1498.155 2802.105 ;
        RECT 1497.150 2801.790 1498.155 2802.090 ;
        RECT 1497.825 2801.775 1498.155 2801.790 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2887.950 323.580 2888.270 323.640 ;
        RECT 2901.750 323.580 2902.070 323.640 ;
        RECT 2887.950 323.440 2902.070 323.580 ;
        RECT 2887.950 323.380 2888.270 323.440 ;
        RECT 2901.750 323.380 2902.070 323.440 ;
      LAYER via ;
        RECT 2887.980 323.380 2888.240 323.640 ;
        RECT 2901.780 323.380 2902.040 323.640 ;
      LAYER met2 ;
        RECT 794.970 2740.555 795.250 2740.925 ;
        RECT 2887.970 2740.555 2888.250 2740.925 ;
        RECT 795.040 2731.680 795.180 2740.555 ;
        RECT 794.990 2722.680 795.550 2731.680 ;
        RECT 2888.040 323.670 2888.180 2740.555 ;
        RECT 2887.980 323.350 2888.240 323.670 ;
        RECT 2901.780 323.350 2902.040 323.670 ;
        RECT 2901.840 322.845 2901.980 323.350 ;
        RECT 2901.770 322.475 2902.050 322.845 ;
      LAYER via2 ;
        RECT 794.970 2740.600 795.250 2740.880 ;
        RECT 2887.970 2740.600 2888.250 2740.880 ;
        RECT 2901.770 322.520 2902.050 322.800 ;
      LAYER met3 ;
        RECT 794.945 2740.890 795.275 2740.905 ;
        RECT 2887.945 2740.890 2888.275 2740.905 ;
        RECT 794.945 2740.590 2888.275 2740.890 ;
        RECT 794.945 2740.575 795.275 2740.590 ;
        RECT 2887.945 2740.575 2888.275 2740.590 ;
        RECT 2901.745 322.810 2902.075 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2901.745 322.510 2924.800 322.810 ;
        RECT 2901.745 322.495 2902.075 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 2750.840 1179.830 2750.900 ;
        RECT 1531.870 2750.840 1532.190 2750.900 ;
        RECT 1179.510 2750.700 1532.190 2750.840 ;
        RECT 1179.510 2750.640 1179.830 2750.700 ;
        RECT 1531.870 2750.640 1532.190 2750.700 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 2750.640 1179.800 2750.900 ;
        RECT 1531.900 2750.640 1532.160 2750.900 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 2750.930 1179.740 3498.270 ;
        RECT 1179.540 2750.610 1179.800 2750.930 ;
        RECT 1531.900 2750.610 1532.160 2750.930 ;
        RECT 1531.960 2731.680 1532.100 2750.610 ;
        RECT 1531.910 2722.680 1532.470 2731.680 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 1566.370 3501.220 1566.690 3501.280 ;
        RECT 851.530 3501.080 1566.690 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 1566.370 3501.020 1566.690 3501.080 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 1566.400 3501.020 1566.660 3501.280 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 1566.400 3500.990 1566.660 3501.310 ;
        RECT 1566.460 2731.970 1566.600 3500.990 ;
        RECT 1566.460 2731.830 1569.360 2731.970 ;
        RECT 1569.220 2731.290 1569.360 2731.830 ;
        RECT 1571.010 2731.290 1571.570 2731.680 ;
        RECT 1569.220 2731.150 1571.570 2731.290 ;
        RECT 1571.010 2722.680 1571.570 2731.150 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.600 527.550 3503.660 ;
        RECT 1607.770 3503.600 1608.090 3503.660 ;
        RECT 527.230 3503.460 1608.090 3503.600 ;
        RECT 527.230 3503.400 527.550 3503.460 ;
        RECT 1607.770 3503.400 1608.090 3503.460 ;
      LAYER via ;
        RECT 527.260 3503.400 527.520 3503.660 ;
        RECT 1607.800 3503.400 1608.060 3503.660 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.690 527.460 3517.600 ;
        RECT 527.260 3503.370 527.520 3503.690 ;
        RECT 1607.800 3503.370 1608.060 3503.690 ;
        RECT 1607.860 2731.290 1608.000 3503.370 ;
        RECT 1609.650 2731.290 1610.210 2731.680 ;
        RECT 1607.860 2731.150 1610.210 2731.290 ;
        RECT 1609.650 2722.680 1610.210 2731.150 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 1642.270 3501.900 1642.590 3501.960 ;
        RECT 202.470 3501.760 1642.590 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 1642.270 3501.700 1642.590 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 1642.300 3501.700 1642.560 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 1642.300 3501.670 1642.560 3501.990 ;
        RECT 1642.360 2731.970 1642.500 3501.670 ;
        RECT 1642.360 2731.830 1646.640 2731.970 ;
        RECT 1646.500 2731.290 1646.640 2731.830 ;
        RECT 1648.290 2731.290 1648.850 2731.680 ;
        RECT 1646.500 2731.150 1648.850 2731.290 ;
        RECT 1648.290 2722.680 1648.850 2731.150 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1683.670 3408.740 1683.990 3408.800 ;
        RECT 17.550 3408.600 1683.990 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1683.670 3408.540 1683.990 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1683.700 3408.540 1683.960 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1683.700 3408.510 1683.960 3408.830 ;
        RECT 1683.760 2730.610 1683.900 3408.510 ;
        RECT 1687.390 2730.610 1687.950 2731.680 ;
        RECT 1683.760 2730.470 1687.950 2730.610 ;
        RECT 1687.390 2722.680 1687.950 2730.470 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 1725.070 3119.060 1725.390 3119.120 ;
        RECT 17.090 3118.920 1725.390 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 1725.070 3118.860 1725.390 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 1725.100 3118.860 1725.360 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 1725.100 3118.830 1725.360 3119.150 ;
        RECT 1725.160 2731.290 1725.300 3118.830 ;
        RECT 1726.030 2731.290 1726.590 2731.680 ;
        RECT 1725.160 2731.150 1726.590 2731.290 ;
        RECT 1726.030 2722.680 1726.590 2731.150 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 1759.570 2836.180 1759.890 2836.240 ;
        RECT 17.090 2836.040 1759.890 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 1759.570 2835.980 1759.890 2836.040 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 1759.600 2835.980 1759.860 2836.240 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 1759.600 2835.950 1759.860 2836.270 ;
        RECT 1759.660 2731.970 1759.800 2835.950 ;
        RECT 1759.660 2731.830 1761.640 2731.970 ;
        RECT 1761.500 2731.290 1761.640 2731.830 ;
        RECT 1764.670 2731.290 1765.230 2731.680 ;
        RECT 1761.500 2731.150 1765.230 2731.290 ;
        RECT 1764.670 2722.680 1765.230 2731.150 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 2723.300 32.590 2723.360 ;
        RECT 1802.350 2723.300 1802.670 2723.360 ;
        RECT 32.270 2723.160 1802.670 2723.300 ;
        RECT 32.270 2723.100 32.590 2723.160 ;
        RECT 1802.350 2723.100 1802.670 2723.160 ;
        RECT 14.790 2549.900 15.110 2549.960 ;
        RECT 32.270 2549.900 32.590 2549.960 ;
        RECT 14.790 2549.760 32.590 2549.900 ;
        RECT 14.790 2549.700 15.110 2549.760 ;
        RECT 32.270 2549.700 32.590 2549.760 ;
      LAYER via ;
        RECT 32.300 2723.100 32.560 2723.360 ;
        RECT 1802.380 2723.100 1802.640 2723.360 ;
        RECT 14.820 2549.700 15.080 2549.960 ;
        RECT 32.300 2549.700 32.560 2549.960 ;
      LAYER met2 ;
        RECT 32.300 2723.070 32.560 2723.390 ;
        RECT 1802.380 2723.130 1802.640 2723.390 ;
        RECT 1803.770 2723.130 1804.330 2731.680 ;
        RECT 1802.380 2723.070 1804.330 2723.130 ;
        RECT 32.360 2549.990 32.500 2723.070 ;
        RECT 1802.440 2722.990 1804.330 2723.070 ;
        RECT 1803.770 2722.680 1804.330 2722.990 ;
        RECT 14.820 2549.845 15.080 2549.990 ;
        RECT 14.810 2549.475 15.090 2549.845 ;
        RECT 32.300 2549.670 32.560 2549.990 ;
      LAYER via2 ;
        RECT 14.810 2549.520 15.090 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 14.785 2549.810 15.115 2549.825 ;
        RECT -4.800 2549.510 15.115 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 14.785 2549.495 15.115 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 2744.040 15.570 2744.100 ;
        RECT 1842.370 2744.040 1842.690 2744.100 ;
        RECT 15.250 2743.900 1842.690 2744.040 ;
        RECT 15.250 2743.840 15.570 2743.900 ;
        RECT 1842.370 2743.840 1842.690 2743.900 ;
      LAYER via ;
        RECT 15.280 2743.840 15.540 2744.100 ;
        RECT 1842.400 2743.840 1842.660 2744.100 ;
      LAYER met2 ;
        RECT 15.280 2743.810 15.540 2744.130 ;
        RECT 1842.400 2743.810 1842.660 2744.130 ;
        RECT 15.340 2262.205 15.480 2743.810 ;
        RECT 1842.460 2731.680 1842.600 2743.810 ;
        RECT 1842.410 2722.680 1842.970 2731.680 ;
        RECT 15.270 2261.835 15.550 2262.205 ;
      LAYER via2 ;
        RECT 15.270 2261.880 15.550 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.245 2262.170 15.575 2262.185 ;
        RECT -4.800 2261.870 15.575 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 15.245 2261.855 15.575 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 2743.360 16.030 2743.420 ;
        RECT 1881.010 2743.360 1881.330 2743.420 ;
        RECT 15.710 2743.220 1881.330 2743.360 ;
        RECT 15.710 2743.160 16.030 2743.220 ;
        RECT 1881.010 2743.160 1881.330 2743.220 ;
      LAYER via ;
        RECT 15.740 2743.160 16.000 2743.420 ;
        RECT 1881.040 2743.160 1881.300 2743.420 ;
      LAYER met2 ;
        RECT 15.740 2743.130 16.000 2743.450 ;
        RECT 1881.040 2743.130 1881.300 2743.450 ;
        RECT 15.800 1975.245 15.940 2743.130 ;
        RECT 1881.100 2731.680 1881.240 2743.130 ;
        RECT 1881.050 2722.680 1881.610 2731.680 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2888.870 558.860 2889.190 558.920 ;
        RECT 2903.130 558.860 2903.450 558.920 ;
        RECT 2888.870 558.720 2903.450 558.860 ;
        RECT 2888.870 558.660 2889.190 558.720 ;
        RECT 2903.130 558.660 2903.450 558.720 ;
      LAYER via ;
        RECT 2888.900 558.660 2889.160 558.920 ;
        RECT 2903.160 558.660 2903.420 558.920 ;
      LAYER met2 ;
        RECT 833.610 2741.915 833.890 2742.285 ;
        RECT 2888.890 2741.915 2889.170 2742.285 ;
        RECT 833.680 2731.680 833.820 2741.915 ;
        RECT 833.630 2722.680 834.190 2731.680 ;
        RECT 2888.960 558.950 2889.100 2741.915 ;
        RECT 2888.900 558.630 2889.160 558.950 ;
        RECT 2903.160 558.630 2903.420 558.950 ;
        RECT 2903.220 557.445 2903.360 558.630 ;
        RECT 2903.150 557.075 2903.430 557.445 ;
      LAYER via2 ;
        RECT 833.610 2741.960 833.890 2742.240 ;
        RECT 2888.890 2741.960 2889.170 2742.240 ;
        RECT 2903.150 557.120 2903.430 557.400 ;
      LAYER met3 ;
        RECT 833.585 2742.250 833.915 2742.265 ;
        RECT 2888.865 2742.250 2889.195 2742.265 ;
        RECT 833.585 2741.950 2889.195 2742.250 ;
        RECT 833.585 2741.935 833.915 2741.950 ;
        RECT 2888.865 2741.935 2889.195 2741.950 ;
        RECT 2903.125 557.410 2903.455 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2903.125 557.110 2924.800 557.410 ;
        RECT 2903.125 557.095 2903.455 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2742.340 16.490 2742.400 ;
        RECT 1920.110 2742.340 1920.430 2742.400 ;
        RECT 16.170 2742.200 1920.430 2742.340 ;
        RECT 16.170 2742.140 16.490 2742.200 ;
        RECT 1920.110 2742.140 1920.430 2742.200 ;
      LAYER via ;
        RECT 16.200 2742.140 16.460 2742.400 ;
        RECT 1920.140 2742.140 1920.400 2742.400 ;
      LAYER met2 ;
        RECT 16.200 2742.110 16.460 2742.430 ;
        RECT 1920.140 2742.110 1920.400 2742.430 ;
        RECT 16.260 1687.605 16.400 2742.110 ;
        RECT 1920.200 2731.680 1920.340 2742.110 ;
        RECT 1920.150 2722.680 1920.710 2731.680 ;
        RECT 16.190 1687.235 16.470 1687.605 ;
      LAYER via2 ;
        RECT 16.190 1687.280 16.470 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.165 1687.570 16.495 1687.585 ;
        RECT -4.800 1687.270 16.495 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.165 1687.255 16.495 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2741.660 20.630 2741.720 ;
        RECT 1958.750 2741.660 1959.070 2741.720 ;
        RECT 20.310 2741.520 1959.070 2741.660 ;
        RECT 20.310 2741.460 20.630 2741.520 ;
        RECT 1958.750 2741.460 1959.070 2741.520 ;
      LAYER via ;
        RECT 20.340 2741.460 20.600 2741.720 ;
        RECT 1958.780 2741.460 1959.040 2741.720 ;
      LAYER met2 ;
        RECT 20.340 2741.430 20.600 2741.750 ;
        RECT 1958.780 2741.430 1959.040 2741.750 ;
        RECT 20.400 1472.045 20.540 2741.430 ;
        RECT 1958.840 2731.680 1958.980 2741.430 ;
        RECT 1958.790 2722.680 1959.350 2731.680 ;
        RECT 20.330 1471.675 20.610 1472.045 ;
      LAYER via2 ;
        RECT 20.330 1471.720 20.610 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 20.305 1472.010 20.635 1472.025 ;
        RECT -4.800 1471.710 20.635 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 20.305 1471.695 20.635 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 2740.300 20.170 2740.360 ;
        RECT 1997.390 2740.300 1997.710 2740.360 ;
        RECT 19.850 2740.160 1997.710 2740.300 ;
        RECT 19.850 2740.100 20.170 2740.160 ;
        RECT 1997.390 2740.100 1997.710 2740.160 ;
      LAYER via ;
        RECT 19.880 2740.100 20.140 2740.360 ;
        RECT 1997.420 2740.100 1997.680 2740.360 ;
      LAYER met2 ;
        RECT 19.880 2740.070 20.140 2740.390 ;
        RECT 1997.420 2740.070 1997.680 2740.390 ;
        RECT 19.940 1256.485 20.080 2740.070 ;
        RECT 1997.480 2731.680 1997.620 2740.070 ;
        RECT 1997.430 2722.680 1997.990 2731.680 ;
        RECT 19.870 1256.115 20.150 1256.485 ;
      LAYER via2 ;
        RECT 19.870 1256.160 20.150 1256.440 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 19.845 1256.450 20.175 1256.465 ;
        RECT -4.800 1256.150 20.175 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 19.845 1256.135 20.175 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.510 2743.955 2036.790 2744.325 ;
        RECT 2036.580 2731.680 2036.720 2743.955 ;
        RECT 2036.530 2722.680 2037.090 2731.680 ;
        RECT 763.690 1075.915 763.970 1076.285 ;
        RECT 763.760 1041.605 763.900 1075.915 ;
        RECT 763.690 1041.235 763.970 1041.605 ;
      LAYER via2 ;
        RECT 2036.510 2744.000 2036.790 2744.280 ;
        RECT 763.690 1075.960 763.970 1076.240 ;
        RECT 763.690 1041.280 763.970 1041.560 ;
      LAYER met3 ;
        RECT 763.870 2744.290 764.250 2744.300 ;
        RECT 2036.485 2744.290 2036.815 2744.305 ;
        RECT 763.870 2743.990 2036.815 2744.290 ;
        RECT 763.870 2743.980 764.250 2743.990 ;
        RECT 2036.485 2743.975 2036.815 2743.990 ;
        RECT 763.665 1076.260 763.995 1076.265 ;
        RECT 763.665 1076.250 764.250 1076.260 ;
        RECT 763.440 1075.950 764.250 1076.250 ;
        RECT 763.665 1075.940 764.250 1075.950 ;
        RECT 763.665 1075.935 763.995 1075.940 ;
        RECT 763.665 1041.570 763.995 1041.585 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 3.070 1041.270 763.995 1041.570 ;
        RECT 3.070 1040.890 3.370 1041.270 ;
        RECT 763.665 1041.255 763.995 1041.270 ;
        RECT -4.800 1040.590 3.370 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
      LAYER via3 ;
        RECT 763.900 2743.980 764.220 2744.300 ;
        RECT 763.900 1075.940 764.220 1076.260 ;
      LAYER met4 ;
        RECT 763.895 2743.975 764.225 2744.305 ;
        RECT 763.910 2698.050 764.210 2743.975 ;
        RECT 762.070 2697.750 764.210 2698.050 ;
        RECT 762.070 1219.050 762.370 2697.750 ;
        RECT 762.070 1218.750 764.210 1219.050 ;
        RECT 763.910 1076.265 764.210 1218.750 ;
        RECT 763.895 1075.935 764.225 1076.265 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2075.150 2742.595 2075.430 2742.965 ;
        RECT 2075.220 2731.680 2075.360 2742.595 ;
        RECT 2075.170 2722.680 2075.730 2731.680 ;
        RECT 760.010 1006.555 760.290 1006.925 ;
        RECT 760.080 983.125 760.220 1006.555 ;
        RECT 760.010 982.755 760.290 983.125 ;
      LAYER via2 ;
        RECT 2075.150 2742.640 2075.430 2742.920 ;
        RECT 760.010 1006.600 760.290 1006.880 ;
        RECT 760.010 982.800 760.290 983.080 ;
      LAYER met3 ;
        RECT 759.270 2742.930 759.650 2742.940 ;
        RECT 2075.125 2742.930 2075.455 2742.945 ;
        RECT 759.270 2742.630 2075.455 2742.930 ;
        RECT 759.270 2742.620 759.650 2742.630 ;
        RECT 2075.125 2742.615 2075.455 2742.630 ;
        RECT 759.270 1732.820 759.650 1733.140 ;
        RECT 759.310 1731.100 759.610 1732.820 ;
        RECT 759.270 1730.780 759.650 1731.100 ;
        RECT 759.270 1676.690 759.650 1676.700 ;
        RECT 759.270 1676.390 761.450 1676.690 ;
        RECT 759.270 1676.380 759.650 1676.390 ;
        RECT 761.150 1676.020 761.450 1676.390 ;
        RECT 761.110 1675.700 761.490 1676.020 ;
        RECT 759.270 1006.890 759.650 1006.900 ;
        RECT 759.985 1006.890 760.315 1006.905 ;
        RECT 759.270 1006.590 760.315 1006.890 ;
        RECT 759.270 1006.580 759.650 1006.590 ;
        RECT 759.985 1006.575 760.315 1006.590 ;
        RECT 759.270 983.090 759.650 983.100 ;
        RECT 759.985 983.090 760.315 983.105 ;
        RECT 759.270 982.790 760.315 983.090 ;
        RECT 759.270 982.780 759.650 982.790 ;
        RECT 759.985 982.775 760.315 982.790 ;
        RECT 759.270 828.050 759.650 828.060 ;
        RECT 3.070 827.750 759.650 828.050 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 3.070 825.330 3.370 827.750 ;
        RECT 759.270 827.740 759.650 827.750 ;
        RECT -4.800 825.030 3.370 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
      LAYER via3 ;
        RECT 759.300 2742.620 759.620 2742.940 ;
        RECT 759.300 1732.820 759.620 1733.140 ;
        RECT 759.300 1730.780 759.620 1731.100 ;
        RECT 759.300 1676.380 759.620 1676.700 ;
        RECT 761.140 1675.700 761.460 1676.020 ;
        RECT 759.300 1006.580 759.620 1006.900 ;
        RECT 759.300 982.780 759.620 983.100 ;
        RECT 759.300 827.740 759.620 828.060 ;
      LAYER met4 ;
        RECT 759.295 2742.615 759.625 2742.945 ;
        RECT 759.310 1733.145 759.610 2742.615 ;
        RECT 759.295 1732.815 759.625 1733.145 ;
        RECT 759.295 1730.775 759.625 1731.105 ;
        RECT 759.310 1676.705 759.610 1730.775 ;
        RECT 759.295 1676.375 759.625 1676.705 ;
        RECT 761.135 1675.695 761.465 1676.025 ;
        RECT 761.150 1635.890 761.450 1675.695 ;
        RECT 759.310 1635.590 761.450 1635.890 ;
        RECT 759.310 1006.905 759.610 1635.590 ;
        RECT 759.295 1006.575 759.625 1006.905 ;
        RECT 759.295 982.775 759.625 983.105 ;
        RECT 759.310 828.065 759.610 982.775 ;
        RECT 759.295 827.735 759.625 828.065 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2112.410 2726.530 2112.690 2726.645 ;
        RECT 2113.810 2726.530 2114.370 2731.680 ;
        RECT 2112.410 2726.390 2114.370 2726.530 ;
        RECT 2112.410 2726.275 2112.690 2726.390 ;
        RECT 2113.810 2722.680 2114.370 2726.390 ;
        RECT 14.810 613.515 15.090 613.885 ;
        RECT 14.880 610.485 15.020 613.515 ;
        RECT 14.810 610.115 15.090 610.485 ;
      LAYER via2 ;
        RECT 2112.410 2726.320 2112.690 2726.600 ;
        RECT 14.810 613.560 15.090 613.840 ;
        RECT 14.810 610.160 15.090 610.440 ;
      LAYER met3 ;
        RECT 761.110 2726.610 761.490 2726.620 ;
        RECT 2112.385 2726.610 2112.715 2726.625 ;
        RECT 761.110 2726.310 2112.715 2726.610 ;
        RECT 761.110 2726.300 761.490 2726.310 ;
        RECT 2112.385 2726.295 2112.715 2726.310 ;
        RECT 761.110 2681.050 761.490 2681.060 ;
        RECT 764.790 2681.050 765.170 2681.060 ;
        RECT 761.110 2680.750 765.170 2681.050 ;
        RECT 761.110 2680.740 761.490 2680.750 ;
        RECT 764.790 2680.740 765.170 2680.750 ;
        RECT 764.790 2552.530 765.170 2552.540 ;
        RECT 763.910 2552.230 765.170 2552.530 ;
        RECT 763.910 2550.490 764.210 2552.230 ;
        RECT 764.790 2552.220 765.170 2552.230 ;
        RECT 764.790 2550.490 765.170 2550.500 ;
        RECT 763.910 2550.190 765.170 2550.490 ;
        RECT 764.790 2550.180 765.170 2550.190 ;
        RECT 764.790 1637.620 765.170 1637.940 ;
        RECT 764.830 1635.900 765.130 1637.620 ;
        RECT 764.790 1635.580 765.170 1635.900 ;
        RECT 764.790 1222.140 765.170 1222.460 ;
        RECT 764.830 1221.100 765.130 1222.140 ;
        RECT 764.790 1220.780 765.170 1221.100 ;
        RECT 14.785 613.850 15.115 613.865 ;
        RECT 764.790 613.850 765.170 613.860 ;
        RECT 14.785 613.550 765.170 613.850 ;
        RECT 14.785 613.535 15.115 613.550 ;
        RECT 764.790 613.540 765.170 613.550 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 14.785 610.450 15.115 610.465 ;
        RECT -4.800 610.150 15.115 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 14.785 610.135 15.115 610.150 ;
      LAYER via3 ;
        RECT 761.140 2726.300 761.460 2726.620 ;
        RECT 761.140 2680.740 761.460 2681.060 ;
        RECT 764.820 2680.740 765.140 2681.060 ;
        RECT 764.820 2552.220 765.140 2552.540 ;
        RECT 764.820 2550.180 765.140 2550.500 ;
        RECT 764.820 1637.620 765.140 1637.940 ;
        RECT 764.820 1635.580 765.140 1635.900 ;
        RECT 764.820 1222.140 765.140 1222.460 ;
        RECT 764.820 1220.780 765.140 1221.100 ;
        RECT 764.820 613.540 765.140 613.860 ;
      LAYER met4 ;
        RECT 761.135 2726.295 761.465 2726.625 ;
        RECT 761.150 2681.065 761.450 2726.295 ;
        RECT 761.135 2680.735 761.465 2681.065 ;
        RECT 764.815 2680.735 765.145 2681.065 ;
        RECT 764.830 2552.545 765.130 2680.735 ;
        RECT 764.815 2552.215 765.145 2552.545 ;
        RECT 764.815 2550.175 765.145 2550.505 ;
        RECT 764.830 1637.945 765.130 2550.175 ;
        RECT 764.815 1637.615 765.145 1637.945 ;
        RECT 764.815 1635.575 765.145 1635.905 ;
        RECT 764.830 1222.465 765.130 1635.575 ;
        RECT 764.815 1222.135 765.145 1222.465 ;
        RECT 764.815 1220.775 765.145 1221.105 ;
        RECT 764.830 613.865 765.130 1220.775 ;
        RECT 764.815 613.535 765.145 613.865 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2152.430 2725.850 2152.710 2725.965 ;
        RECT 2152.910 2725.850 2153.470 2731.680 ;
        RECT 2152.430 2725.710 2153.470 2725.850 ;
        RECT 2152.430 2725.595 2152.710 2725.710 ;
        RECT 2152.910 2722.680 2153.470 2725.710 ;
        RECT 16.650 399.995 16.930 400.365 ;
        RECT 16.720 394.925 16.860 399.995 ;
        RECT 16.650 394.555 16.930 394.925 ;
      LAYER via2 ;
        RECT 2152.430 2725.640 2152.710 2725.920 ;
        RECT 16.650 400.040 16.930 400.320 ;
        RECT 16.650 394.600 16.930 394.880 ;
      LAYER met3 ;
        RECT 764.790 2725.930 765.170 2725.940 ;
        RECT 2152.405 2725.930 2152.735 2725.945 ;
        RECT 764.790 2725.630 2152.735 2725.930 ;
        RECT 764.790 2725.620 765.170 2725.630 ;
        RECT 2152.405 2725.615 2152.735 2725.630 ;
        RECT 763.870 2608.290 764.250 2608.300 ;
        RECT 762.990 2607.990 764.250 2608.290 ;
        RECT 762.990 2601.500 763.290 2607.990 ;
        RECT 763.870 2607.980 764.250 2607.990 ;
        RECT 762.950 2601.180 763.330 2601.500 ;
        RECT 760.190 2600.810 760.570 2600.820 ;
        RECT 762.950 2600.810 763.330 2600.820 ;
        RECT 760.190 2600.510 763.330 2600.810 ;
        RECT 760.190 2600.500 760.570 2600.510 ;
        RECT 762.950 2600.500 763.330 2600.510 ;
        RECT 760.190 2553.210 760.570 2553.220 ;
        RECT 763.870 2553.210 764.250 2553.220 ;
        RECT 760.190 2552.910 764.250 2553.210 ;
        RECT 760.190 2552.900 760.570 2552.910 ;
        RECT 763.870 2552.900 764.250 2552.910 ;
        RECT 762.950 2457.330 763.330 2457.340 ;
        RECT 762.950 2457.030 764.210 2457.330 ;
        RECT 762.950 2457.020 763.330 2457.030 ;
        RECT 763.910 2456.660 764.210 2457.030 ;
        RECT 763.870 2456.340 764.250 2456.660 ;
        RECT 763.870 2455.970 764.250 2455.980 ;
        RECT 763.870 2455.670 765.130 2455.970 ;
        RECT 763.870 2455.660 764.250 2455.670 ;
        RECT 760.190 2454.610 760.570 2454.620 ;
        RECT 764.830 2454.610 765.130 2455.670 ;
        RECT 760.190 2454.310 765.130 2454.610 ;
        RECT 760.190 2454.300 760.570 2454.310 ;
        RECT 760.190 2408.370 760.570 2408.380 ;
        RECT 763.870 2408.370 764.250 2408.380 ;
        RECT 760.190 2408.070 764.250 2408.370 ;
        RECT 760.190 2408.060 760.570 2408.070 ;
        RECT 763.870 2408.060 764.250 2408.070 ;
        RECT 761.110 2407.690 761.490 2407.700 ;
        RECT 763.870 2407.690 764.250 2407.700 ;
        RECT 761.110 2407.390 764.250 2407.690 ;
        RECT 761.110 2407.380 761.490 2407.390 ;
        RECT 763.870 2407.380 764.250 2407.390 ;
        RECT 761.110 2360.090 761.490 2360.100 ;
        RECT 763.870 2360.090 764.250 2360.100 ;
        RECT 761.110 2359.790 764.250 2360.090 ;
        RECT 761.110 2359.780 761.490 2359.790 ;
        RECT 763.870 2359.780 764.250 2359.790 ;
        RECT 763.870 2317.930 764.250 2317.940 ;
        RECT 765.710 2317.930 766.090 2317.940 ;
        RECT 763.870 2317.630 766.090 2317.930 ;
        RECT 763.870 2317.620 764.250 2317.630 ;
        RECT 765.710 2317.620 766.090 2317.630 ;
        RECT 763.870 2271.010 764.250 2271.020 ;
        RECT 765.710 2271.010 766.090 2271.020 ;
        RECT 763.870 2270.710 766.090 2271.010 ;
        RECT 763.870 2270.700 764.250 2270.710 ;
        RECT 765.710 2270.700 766.090 2270.710 ;
        RECT 761.110 2262.850 761.490 2262.860 ;
        RECT 763.870 2262.850 764.250 2262.860 ;
        RECT 761.110 2262.550 764.250 2262.850 ;
        RECT 761.110 2262.540 761.490 2262.550 ;
        RECT 763.870 2262.540 764.250 2262.550 ;
        RECT 761.110 2215.930 761.490 2215.940 ;
        RECT 761.110 2215.630 763.290 2215.930 ;
        RECT 761.110 2215.620 761.490 2215.630 ;
        RECT 762.990 2215.260 763.290 2215.630 ;
        RECT 762.950 2214.940 763.330 2215.260 ;
        RECT 761.110 2118.010 761.490 2118.020 ;
        RECT 763.870 2118.010 764.250 2118.020 ;
        RECT 761.110 2117.710 764.250 2118.010 ;
        RECT 761.110 2117.700 761.490 2117.710 ;
        RECT 763.870 2117.700 764.250 2117.710 ;
        RECT 761.110 2071.090 761.490 2071.100 ;
        RECT 761.110 2070.790 764.210 2071.090 ;
        RECT 761.110 2070.780 761.490 2070.790 ;
        RECT 763.910 2070.420 764.210 2070.790 ;
        RECT 763.870 2070.100 764.250 2070.420 ;
        RECT 761.110 2021.450 761.490 2021.460 ;
        RECT 763.870 2021.450 764.250 2021.460 ;
        RECT 761.110 2021.150 764.250 2021.450 ;
        RECT 761.110 2021.140 761.490 2021.150 ;
        RECT 763.870 2021.140 764.250 2021.150 ;
        RECT 761.110 1974.530 761.490 1974.540 ;
        RECT 761.110 1974.230 764.210 1974.530 ;
        RECT 761.110 1974.220 761.490 1974.230 ;
        RECT 763.910 1973.860 764.210 1974.230 ;
        RECT 763.870 1973.540 764.250 1973.860 ;
        RECT 761.110 1828.330 761.490 1828.340 ;
        RECT 763.870 1828.330 764.250 1828.340 ;
        RECT 761.110 1828.030 764.250 1828.330 ;
        RECT 761.110 1828.020 761.490 1828.030 ;
        RECT 763.870 1828.020 764.250 1828.030 ;
        RECT 761.110 1781.410 761.490 1781.420 ;
        RECT 761.110 1781.110 764.210 1781.410 ;
        RECT 761.110 1781.100 761.490 1781.110 ;
        RECT 763.910 1780.740 764.210 1781.110 ;
        RECT 763.870 1780.420 764.250 1780.740 ;
        RECT 763.870 1637.620 764.250 1637.940 ;
        RECT 763.910 1635.900 764.210 1637.620 ;
        RECT 763.870 1635.580 764.250 1635.900 ;
        RECT 761.110 1635.210 761.490 1635.220 ;
        RECT 763.870 1635.210 764.250 1635.220 ;
        RECT 761.110 1634.910 764.250 1635.210 ;
        RECT 761.110 1634.900 761.490 1634.910 ;
        RECT 763.870 1634.900 764.250 1634.910 ;
        RECT 761.110 1588.290 761.490 1588.300 ;
        RECT 761.110 1587.990 764.210 1588.290 ;
        RECT 761.110 1587.980 761.490 1587.990 ;
        RECT 763.910 1587.620 764.210 1587.990 ;
        RECT 763.870 1587.300 764.250 1587.620 ;
        RECT 761.110 1538.650 761.490 1538.660 ;
        RECT 763.870 1538.650 764.250 1538.660 ;
        RECT 761.110 1538.350 764.250 1538.650 ;
        RECT 761.110 1538.340 761.490 1538.350 ;
        RECT 763.870 1538.340 764.250 1538.350 ;
        RECT 761.110 1491.730 761.490 1491.740 ;
        RECT 761.110 1491.430 764.210 1491.730 ;
        RECT 761.110 1491.420 761.490 1491.430 ;
        RECT 763.910 1491.060 764.210 1491.430 ;
        RECT 763.870 1490.740 764.250 1491.060 ;
        RECT 761.110 1442.090 761.490 1442.100 ;
        RECT 763.870 1442.090 764.250 1442.100 ;
        RECT 761.110 1441.790 764.250 1442.090 ;
        RECT 761.110 1441.780 761.490 1441.790 ;
        RECT 763.870 1441.780 764.250 1441.790 ;
        RECT 761.110 1395.170 761.490 1395.180 ;
        RECT 761.110 1394.870 764.210 1395.170 ;
        RECT 761.110 1394.860 761.490 1394.870 ;
        RECT 763.910 1394.500 764.210 1394.870 ;
        RECT 763.870 1394.180 764.250 1394.500 ;
        RECT 763.870 1296.940 764.250 1297.260 ;
        RECT 762.950 1296.570 763.330 1296.580 ;
        RECT 763.910 1296.570 764.210 1296.940 ;
        RECT 762.950 1296.270 764.210 1296.570 ;
        RECT 762.950 1296.260 763.330 1296.270 ;
        RECT 762.950 1242.540 763.330 1242.860 ;
        RECT 762.990 1242.170 763.290 1242.540 ;
        RECT 763.870 1242.170 764.250 1242.180 ;
        RECT 762.990 1241.870 764.250 1242.170 ;
        RECT 763.870 1241.860 764.250 1241.870 ;
        RECT 763.870 1241.490 764.250 1241.500 ;
        RECT 767.550 1241.490 767.930 1241.500 ;
        RECT 763.870 1241.190 767.930 1241.490 ;
        RECT 763.870 1241.180 764.250 1241.190 ;
        RECT 767.550 1241.180 767.930 1241.190 ;
        RECT 765.710 1193.890 766.090 1193.900 ;
        RECT 767.550 1193.890 767.930 1193.900 ;
        RECT 765.710 1193.590 767.930 1193.890 ;
        RECT 765.710 1193.580 766.090 1193.590 ;
        RECT 767.550 1193.580 767.930 1193.590 ;
        RECT 765.710 1111.300 766.090 1111.620 ;
        RECT 765.750 1110.250 766.050 1111.300 ;
        RECT 766.630 1110.250 767.010 1110.260 ;
        RECT 765.750 1109.950 767.010 1110.250 ;
        RECT 766.630 1109.940 767.010 1109.950 ;
        RECT 763.870 1075.570 764.250 1075.580 ;
        RECT 765.710 1075.570 766.090 1075.580 ;
        RECT 763.870 1075.270 766.090 1075.570 ;
        RECT 763.870 1075.260 764.250 1075.270 ;
        RECT 765.710 1075.260 766.090 1075.270 ;
        RECT 16.625 400.330 16.955 400.345 ;
        RECT 763.870 400.330 764.250 400.340 ;
        RECT 16.625 400.030 764.250 400.330 ;
        RECT 16.625 400.015 16.955 400.030 ;
        RECT 763.870 400.020 764.250 400.030 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.625 394.890 16.955 394.905 ;
        RECT -4.800 394.590 16.955 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.625 394.575 16.955 394.590 ;
      LAYER via3 ;
        RECT 764.820 2725.620 765.140 2725.940 ;
        RECT 763.900 2607.980 764.220 2608.300 ;
        RECT 762.980 2601.180 763.300 2601.500 ;
        RECT 760.220 2600.500 760.540 2600.820 ;
        RECT 762.980 2600.500 763.300 2600.820 ;
        RECT 760.220 2552.900 760.540 2553.220 ;
        RECT 763.900 2552.900 764.220 2553.220 ;
        RECT 762.980 2457.020 763.300 2457.340 ;
        RECT 763.900 2456.340 764.220 2456.660 ;
        RECT 763.900 2455.660 764.220 2455.980 ;
        RECT 760.220 2454.300 760.540 2454.620 ;
        RECT 760.220 2408.060 760.540 2408.380 ;
        RECT 763.900 2408.060 764.220 2408.380 ;
        RECT 761.140 2407.380 761.460 2407.700 ;
        RECT 763.900 2407.380 764.220 2407.700 ;
        RECT 761.140 2359.780 761.460 2360.100 ;
        RECT 763.900 2359.780 764.220 2360.100 ;
        RECT 763.900 2317.620 764.220 2317.940 ;
        RECT 765.740 2317.620 766.060 2317.940 ;
        RECT 763.900 2270.700 764.220 2271.020 ;
        RECT 765.740 2270.700 766.060 2271.020 ;
        RECT 761.140 2262.540 761.460 2262.860 ;
        RECT 763.900 2262.540 764.220 2262.860 ;
        RECT 761.140 2215.620 761.460 2215.940 ;
        RECT 762.980 2214.940 763.300 2215.260 ;
        RECT 761.140 2117.700 761.460 2118.020 ;
        RECT 763.900 2117.700 764.220 2118.020 ;
        RECT 761.140 2070.780 761.460 2071.100 ;
        RECT 763.900 2070.100 764.220 2070.420 ;
        RECT 761.140 2021.140 761.460 2021.460 ;
        RECT 763.900 2021.140 764.220 2021.460 ;
        RECT 761.140 1974.220 761.460 1974.540 ;
        RECT 763.900 1973.540 764.220 1973.860 ;
        RECT 761.140 1828.020 761.460 1828.340 ;
        RECT 763.900 1828.020 764.220 1828.340 ;
        RECT 761.140 1781.100 761.460 1781.420 ;
        RECT 763.900 1780.420 764.220 1780.740 ;
        RECT 763.900 1637.620 764.220 1637.940 ;
        RECT 763.900 1635.580 764.220 1635.900 ;
        RECT 761.140 1634.900 761.460 1635.220 ;
        RECT 763.900 1634.900 764.220 1635.220 ;
        RECT 761.140 1587.980 761.460 1588.300 ;
        RECT 763.900 1587.300 764.220 1587.620 ;
        RECT 761.140 1538.340 761.460 1538.660 ;
        RECT 763.900 1538.340 764.220 1538.660 ;
        RECT 761.140 1491.420 761.460 1491.740 ;
        RECT 763.900 1490.740 764.220 1491.060 ;
        RECT 761.140 1441.780 761.460 1442.100 ;
        RECT 763.900 1441.780 764.220 1442.100 ;
        RECT 761.140 1394.860 761.460 1395.180 ;
        RECT 763.900 1394.180 764.220 1394.500 ;
        RECT 763.900 1296.940 764.220 1297.260 ;
        RECT 762.980 1296.260 763.300 1296.580 ;
        RECT 762.980 1242.540 763.300 1242.860 ;
        RECT 763.900 1241.860 764.220 1242.180 ;
        RECT 763.900 1241.180 764.220 1241.500 ;
        RECT 767.580 1241.180 767.900 1241.500 ;
        RECT 765.740 1193.580 766.060 1193.900 ;
        RECT 767.580 1193.580 767.900 1193.900 ;
        RECT 765.740 1111.300 766.060 1111.620 ;
        RECT 766.660 1109.940 766.980 1110.260 ;
        RECT 763.900 1075.260 764.220 1075.580 ;
        RECT 765.740 1075.260 766.060 1075.580 ;
        RECT 763.900 400.020 764.220 400.340 ;
      LAYER met4 ;
        RECT 764.815 2725.615 765.145 2725.945 ;
        RECT 764.830 2687.850 765.130 2725.615 ;
        RECT 762.990 2687.550 765.130 2687.850 ;
        RECT 762.990 2657.250 763.290 2687.550 ;
        RECT 762.990 2656.950 764.210 2657.250 ;
        RECT 763.910 2608.305 764.210 2656.950 ;
        RECT 763.895 2607.975 764.225 2608.305 ;
        RECT 762.975 2601.175 763.305 2601.505 ;
        RECT 762.990 2600.825 763.290 2601.175 ;
        RECT 760.215 2600.495 760.545 2600.825 ;
        RECT 762.975 2600.495 763.305 2600.825 ;
        RECT 760.230 2553.225 760.530 2600.495 ;
        RECT 760.215 2552.895 760.545 2553.225 ;
        RECT 763.895 2552.895 764.225 2553.225 ;
        RECT 763.910 2504.250 764.210 2552.895 ;
        RECT 762.990 2503.950 764.210 2504.250 ;
        RECT 762.990 2457.345 763.290 2503.950 ;
        RECT 762.975 2457.015 763.305 2457.345 ;
        RECT 763.895 2456.335 764.225 2456.665 ;
        RECT 763.910 2455.985 764.210 2456.335 ;
        RECT 763.895 2455.655 764.225 2455.985 ;
        RECT 760.215 2454.295 760.545 2454.625 ;
        RECT 760.230 2408.385 760.530 2454.295 ;
        RECT 760.215 2408.055 760.545 2408.385 ;
        RECT 763.895 2408.055 764.225 2408.385 ;
        RECT 763.910 2407.705 764.210 2408.055 ;
        RECT 761.135 2407.375 761.465 2407.705 ;
        RECT 763.895 2407.375 764.225 2407.705 ;
        RECT 761.150 2360.105 761.450 2407.375 ;
        RECT 761.135 2359.775 761.465 2360.105 ;
        RECT 763.895 2359.775 764.225 2360.105 ;
        RECT 763.910 2317.945 764.210 2359.775 ;
        RECT 763.895 2317.615 764.225 2317.945 ;
        RECT 765.735 2317.615 766.065 2317.945 ;
        RECT 765.750 2271.025 766.050 2317.615 ;
        RECT 763.895 2270.695 764.225 2271.025 ;
        RECT 765.735 2270.695 766.065 2271.025 ;
        RECT 763.910 2262.865 764.210 2270.695 ;
        RECT 761.135 2262.535 761.465 2262.865 ;
        RECT 763.895 2262.535 764.225 2262.865 ;
        RECT 761.150 2215.945 761.450 2262.535 ;
        RECT 761.135 2215.615 761.465 2215.945 ;
        RECT 762.975 2215.250 763.305 2215.265 ;
        RECT 762.975 2214.950 764.210 2215.250 ;
        RECT 762.975 2214.935 763.305 2214.950 ;
        RECT 763.910 2118.025 764.210 2214.950 ;
        RECT 761.135 2117.695 761.465 2118.025 ;
        RECT 763.895 2117.695 764.225 2118.025 ;
        RECT 761.150 2071.105 761.450 2117.695 ;
        RECT 761.135 2070.775 761.465 2071.105 ;
        RECT 763.895 2070.095 764.225 2070.425 ;
        RECT 763.910 2021.465 764.210 2070.095 ;
        RECT 761.135 2021.135 761.465 2021.465 ;
        RECT 763.895 2021.135 764.225 2021.465 ;
        RECT 761.150 1974.545 761.450 2021.135 ;
        RECT 761.135 1974.215 761.465 1974.545 ;
        RECT 763.895 1973.535 764.225 1973.865 ;
        RECT 763.910 1828.345 764.210 1973.535 ;
        RECT 761.135 1828.015 761.465 1828.345 ;
        RECT 763.895 1828.015 764.225 1828.345 ;
        RECT 761.150 1781.425 761.450 1828.015 ;
        RECT 761.135 1781.095 761.465 1781.425 ;
        RECT 763.895 1780.415 764.225 1780.745 ;
        RECT 763.910 1637.945 764.210 1780.415 ;
        RECT 763.895 1637.615 764.225 1637.945 ;
        RECT 763.895 1635.575 764.225 1635.905 ;
        RECT 763.910 1635.225 764.210 1635.575 ;
        RECT 761.135 1634.895 761.465 1635.225 ;
        RECT 763.895 1634.895 764.225 1635.225 ;
        RECT 761.150 1588.305 761.450 1634.895 ;
        RECT 761.135 1587.975 761.465 1588.305 ;
        RECT 763.895 1587.295 764.225 1587.625 ;
        RECT 763.910 1538.665 764.210 1587.295 ;
        RECT 761.135 1538.335 761.465 1538.665 ;
        RECT 763.895 1538.335 764.225 1538.665 ;
        RECT 761.150 1491.745 761.450 1538.335 ;
        RECT 761.135 1491.415 761.465 1491.745 ;
        RECT 763.895 1490.735 764.225 1491.065 ;
        RECT 763.910 1442.105 764.210 1490.735 ;
        RECT 761.135 1441.775 761.465 1442.105 ;
        RECT 763.895 1441.775 764.225 1442.105 ;
        RECT 761.150 1395.185 761.450 1441.775 ;
        RECT 761.135 1394.855 761.465 1395.185 ;
        RECT 763.895 1394.175 764.225 1394.505 ;
        RECT 763.910 1297.265 764.210 1394.175 ;
        RECT 763.895 1296.935 764.225 1297.265 ;
        RECT 762.975 1296.255 763.305 1296.585 ;
        RECT 762.990 1242.865 763.290 1296.255 ;
        RECT 762.975 1242.535 763.305 1242.865 ;
        RECT 763.895 1241.855 764.225 1242.185 ;
        RECT 763.910 1241.505 764.210 1241.855 ;
        RECT 763.895 1241.175 764.225 1241.505 ;
        RECT 767.575 1241.175 767.905 1241.505 ;
        RECT 767.590 1193.905 767.890 1241.175 ;
        RECT 765.735 1193.575 766.065 1193.905 ;
        RECT 767.575 1193.575 767.905 1193.905 ;
        RECT 765.750 1111.625 766.050 1193.575 ;
        RECT 765.735 1111.295 766.065 1111.625 ;
        RECT 766.655 1109.935 766.985 1110.265 ;
        RECT 766.670 1103.450 766.970 1109.935 ;
        RECT 765.750 1103.150 766.970 1103.450 ;
        RECT 765.750 1075.585 766.050 1103.150 ;
        RECT 763.895 1075.255 764.225 1075.585 ;
        RECT 765.735 1075.255 766.065 1075.585 ;
        RECT 763.910 400.345 764.210 1075.255 ;
        RECT 763.895 400.015 764.225 400.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2191.125 2718.385 2191.295 2723.315 ;
        RECT 62.245 2713.965 62.415 2714.815 ;
        RECT 96.745 2714.645 96.915 2715.495 ;
        RECT 144.585 2714.305 144.755 2715.495 ;
        RECT 158.845 2713.965 159.015 2714.815 ;
        RECT 193.345 2714.645 193.515 2715.495 ;
        RECT 241.185 2714.305 241.355 2715.495 ;
        RECT 255.445 2713.965 255.615 2714.815 ;
        RECT 289.945 2714.645 290.115 2715.495 ;
        RECT 337.785 2714.305 337.955 2715.495 ;
        RECT 352.045 2713.965 352.215 2714.815 ;
        RECT 386.545 2714.645 386.715 2715.495 ;
        RECT 434.385 2714.305 434.555 2715.495 ;
        RECT 448.645 2713.965 448.815 2714.815 ;
        RECT 483.145 2714.645 483.315 2715.495 ;
        RECT 530.985 2714.305 531.155 2715.495 ;
        RECT 545.245 2713.965 545.415 2714.815 ;
        RECT 579.745 2714.645 579.915 2715.495 ;
        RECT 627.585 2714.305 627.755 2715.495 ;
        RECT 724.645 2714.985 724.815 2715.835 ;
        RECT 641.845 2713.965 642.015 2714.815 ;
        RECT 689.685 2714.645 690.315 2714.815 ;
        RECT 772.485 2714.305 772.655 2715.835 ;
        RECT 773.405 2714.475 773.575 2714.815 ;
        RECT 821.245 2714.645 821.415 2716.175 ;
        RECT 772.945 2714.305 773.575 2714.475 ;
        RECT 844.705 2714.305 844.875 2716.175 ;
        RECT 882.425 2714.305 882.595 2715.835 ;
        RECT 917.385 2714.645 917.555 2715.835 ;
        RECT 917.845 2714.645 918.015 2716.175 ;
        RECT 941.305 2714.305 941.475 2716.175 ;
        RECT 966.605 2714.305 966.775 2715.835 ;
        RECT 1013.985 2714.645 1014.155 2715.835 ;
        RECT 1014.445 2714.645 1014.615 2716.175 ;
        RECT 1037.905 2714.305 1038.075 2716.175 ;
        RECT 1055.845 2714.305 1056.015 2715.835 ;
        RECT 1103.685 2714.645 1103.855 2715.835 ;
        RECT 1249.045 2715.325 1249.215 2716.175 ;
        RECT 1296.885 2714.985 1297.055 2716.175 ;
        RECT 1325.865 2714.305 1326.035 2715.155 ;
        RECT 1365.425 2714.305 1365.595 2715.835 ;
        RECT 1400.385 2714.645 1400.555 2715.835 ;
        RECT 1400.845 2714.645 1401.015 2716.175 ;
        RECT 1424.305 2714.305 1424.475 2716.175 ;
        RECT 1462.025 2714.305 1462.195 2715.835 ;
        RECT 1496.985 2714.645 1497.155 2715.835 ;
        RECT 1558.625 2714.305 1558.795 2715.835 ;
        RECT 1593.585 2714.645 1593.755 2715.835 ;
        RECT 1594.045 2714.645 1594.215 2716.175 ;
        RECT 1617.505 2714.305 1617.675 2716.175 ;
        RECT 1635.445 2714.305 1635.615 2715.495 ;
        RECT 2124.885 2715.325 2125.055 2716.175 ;
        RECT 1848.885 2714.985 1850.435 2715.155 ;
        RECT 1945.485 2714.985 1946.115 2715.155 ;
        RECT 1993.785 2714.985 1994.875 2715.155 ;
        RECT 1848.885 2714.305 1849.055 2714.985 ;
      LAYER mcon ;
        RECT 2191.125 2723.145 2191.295 2723.315 ;
        RECT 821.245 2716.005 821.415 2716.175 ;
        RECT 724.645 2715.665 724.815 2715.835 ;
        RECT 96.745 2715.325 96.915 2715.495 ;
        RECT 62.245 2714.645 62.415 2714.815 ;
        RECT 144.585 2715.325 144.755 2715.495 ;
        RECT 193.345 2715.325 193.515 2715.495 ;
        RECT 158.845 2714.645 159.015 2714.815 ;
        RECT 241.185 2715.325 241.355 2715.495 ;
        RECT 289.945 2715.325 290.115 2715.495 ;
        RECT 255.445 2714.645 255.615 2714.815 ;
        RECT 337.785 2715.325 337.955 2715.495 ;
        RECT 386.545 2715.325 386.715 2715.495 ;
        RECT 352.045 2714.645 352.215 2714.815 ;
        RECT 434.385 2715.325 434.555 2715.495 ;
        RECT 483.145 2715.325 483.315 2715.495 ;
        RECT 448.645 2714.645 448.815 2714.815 ;
        RECT 530.985 2715.325 531.155 2715.495 ;
        RECT 579.745 2715.325 579.915 2715.495 ;
        RECT 545.245 2714.645 545.415 2714.815 ;
        RECT 627.585 2715.325 627.755 2715.495 ;
        RECT 772.485 2715.665 772.655 2715.835 ;
        RECT 641.845 2714.645 642.015 2714.815 ;
        RECT 690.145 2714.645 690.315 2714.815 ;
        RECT 773.405 2714.645 773.575 2714.815 ;
        RECT 844.705 2716.005 844.875 2716.175 ;
        RECT 917.845 2716.005 918.015 2716.175 ;
        RECT 882.425 2715.665 882.595 2715.835 ;
        RECT 917.385 2715.665 917.555 2715.835 ;
        RECT 941.305 2716.005 941.475 2716.175 ;
        RECT 1014.445 2716.005 1014.615 2716.175 ;
        RECT 966.605 2715.665 966.775 2715.835 ;
        RECT 1013.985 2715.665 1014.155 2715.835 ;
        RECT 1037.905 2716.005 1038.075 2716.175 ;
        RECT 1249.045 2716.005 1249.215 2716.175 ;
        RECT 1055.845 2715.665 1056.015 2715.835 ;
        RECT 1103.685 2715.665 1103.855 2715.835 ;
        RECT 1296.885 2716.005 1297.055 2716.175 ;
        RECT 1400.845 2716.005 1401.015 2716.175 ;
        RECT 1365.425 2715.665 1365.595 2715.835 ;
        RECT 1325.865 2714.985 1326.035 2715.155 ;
        RECT 1400.385 2715.665 1400.555 2715.835 ;
        RECT 1424.305 2716.005 1424.475 2716.175 ;
        RECT 1594.045 2716.005 1594.215 2716.175 ;
        RECT 1462.025 2715.665 1462.195 2715.835 ;
        RECT 1496.985 2715.665 1497.155 2715.835 ;
        RECT 1558.625 2715.665 1558.795 2715.835 ;
        RECT 1593.585 2715.665 1593.755 2715.835 ;
        RECT 1617.505 2716.005 1617.675 2716.175 ;
        RECT 2124.885 2716.005 2125.055 2716.175 ;
        RECT 1635.445 2715.325 1635.615 2715.495 ;
        RECT 1850.265 2714.985 1850.435 2715.155 ;
        RECT 1945.945 2714.985 1946.115 2715.155 ;
        RECT 1994.705 2714.985 1994.875 2715.155 ;
      LAYER met1 ;
        RECT 2191.050 2723.300 2191.370 2723.360 ;
        RECT 2190.855 2723.160 2191.370 2723.300 ;
        RECT 2191.050 2723.100 2191.370 2723.160 ;
        RECT 2191.065 2718.540 2191.355 2718.585 ;
        RECT 2187.000 2718.400 2191.355 2718.540 ;
        RECT 821.185 2716.160 821.475 2716.205 ;
        RECT 844.645 2716.160 844.935 2716.205 ;
        RECT 821.185 2716.020 844.935 2716.160 ;
        RECT 821.185 2715.975 821.475 2716.020 ;
        RECT 844.645 2715.975 844.935 2716.020 ;
        RECT 917.785 2716.160 918.075 2716.205 ;
        RECT 941.245 2716.160 941.535 2716.205 ;
        RECT 917.785 2716.020 941.535 2716.160 ;
        RECT 917.785 2715.975 918.075 2716.020 ;
        RECT 941.245 2715.975 941.535 2716.020 ;
        RECT 1014.385 2716.160 1014.675 2716.205 ;
        RECT 1037.845 2716.160 1038.135 2716.205 ;
        RECT 1014.385 2716.020 1038.135 2716.160 ;
        RECT 1014.385 2715.975 1014.675 2716.020 ;
        RECT 1037.845 2715.975 1038.135 2716.020 ;
        RECT 1248.985 2716.160 1249.275 2716.205 ;
        RECT 1296.825 2716.160 1297.115 2716.205 ;
        RECT 1248.985 2716.020 1297.115 2716.160 ;
        RECT 1248.985 2715.975 1249.275 2716.020 ;
        RECT 1296.825 2715.975 1297.115 2716.020 ;
        RECT 1400.785 2716.160 1401.075 2716.205 ;
        RECT 1424.245 2716.160 1424.535 2716.205 ;
        RECT 1400.785 2716.020 1424.535 2716.160 ;
        RECT 1400.785 2715.975 1401.075 2716.020 ;
        RECT 1424.245 2715.975 1424.535 2716.020 ;
        RECT 1593.985 2716.160 1594.275 2716.205 ;
        RECT 1617.445 2716.160 1617.735 2716.205 ;
        RECT 2124.825 2716.160 2125.115 2716.205 ;
        RECT 1593.985 2716.020 1617.735 2716.160 ;
        RECT 1593.985 2715.975 1594.275 2716.020 ;
        RECT 1617.445 2715.975 1617.735 2716.020 ;
        RECT 2089.940 2716.020 2125.115 2716.160 ;
        RECT 724.585 2715.820 724.875 2715.865 ;
        RECT 772.425 2715.820 772.715 2715.865 ;
        RECT 724.585 2715.680 772.715 2715.820 ;
        RECT 724.585 2715.635 724.875 2715.680 ;
        RECT 772.425 2715.635 772.715 2715.680 ;
        RECT 882.365 2715.820 882.655 2715.865 ;
        RECT 917.325 2715.820 917.615 2715.865 ;
        RECT 882.365 2715.680 917.615 2715.820 ;
        RECT 882.365 2715.635 882.655 2715.680 ;
        RECT 917.325 2715.635 917.615 2715.680 ;
        RECT 966.545 2715.820 966.835 2715.865 ;
        RECT 1013.925 2715.820 1014.215 2715.865 ;
        RECT 966.545 2715.680 1014.215 2715.820 ;
        RECT 966.545 2715.635 966.835 2715.680 ;
        RECT 1013.925 2715.635 1014.215 2715.680 ;
        RECT 1055.785 2715.820 1056.075 2715.865 ;
        RECT 1103.625 2715.820 1103.915 2715.865 ;
        RECT 1055.785 2715.680 1103.915 2715.820 ;
        RECT 1055.785 2715.635 1056.075 2715.680 ;
        RECT 1103.625 2715.635 1103.915 2715.680 ;
        RECT 1365.365 2715.820 1365.655 2715.865 ;
        RECT 1400.325 2715.820 1400.615 2715.865 ;
        RECT 1365.365 2715.680 1400.615 2715.820 ;
        RECT 1365.365 2715.635 1365.655 2715.680 ;
        RECT 1400.325 2715.635 1400.615 2715.680 ;
        RECT 1461.965 2715.820 1462.255 2715.865 ;
        RECT 1496.925 2715.820 1497.215 2715.865 ;
        RECT 1461.965 2715.680 1497.215 2715.820 ;
        RECT 1461.965 2715.635 1462.255 2715.680 ;
        RECT 1496.925 2715.635 1497.215 2715.680 ;
        RECT 1558.565 2715.820 1558.855 2715.865 ;
        RECT 1593.525 2715.820 1593.815 2715.865 ;
        RECT 1558.565 2715.680 1593.815 2715.820 ;
        RECT 1558.565 2715.635 1558.855 2715.680 ;
        RECT 1593.525 2715.635 1593.815 2715.680 ;
        RECT 96.685 2715.480 96.975 2715.525 ;
        RECT 144.525 2715.480 144.815 2715.525 ;
        RECT 96.685 2715.340 144.815 2715.480 ;
        RECT 96.685 2715.295 96.975 2715.340 ;
        RECT 144.525 2715.295 144.815 2715.340 ;
        RECT 193.285 2715.480 193.575 2715.525 ;
        RECT 241.125 2715.480 241.415 2715.525 ;
        RECT 193.285 2715.340 241.415 2715.480 ;
        RECT 193.285 2715.295 193.575 2715.340 ;
        RECT 241.125 2715.295 241.415 2715.340 ;
        RECT 289.885 2715.480 290.175 2715.525 ;
        RECT 337.725 2715.480 338.015 2715.525 ;
        RECT 289.885 2715.340 338.015 2715.480 ;
        RECT 289.885 2715.295 290.175 2715.340 ;
        RECT 337.725 2715.295 338.015 2715.340 ;
        RECT 386.485 2715.480 386.775 2715.525 ;
        RECT 434.325 2715.480 434.615 2715.525 ;
        RECT 386.485 2715.340 434.615 2715.480 ;
        RECT 386.485 2715.295 386.775 2715.340 ;
        RECT 434.325 2715.295 434.615 2715.340 ;
        RECT 483.085 2715.480 483.375 2715.525 ;
        RECT 530.925 2715.480 531.215 2715.525 ;
        RECT 483.085 2715.340 531.215 2715.480 ;
        RECT 483.085 2715.295 483.375 2715.340 ;
        RECT 530.925 2715.295 531.215 2715.340 ;
        RECT 579.685 2715.480 579.975 2715.525 ;
        RECT 627.525 2715.480 627.815 2715.525 ;
        RECT 1248.985 2715.480 1249.275 2715.525 ;
        RECT 579.685 2715.340 627.815 2715.480 ;
        RECT 579.685 2715.295 579.975 2715.340 ;
        RECT 627.525 2715.295 627.815 2715.340 ;
        RECT 1172.240 2715.340 1249.275 2715.480 ;
        RECT 724.585 2715.140 724.875 2715.185 ;
        RECT 691.080 2715.000 724.875 2715.140 ;
        RECT 62.185 2714.800 62.475 2714.845 ;
        RECT 96.685 2714.800 96.975 2714.845 ;
        RECT 62.185 2714.660 96.975 2714.800 ;
        RECT 62.185 2714.615 62.475 2714.660 ;
        RECT 96.685 2714.615 96.975 2714.660 ;
        RECT 158.785 2714.800 159.075 2714.845 ;
        RECT 193.285 2714.800 193.575 2714.845 ;
        RECT 158.785 2714.660 193.575 2714.800 ;
        RECT 158.785 2714.615 159.075 2714.660 ;
        RECT 193.285 2714.615 193.575 2714.660 ;
        RECT 255.385 2714.800 255.675 2714.845 ;
        RECT 289.885 2714.800 290.175 2714.845 ;
        RECT 255.385 2714.660 290.175 2714.800 ;
        RECT 255.385 2714.615 255.675 2714.660 ;
        RECT 289.885 2714.615 290.175 2714.660 ;
        RECT 351.985 2714.800 352.275 2714.845 ;
        RECT 386.485 2714.800 386.775 2714.845 ;
        RECT 351.985 2714.660 386.775 2714.800 ;
        RECT 351.985 2714.615 352.275 2714.660 ;
        RECT 386.485 2714.615 386.775 2714.660 ;
        RECT 448.585 2714.800 448.875 2714.845 ;
        RECT 483.085 2714.800 483.375 2714.845 ;
        RECT 448.585 2714.660 483.375 2714.800 ;
        RECT 448.585 2714.615 448.875 2714.660 ;
        RECT 483.085 2714.615 483.375 2714.660 ;
        RECT 545.185 2714.800 545.475 2714.845 ;
        RECT 579.685 2714.800 579.975 2714.845 ;
        RECT 545.185 2714.660 579.975 2714.800 ;
        RECT 545.185 2714.615 545.475 2714.660 ;
        RECT 579.685 2714.615 579.975 2714.660 ;
        RECT 641.785 2714.800 642.075 2714.845 ;
        RECT 689.625 2714.800 689.915 2714.845 ;
        RECT 641.785 2714.660 689.915 2714.800 ;
        RECT 641.785 2714.615 642.075 2714.660 ;
        RECT 689.625 2714.615 689.915 2714.660 ;
        RECT 690.085 2714.800 690.375 2714.845 ;
        RECT 691.080 2714.800 691.220 2715.000 ;
        RECT 724.585 2714.955 724.875 2715.000 ;
        RECT 690.085 2714.660 691.220 2714.800 ;
        RECT 773.345 2714.800 773.635 2714.845 ;
        RECT 821.185 2714.800 821.475 2714.845 ;
        RECT 773.345 2714.660 821.475 2714.800 ;
        RECT 690.085 2714.615 690.375 2714.660 ;
        RECT 773.345 2714.615 773.635 2714.660 ;
        RECT 821.185 2714.615 821.475 2714.660 ;
        RECT 917.325 2714.800 917.615 2714.845 ;
        RECT 917.785 2714.800 918.075 2714.845 ;
        RECT 917.325 2714.660 918.075 2714.800 ;
        RECT 917.325 2714.615 917.615 2714.660 ;
        RECT 917.785 2714.615 918.075 2714.660 ;
        RECT 1013.925 2714.800 1014.215 2714.845 ;
        RECT 1014.385 2714.800 1014.675 2714.845 ;
        RECT 1013.925 2714.660 1014.675 2714.800 ;
        RECT 1013.925 2714.615 1014.215 2714.660 ;
        RECT 1014.385 2714.615 1014.675 2714.660 ;
        RECT 1103.625 2714.800 1103.915 2714.845 ;
        RECT 1172.240 2714.800 1172.380 2715.340 ;
        RECT 1248.985 2715.295 1249.275 2715.340 ;
        RECT 1635.385 2715.480 1635.675 2715.525 ;
        RECT 2089.940 2715.480 2090.080 2716.020 ;
        RECT 2124.825 2715.975 2125.115 2716.020 ;
        RECT 2187.000 2715.820 2187.140 2718.400 ;
        RECT 2191.065 2718.355 2191.355 2718.400 ;
        RECT 2139.160 2715.680 2187.140 2715.820 ;
        RECT 1635.385 2715.340 1683.440 2715.480 ;
        RECT 1635.385 2715.295 1635.675 2715.340 ;
        RECT 1296.825 2715.140 1297.115 2715.185 ;
        RECT 1325.805 2715.140 1326.095 2715.185 ;
        RECT 1296.825 2715.000 1326.095 2715.140 ;
        RECT 1296.825 2714.955 1297.115 2715.000 ;
        RECT 1325.805 2714.955 1326.095 2715.000 ;
        RECT 1497.460 2715.000 1521.060 2715.140 ;
        RECT 1103.625 2714.660 1172.380 2714.800 ;
        RECT 1400.325 2714.800 1400.615 2714.845 ;
        RECT 1400.785 2714.800 1401.075 2714.845 ;
        RECT 1400.325 2714.660 1401.075 2714.800 ;
        RECT 1103.625 2714.615 1103.915 2714.660 ;
        RECT 1400.325 2714.615 1400.615 2714.660 ;
        RECT 1400.785 2714.615 1401.075 2714.660 ;
        RECT 1496.925 2714.800 1497.215 2714.845 ;
        RECT 1497.460 2714.800 1497.600 2715.000 ;
        RECT 1496.925 2714.660 1497.600 2714.800 ;
        RECT 1496.925 2714.615 1497.215 2714.660 ;
        RECT 144.525 2714.460 144.815 2714.505 ;
        RECT 241.125 2714.460 241.415 2714.505 ;
        RECT 337.725 2714.460 338.015 2714.505 ;
        RECT 434.325 2714.460 434.615 2714.505 ;
        RECT 530.925 2714.460 531.215 2714.505 ;
        RECT 627.525 2714.460 627.815 2714.505 ;
        RECT 772.425 2714.460 772.715 2714.505 ;
        RECT 772.885 2714.460 773.175 2714.505 ;
        RECT 144.525 2714.320 158.540 2714.460 ;
        RECT 144.525 2714.275 144.815 2714.320 ;
        RECT 17.550 2714.120 17.870 2714.180 ;
        RECT 62.185 2714.120 62.475 2714.165 ;
        RECT 17.550 2713.980 62.475 2714.120 ;
        RECT 158.400 2714.120 158.540 2714.320 ;
        RECT 241.125 2714.320 255.140 2714.460 ;
        RECT 241.125 2714.275 241.415 2714.320 ;
        RECT 158.785 2714.120 159.075 2714.165 ;
        RECT 158.400 2713.980 159.075 2714.120 ;
        RECT 255.000 2714.120 255.140 2714.320 ;
        RECT 337.725 2714.320 351.740 2714.460 ;
        RECT 337.725 2714.275 338.015 2714.320 ;
        RECT 255.385 2714.120 255.675 2714.165 ;
        RECT 255.000 2713.980 255.675 2714.120 ;
        RECT 351.600 2714.120 351.740 2714.320 ;
        RECT 434.325 2714.320 448.340 2714.460 ;
        RECT 434.325 2714.275 434.615 2714.320 ;
        RECT 351.985 2714.120 352.275 2714.165 ;
        RECT 351.600 2713.980 352.275 2714.120 ;
        RECT 448.200 2714.120 448.340 2714.320 ;
        RECT 530.925 2714.320 544.940 2714.460 ;
        RECT 530.925 2714.275 531.215 2714.320 ;
        RECT 448.585 2714.120 448.875 2714.165 ;
        RECT 448.200 2713.980 448.875 2714.120 ;
        RECT 544.800 2714.120 544.940 2714.320 ;
        RECT 627.525 2714.320 641.540 2714.460 ;
        RECT 627.525 2714.275 627.815 2714.320 ;
        RECT 545.185 2714.120 545.475 2714.165 ;
        RECT 544.800 2713.980 545.475 2714.120 ;
        RECT 641.400 2714.120 641.540 2714.320 ;
        RECT 772.425 2714.320 773.175 2714.460 ;
        RECT 772.425 2714.275 772.715 2714.320 ;
        RECT 772.885 2714.275 773.175 2714.320 ;
        RECT 844.645 2714.275 844.935 2714.505 ;
        RECT 882.365 2714.275 882.655 2714.505 ;
        RECT 941.245 2714.275 941.535 2714.505 ;
        RECT 966.545 2714.275 966.835 2714.505 ;
        RECT 1037.845 2714.275 1038.135 2714.505 ;
        RECT 1055.785 2714.275 1056.075 2714.505 ;
        RECT 1325.805 2714.275 1326.095 2714.505 ;
        RECT 1365.365 2714.275 1365.655 2714.505 ;
        RECT 1424.245 2714.275 1424.535 2714.505 ;
        RECT 1461.965 2714.275 1462.255 2714.505 ;
        RECT 641.785 2714.120 642.075 2714.165 ;
        RECT 641.400 2713.980 642.075 2714.120 ;
        RECT 844.720 2714.120 844.860 2714.275 ;
        RECT 882.440 2714.120 882.580 2714.275 ;
        RECT 844.720 2713.980 882.580 2714.120 ;
        RECT 941.320 2714.120 941.460 2714.275 ;
        RECT 966.620 2714.120 966.760 2714.275 ;
        RECT 941.320 2713.980 966.760 2714.120 ;
        RECT 1037.920 2714.120 1038.060 2714.275 ;
        RECT 1055.860 2714.120 1056.000 2714.275 ;
        RECT 1037.920 2713.980 1056.000 2714.120 ;
        RECT 1325.880 2714.120 1326.020 2714.275 ;
        RECT 1365.440 2714.120 1365.580 2714.275 ;
        RECT 1325.880 2713.980 1365.580 2714.120 ;
        RECT 1424.320 2714.120 1424.460 2714.275 ;
        RECT 1462.040 2714.120 1462.180 2714.275 ;
        RECT 1424.320 2713.980 1462.180 2714.120 ;
        RECT 1520.920 2714.120 1521.060 2715.000 ;
        RECT 1593.525 2714.800 1593.815 2714.845 ;
        RECT 1593.985 2714.800 1594.275 2714.845 ;
        RECT 1593.525 2714.660 1594.275 2714.800 ;
        RECT 1683.300 2714.800 1683.440 2715.340 ;
        RECT 1732.520 2715.340 1779.580 2715.480 ;
        RECT 1732.520 2714.800 1732.660 2715.340 ;
        RECT 1683.300 2714.660 1732.660 2714.800 ;
        RECT 1593.525 2714.615 1593.815 2714.660 ;
        RECT 1593.985 2714.615 1594.275 2714.660 ;
        RECT 1558.565 2714.275 1558.855 2714.505 ;
        RECT 1617.445 2714.275 1617.735 2714.505 ;
        RECT 1635.385 2714.275 1635.675 2714.505 ;
        RECT 1558.640 2714.120 1558.780 2714.275 ;
        RECT 1520.920 2713.980 1558.780 2714.120 ;
        RECT 1617.520 2714.120 1617.660 2714.275 ;
        RECT 1635.460 2714.120 1635.600 2714.275 ;
        RECT 1617.520 2713.980 1635.600 2714.120 ;
        RECT 1779.440 2714.120 1779.580 2715.340 ;
        RECT 2043.480 2715.340 2090.080 2715.480 ;
        RECT 2124.825 2715.480 2125.115 2715.525 ;
        RECT 2139.160 2715.480 2139.300 2715.680 ;
        RECT 2124.825 2715.340 2139.300 2715.480 ;
        RECT 1850.205 2715.140 1850.495 2715.185 ;
        RECT 1945.425 2715.140 1945.715 2715.185 ;
        RECT 1850.205 2715.000 1945.715 2715.140 ;
        RECT 1850.205 2714.955 1850.495 2715.000 ;
        RECT 1945.425 2714.955 1945.715 2715.000 ;
        RECT 1945.885 2715.140 1946.175 2715.185 ;
        RECT 1993.725 2715.140 1994.015 2715.185 ;
        RECT 1945.885 2715.000 1994.015 2715.140 ;
        RECT 1945.885 2714.955 1946.175 2715.000 ;
        RECT 1993.725 2714.955 1994.015 2715.000 ;
        RECT 1994.645 2715.140 1994.935 2715.185 ;
        RECT 2043.480 2715.140 2043.620 2715.340 ;
        RECT 2124.825 2715.295 2125.115 2715.340 ;
        RECT 1994.645 2715.000 2004.520 2715.140 ;
        RECT 1994.645 2714.955 1994.935 2715.000 ;
        RECT 2004.380 2714.800 2004.520 2715.000 ;
        RECT 2042.560 2715.000 2043.620 2715.140 ;
        RECT 2042.560 2714.800 2042.700 2715.000 ;
        RECT 2004.380 2714.660 2042.700 2714.800 ;
        RECT 1848.825 2714.460 1849.115 2714.505 ;
        RECT 1848.440 2714.320 1849.115 2714.460 ;
        RECT 1848.440 2714.120 1848.580 2714.320 ;
        RECT 1848.825 2714.275 1849.115 2714.320 ;
        RECT 1779.440 2713.980 1848.580 2714.120 ;
        RECT 17.550 2713.920 17.870 2713.980 ;
        RECT 62.185 2713.935 62.475 2713.980 ;
        RECT 158.785 2713.935 159.075 2713.980 ;
        RECT 255.385 2713.935 255.675 2713.980 ;
        RECT 351.985 2713.935 352.275 2713.980 ;
        RECT 448.585 2713.935 448.875 2713.980 ;
        RECT 545.185 2713.935 545.475 2713.980 ;
        RECT 641.785 2713.935 642.075 2713.980 ;
      LAYER via ;
        RECT 2191.080 2723.100 2191.340 2723.360 ;
        RECT 17.580 2713.920 17.840 2714.180 ;
      LAYER met2 ;
        RECT 2191.080 2723.130 2191.340 2723.390 ;
        RECT 2191.550 2723.130 2192.110 2731.680 ;
        RECT 2191.080 2723.070 2192.110 2723.130 ;
        RECT 2191.140 2722.990 2192.110 2723.070 ;
        RECT 2191.550 2722.680 2192.110 2722.990 ;
        RECT 17.580 2713.890 17.840 2714.210 ;
        RECT 17.640 179.365 17.780 2713.890 ;
        RECT 17.570 178.995 17.850 179.365 ;
      LAYER via2 ;
        RECT 17.570 179.040 17.850 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.545 179.330 17.875 179.345 ;
        RECT -4.800 179.030 17.875 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.545 179.015 17.875 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 874.605 2721.445 874.775 2723.655 ;
      LAYER mcon ;
        RECT 874.605 2723.485 874.775 2723.655 ;
      LAYER met1 ;
        RECT 874.530 2723.640 874.850 2723.700 ;
        RECT 874.335 2723.500 874.850 2723.640 ;
        RECT 874.530 2723.440 874.850 2723.500 ;
        RECT 874.545 2721.600 874.835 2721.645 ;
        RECT 2889.790 2721.600 2890.110 2721.660 ;
        RECT 874.545 2721.460 2890.110 2721.600 ;
        RECT 874.545 2721.415 874.835 2721.460 ;
        RECT 2889.790 2721.400 2890.110 2721.460 ;
        RECT 2889.790 793.460 2890.110 793.520 ;
        RECT 2900.370 793.460 2900.690 793.520 ;
        RECT 2889.790 793.320 2900.690 793.460 ;
        RECT 2889.790 793.260 2890.110 793.320 ;
        RECT 2900.370 793.260 2900.690 793.320 ;
      LAYER via ;
        RECT 874.560 2723.440 874.820 2723.700 ;
        RECT 2889.820 2721.400 2890.080 2721.660 ;
        RECT 2889.820 793.260 2890.080 793.520 ;
        RECT 2900.400 793.260 2900.660 793.520 ;
      LAYER met2 ;
        RECT 872.730 2723.810 873.290 2731.680 ;
        RECT 872.730 2723.730 874.760 2723.810 ;
        RECT 872.730 2723.670 874.820 2723.730 ;
        RECT 872.730 2722.680 873.290 2723.670 ;
        RECT 874.560 2723.410 874.820 2723.670 ;
        RECT 2889.820 2721.370 2890.080 2721.690 ;
        RECT 2889.880 793.550 2890.020 2721.370 ;
        RECT 2889.820 793.230 2890.080 793.550 ;
        RECT 2900.400 793.230 2900.660 793.550 ;
        RECT 2900.460 792.045 2900.600 793.230 ;
        RECT 2900.390 791.675 2900.670 792.045 ;
      LAYER via2 ;
        RECT 2900.390 791.720 2900.670 792.000 ;
      LAYER met3 ;
        RECT 2900.365 792.010 2900.695 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.365 791.710 2924.800 792.010 ;
        RECT 2900.365 791.695 2900.695 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 913.245 2722.125 913.415 2723.655 ;
      LAYER mcon ;
        RECT 913.245 2723.485 913.415 2723.655 ;
      LAYER met1 ;
        RECT 913.170 2723.640 913.490 2723.700 ;
        RECT 912.975 2723.500 913.490 2723.640 ;
        RECT 913.170 2723.440 913.490 2723.500 ;
        RECT 913.185 2722.280 913.475 2722.325 ;
        RECT 2890.250 2722.280 2890.570 2722.340 ;
        RECT 913.185 2722.140 2890.570 2722.280 ;
        RECT 913.185 2722.095 913.475 2722.140 ;
        RECT 2890.250 2722.080 2890.570 2722.140 ;
        RECT 2890.250 1028.060 2890.570 1028.120 ;
        RECT 2904.050 1028.060 2904.370 1028.120 ;
        RECT 2890.250 1027.920 2904.370 1028.060 ;
        RECT 2890.250 1027.860 2890.570 1027.920 ;
        RECT 2904.050 1027.860 2904.370 1027.920 ;
      LAYER via ;
        RECT 913.200 2723.440 913.460 2723.700 ;
        RECT 2890.280 2722.080 2890.540 2722.340 ;
        RECT 2890.280 1027.860 2890.540 1028.120 ;
        RECT 2904.080 1027.860 2904.340 1028.120 ;
      LAYER met2 ;
        RECT 911.370 2723.810 911.930 2731.680 ;
        RECT 911.370 2723.730 913.400 2723.810 ;
        RECT 911.370 2723.670 913.460 2723.730 ;
        RECT 911.370 2722.680 911.930 2723.670 ;
        RECT 913.200 2723.410 913.460 2723.670 ;
        RECT 2890.280 2722.050 2890.540 2722.370 ;
        RECT 2890.340 1028.150 2890.480 2722.050 ;
        RECT 2890.280 1027.830 2890.540 1028.150 ;
        RECT 2904.080 1027.830 2904.340 1028.150 ;
        RECT 2904.140 1026.645 2904.280 1027.830 ;
        RECT 2904.070 1026.275 2904.350 1026.645 ;
      LAYER via2 ;
        RECT 2904.070 1026.320 2904.350 1026.600 ;
      LAYER met3 ;
        RECT 2904.045 1026.610 2904.375 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2904.045 1026.310 2924.800 1026.610 ;
        RECT 2904.045 1026.295 2904.375 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.990 2743.275 950.270 2743.645 ;
        RECT 950.060 2731.680 950.200 2743.275 ;
        RECT 950.010 2722.680 950.570 2731.680 ;
      LAYER via2 ;
        RECT 949.990 2743.320 950.270 2743.600 ;
      LAYER met3 ;
        RECT 949.965 2743.610 950.295 2743.625 ;
        RECT 2232.190 2743.610 2232.570 2743.620 ;
        RECT 949.965 2743.310 2232.570 2743.610 ;
        RECT 949.965 2743.295 950.295 2743.310 ;
        RECT 2232.190 2743.300 2232.570 2743.310 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2916.710 1260.910 2924.800 1261.210 ;
        RECT 2234.030 1257.810 2234.410 1257.820 ;
        RECT 2234.030 1257.510 2256.450 1257.810 ;
        RECT 2234.030 1257.500 2234.410 1257.510 ;
        RECT 2256.150 1257.130 2256.450 1257.510 ;
        RECT 2304.910 1257.510 2353.050 1257.810 ;
        RECT 2256.150 1256.830 2304.290 1257.130 ;
        RECT 2303.990 1256.450 2304.290 1256.830 ;
        RECT 2304.910 1256.450 2305.210 1257.510 ;
        RECT 2352.750 1257.130 2353.050 1257.510 ;
        RECT 2401.510 1257.510 2449.650 1257.810 ;
        RECT 2352.750 1256.830 2400.890 1257.130 ;
        RECT 2303.990 1256.150 2305.210 1256.450 ;
        RECT 2400.590 1256.450 2400.890 1256.830 ;
        RECT 2401.510 1256.450 2401.810 1257.510 ;
        RECT 2449.350 1257.130 2449.650 1257.510 ;
        RECT 2498.110 1257.510 2546.250 1257.810 ;
        RECT 2449.350 1256.830 2497.490 1257.130 ;
        RECT 2400.590 1256.150 2401.810 1256.450 ;
        RECT 2497.190 1256.450 2497.490 1256.830 ;
        RECT 2498.110 1256.450 2498.410 1257.510 ;
        RECT 2545.950 1257.130 2546.250 1257.510 ;
        RECT 2594.710 1257.510 2642.850 1257.810 ;
        RECT 2545.950 1256.830 2594.090 1257.130 ;
        RECT 2497.190 1256.150 2498.410 1256.450 ;
        RECT 2593.790 1256.450 2594.090 1256.830 ;
        RECT 2594.710 1256.450 2595.010 1257.510 ;
        RECT 2642.550 1257.130 2642.850 1257.510 ;
        RECT 2691.310 1257.510 2739.450 1257.810 ;
        RECT 2642.550 1256.830 2690.690 1257.130 ;
        RECT 2593.790 1256.150 2595.010 1256.450 ;
        RECT 2690.390 1256.450 2690.690 1256.830 ;
        RECT 2691.310 1256.450 2691.610 1257.510 ;
        RECT 2739.150 1257.130 2739.450 1257.510 ;
        RECT 2787.910 1257.510 2836.050 1257.810 ;
        RECT 2739.150 1256.830 2787.290 1257.130 ;
        RECT 2690.390 1256.150 2691.610 1256.450 ;
        RECT 2786.990 1256.450 2787.290 1256.830 ;
        RECT 2787.910 1256.450 2788.210 1257.510 ;
        RECT 2835.750 1257.130 2836.050 1257.510 ;
        RECT 2916.710 1257.130 2917.010 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2835.750 1256.830 2883.890 1257.130 ;
        RECT 2786.990 1256.150 2788.210 1256.450 ;
        RECT 2883.590 1256.450 2883.890 1256.830 ;
        RECT 2884.510 1256.830 2917.010 1257.130 ;
        RECT 2884.510 1256.450 2884.810 1256.830 ;
        RECT 2883.590 1256.150 2884.810 1256.450 ;
      LAYER via3 ;
        RECT 2232.220 2743.300 2232.540 2743.620 ;
        RECT 2234.060 1257.500 2234.380 1257.820 ;
      LAYER met4 ;
        RECT 2232.215 2743.295 2232.545 2743.625 ;
        RECT 2232.230 1273.450 2232.530 2743.295 ;
        RECT 2232.230 1273.150 2234.370 1273.450 ;
        RECT 2234.070 1257.825 2234.370 1273.150 ;
        RECT 2234.055 1257.495 2234.385 1257.825 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.090 2744.635 989.370 2745.005 ;
        RECT 989.160 2731.680 989.300 2744.635 ;
        RECT 989.110 2722.680 989.670 2731.680 ;
      LAYER via2 ;
        RECT 989.090 2744.680 989.370 2744.960 ;
      LAYER met3 ;
        RECT 989.065 2744.970 989.395 2744.985 ;
        RECT 2233.110 2744.970 2233.490 2744.980 ;
        RECT 989.065 2744.670 2233.490 2744.970 ;
        RECT 989.065 2744.655 989.395 2744.670 ;
        RECT 2233.110 2744.660 2233.490 2744.670 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2916.710 1495.510 2924.800 1495.810 ;
        RECT 2233.110 1492.410 2233.490 1492.420 ;
        RECT 2233.110 1492.110 2256.450 1492.410 ;
        RECT 2233.110 1492.100 2233.490 1492.110 ;
        RECT 2256.150 1491.730 2256.450 1492.110 ;
        RECT 2304.910 1492.110 2353.050 1492.410 ;
        RECT 2256.150 1491.430 2304.290 1491.730 ;
        RECT 2303.990 1491.050 2304.290 1491.430 ;
        RECT 2304.910 1491.050 2305.210 1492.110 ;
        RECT 2352.750 1491.730 2353.050 1492.110 ;
        RECT 2401.510 1492.110 2449.650 1492.410 ;
        RECT 2352.750 1491.430 2400.890 1491.730 ;
        RECT 2303.990 1490.750 2305.210 1491.050 ;
        RECT 2400.590 1491.050 2400.890 1491.430 ;
        RECT 2401.510 1491.050 2401.810 1492.110 ;
        RECT 2449.350 1491.730 2449.650 1492.110 ;
        RECT 2498.110 1492.110 2546.250 1492.410 ;
        RECT 2449.350 1491.430 2497.490 1491.730 ;
        RECT 2400.590 1490.750 2401.810 1491.050 ;
        RECT 2497.190 1491.050 2497.490 1491.430 ;
        RECT 2498.110 1491.050 2498.410 1492.110 ;
        RECT 2545.950 1491.730 2546.250 1492.110 ;
        RECT 2594.710 1492.110 2642.850 1492.410 ;
        RECT 2545.950 1491.430 2594.090 1491.730 ;
        RECT 2497.190 1490.750 2498.410 1491.050 ;
        RECT 2593.790 1491.050 2594.090 1491.430 ;
        RECT 2594.710 1491.050 2595.010 1492.110 ;
        RECT 2642.550 1491.730 2642.850 1492.110 ;
        RECT 2691.310 1492.110 2739.450 1492.410 ;
        RECT 2642.550 1491.430 2690.690 1491.730 ;
        RECT 2593.790 1490.750 2595.010 1491.050 ;
        RECT 2690.390 1491.050 2690.690 1491.430 ;
        RECT 2691.310 1491.050 2691.610 1492.110 ;
        RECT 2739.150 1491.730 2739.450 1492.110 ;
        RECT 2787.910 1492.110 2836.050 1492.410 ;
        RECT 2739.150 1491.430 2787.290 1491.730 ;
        RECT 2690.390 1490.750 2691.610 1491.050 ;
        RECT 2786.990 1491.050 2787.290 1491.430 ;
        RECT 2787.910 1491.050 2788.210 1492.110 ;
        RECT 2835.750 1491.730 2836.050 1492.110 ;
        RECT 2916.710 1491.730 2917.010 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2835.750 1491.430 2883.890 1491.730 ;
        RECT 2786.990 1490.750 2788.210 1491.050 ;
        RECT 2883.590 1491.050 2883.890 1491.430 ;
        RECT 2884.510 1491.430 2917.010 1491.730 ;
        RECT 2884.510 1491.050 2884.810 1491.430 ;
        RECT 2883.590 1490.750 2884.810 1491.050 ;
      LAYER via3 ;
        RECT 2233.140 2744.660 2233.460 2744.980 ;
        RECT 2233.140 1492.100 2233.460 1492.420 ;
      LAYER met4 ;
        RECT 2233.135 2744.655 2233.465 2744.985 ;
        RECT 2233.150 1492.425 2233.450 2744.655 ;
        RECT 2233.135 1492.095 2233.465 1492.425 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.270 2723.130 1027.550 2723.245 ;
        RECT 1027.750 2723.130 1028.310 2731.680 ;
        RECT 1027.270 2722.990 1028.310 2723.130 ;
        RECT 1027.270 2722.875 1027.550 2722.990 ;
        RECT 1027.750 2722.680 1028.310 2722.990 ;
        RECT 2900.850 2716.075 2901.130 2716.445 ;
        RECT 2900.920 1730.445 2901.060 2716.075 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
      LAYER via2 ;
        RECT 1027.270 2722.920 1027.550 2723.200 ;
        RECT 2900.850 2716.120 2901.130 2716.400 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
        RECT 1027.245 2723.220 1027.575 2723.225 ;
        RECT 1026.990 2723.210 1027.575 2723.220 ;
        RECT 1026.790 2722.910 1027.575 2723.210 ;
        RECT 1026.990 2722.900 1027.575 2722.910 ;
        RECT 1027.245 2722.895 1027.575 2722.900 ;
        RECT 1134.630 2719.810 1135.010 2719.820 ;
        RECT 1158.550 2719.810 1158.930 2719.820 ;
        RECT 1134.630 2719.510 1158.930 2719.810 ;
        RECT 1134.630 2719.500 1135.010 2719.510 ;
        RECT 1158.550 2719.500 1158.930 2719.510 ;
        RECT 1026.990 2716.410 1027.370 2716.420 ;
        RECT 1134.630 2716.410 1135.010 2716.420 ;
        RECT 1026.990 2716.110 1135.010 2716.410 ;
        RECT 1026.990 2716.100 1027.370 2716.110 ;
        RECT 1134.630 2716.100 1135.010 2716.110 ;
        RECT 1158.550 2716.410 1158.930 2716.420 ;
        RECT 2900.825 2716.410 2901.155 2716.425 ;
        RECT 1158.550 2716.110 2901.155 2716.410 ;
        RECT 1158.550 2716.100 1158.930 2716.110 ;
        RECT 2900.825 2716.095 2901.155 2716.110 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
      LAYER via3 ;
        RECT 1027.020 2722.900 1027.340 2723.220 ;
        RECT 1134.660 2719.500 1134.980 2719.820 ;
        RECT 1158.580 2719.500 1158.900 2719.820 ;
        RECT 1027.020 2716.100 1027.340 2716.420 ;
        RECT 1134.660 2716.100 1134.980 2716.420 ;
        RECT 1158.580 2716.100 1158.900 2716.420 ;
      LAYER met4 ;
        RECT 1027.015 2722.895 1027.345 2723.225 ;
        RECT 1027.030 2716.425 1027.330 2722.895 ;
        RECT 1134.655 2719.495 1134.985 2719.825 ;
        RECT 1158.575 2719.495 1158.905 2719.825 ;
        RECT 1134.670 2716.425 1134.970 2719.495 ;
        RECT 1158.590 2716.425 1158.890 2719.495 ;
        RECT 1027.015 2716.095 1027.345 2716.425 ;
        RECT 1134.655 2716.095 1134.985 2716.425 ;
        RECT 1158.575 2716.095 1158.905 2716.425 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1066.390 2723.130 1066.950 2731.680 ;
        RECT 1067.290 2723.130 1067.570 2723.245 ;
        RECT 1066.390 2722.990 1067.570 2723.130 ;
        RECT 1066.390 2722.680 1066.950 2722.990 ;
        RECT 1067.290 2722.875 1067.570 2722.990 ;
        RECT 2899.010 2717.435 2899.290 2717.805 ;
        RECT 2899.080 1965.045 2899.220 2717.435 ;
        RECT 2899.010 1964.675 2899.290 1965.045 ;
      LAYER via2 ;
        RECT 1067.290 2722.920 1067.570 2723.200 ;
        RECT 2899.010 2717.480 2899.290 2717.760 ;
        RECT 2899.010 1964.720 2899.290 1965.000 ;
      LAYER met3 ;
        RECT 1067.265 2723.220 1067.595 2723.225 ;
        RECT 1067.265 2723.210 1067.850 2723.220 ;
        RECT 1067.265 2722.910 1068.050 2723.210 ;
        RECT 1067.265 2722.900 1067.850 2722.910 ;
        RECT 1067.265 2722.895 1067.595 2722.900 ;
        RECT 1067.470 2717.770 1067.850 2717.780 ;
        RECT 2898.985 2717.770 2899.315 2717.785 ;
        RECT 1067.470 2717.470 2899.315 2717.770 ;
        RECT 1067.470 2717.460 1067.850 2717.470 ;
        RECT 2898.985 2717.455 2899.315 2717.470 ;
        RECT 2898.985 1965.010 2899.315 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.985 1964.710 2924.800 1965.010 ;
        RECT 2898.985 1964.695 2899.315 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
      LAYER via3 ;
        RECT 1067.500 2722.900 1067.820 2723.220 ;
        RECT 1067.500 2717.460 1067.820 2717.780 ;
      LAYER met4 ;
        RECT 1067.495 2722.895 1067.825 2723.225 ;
        RECT 1067.510 2717.785 1067.810 2722.895 ;
        RECT 1067.495 2717.455 1067.825 2717.785 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1105.490 2723.130 1106.050 2731.680 ;
        RECT 1106.390 2723.130 1106.670 2723.245 ;
        RECT 1105.490 2722.990 1106.670 2723.130 ;
        RECT 1105.490 2722.680 1106.050 2722.990 ;
        RECT 1106.390 2722.875 1106.670 2722.990 ;
        RECT 2898.090 2718.115 2898.370 2718.485 ;
        RECT 2898.160 2199.645 2898.300 2718.115 ;
        RECT 2898.090 2199.275 2898.370 2199.645 ;
      LAYER via2 ;
        RECT 1106.390 2722.920 1106.670 2723.200 ;
        RECT 2898.090 2718.160 2898.370 2718.440 ;
        RECT 2898.090 2199.320 2898.370 2199.600 ;
      LAYER met3 ;
        RECT 1106.365 2723.210 1106.695 2723.225 ;
        RECT 1107.030 2723.210 1107.410 2723.220 ;
        RECT 1106.365 2722.910 1107.410 2723.210 ;
        RECT 1106.365 2722.895 1106.695 2722.910 ;
        RECT 1107.030 2722.900 1107.410 2722.910 ;
        RECT 1107.030 2718.450 1107.410 2718.460 ;
        RECT 2898.065 2718.450 2898.395 2718.465 ;
        RECT 1107.030 2718.150 2898.395 2718.450 ;
        RECT 1107.030 2718.140 1107.410 2718.150 ;
        RECT 2898.065 2718.135 2898.395 2718.150 ;
        RECT 2898.065 2199.610 2898.395 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.065 2199.310 2924.800 2199.610 ;
        RECT 2898.065 2199.295 2898.395 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
      LAYER via3 ;
        RECT 1107.060 2722.900 1107.380 2723.220 ;
        RECT 1107.060 2718.140 1107.380 2718.460 ;
      LAYER met4 ;
        RECT 1107.055 2722.895 1107.385 2723.225 ;
        RECT 1107.070 2718.465 1107.370 2722.895 ;
        RECT 1107.055 2718.135 1107.385 2718.465 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1703.450 201.180 1703.770 201.240 ;
        RECT 1704.830 201.180 1705.150 201.240 ;
        RECT 1703.450 201.040 1705.150 201.180 ;
        RECT 1703.450 200.980 1703.770 201.040 ;
        RECT 1704.830 200.980 1705.150 201.040 ;
        RECT 1007.470 200.840 1007.790 200.900 ;
        RECT 1096.710 200.840 1097.030 200.900 ;
        RECT 1007.470 200.700 1097.030 200.840 ;
        RECT 1007.470 200.640 1007.790 200.700 ;
        RECT 1096.710 200.640 1097.030 200.700 ;
        RECT 1606.390 200.840 1606.710 200.900 ;
        RECT 1607.770 200.840 1608.090 200.900 ;
        RECT 1606.390 200.700 1608.090 200.840 ;
        RECT 1606.390 200.640 1606.710 200.700 ;
        RECT 1607.770 200.640 1608.090 200.700 ;
        RECT 1799.590 200.840 1799.910 200.900 ;
        RECT 1800.970 200.840 1801.290 200.900 ;
        RECT 1799.590 200.700 1801.290 200.840 ;
        RECT 1799.590 200.640 1799.910 200.700 ;
        RECT 1800.970 200.640 1801.290 200.700 ;
        RECT 2221.870 200.500 2222.190 200.560 ;
        RECT 2236.130 200.500 2236.450 200.560 ;
        RECT 2221.870 200.360 2236.450 200.500 ;
        RECT 2221.870 200.300 2222.190 200.360 ;
        RECT 2236.130 200.300 2236.450 200.360 ;
        RECT 2380.110 200.500 2380.430 200.560 ;
        RECT 2414.610 200.500 2414.930 200.560 ;
        RECT 2380.110 200.360 2414.930 200.500 ;
        RECT 2380.110 200.300 2380.430 200.360 ;
        RECT 2414.610 200.300 2414.930 200.360 ;
      LAYER via ;
        RECT 1703.480 200.980 1703.740 201.240 ;
        RECT 1704.860 200.980 1705.120 201.240 ;
        RECT 1007.500 200.640 1007.760 200.900 ;
        RECT 1096.740 200.640 1097.000 200.900 ;
        RECT 1606.420 200.640 1606.680 200.900 ;
        RECT 1607.800 200.640 1608.060 200.900 ;
        RECT 1799.620 200.640 1799.880 200.900 ;
        RECT 1801.000 200.640 1801.260 200.900 ;
        RECT 2221.900 200.300 2222.160 200.560 ;
        RECT 2236.160 200.300 2236.420 200.560 ;
        RECT 2380.140 200.300 2380.400 200.560 ;
        RECT 2414.640 200.300 2414.900 200.560 ;
      LAYER met2 ;
        RECT 769.230 2723.130 769.790 2731.680 ;
        RECT 770.130 2723.130 770.410 2723.245 ;
        RECT 769.230 2722.990 770.410 2723.130 ;
        RECT 769.230 2722.680 769.790 2722.990 ;
        RECT 770.130 2722.875 770.410 2722.990 ;
        RECT 1193.330 202.795 1193.610 203.165 ;
        RECT 1200.230 202.795 1200.510 203.165 ;
        RECT 881.910 201.690 882.190 201.805 ;
        RECT 882.830 201.690 883.110 201.805 ;
        RECT 881.910 201.550 883.110 201.690 ;
        RECT 881.910 201.435 882.190 201.550 ;
        RECT 882.830 201.435 883.110 201.550 ;
        RECT 1145.030 201.435 1145.310 201.805 ;
        RECT 1007.490 200.755 1007.770 201.125 ;
        RECT 1007.500 200.610 1007.760 200.755 ;
        RECT 1096.740 200.610 1097.000 200.930 ;
        RECT 1096.800 200.445 1096.940 200.610 ;
        RECT 1096.730 200.075 1097.010 200.445 ;
        RECT 1145.100 199.085 1145.240 201.435 ;
        RECT 1193.400 200.445 1193.540 202.795 ;
        RECT 1200.300 201.805 1200.440 202.795 ;
        RECT 2359.430 202.115 2359.710 202.485 ;
        RECT 1200.230 201.435 1200.510 201.805 ;
        RECT 2236.150 201.435 2236.430 201.805 ;
        RECT 1703.480 201.125 1703.740 201.270 ;
        RECT 1704.860 201.125 1705.120 201.270 ;
        RECT 1510.730 201.010 1511.010 201.125 ;
        RECT 1511.650 201.010 1511.930 201.125 ;
        RECT 1510.730 200.870 1511.930 201.010 ;
        RECT 1510.730 200.755 1511.010 200.870 ;
        RECT 1511.650 200.755 1511.930 200.870 ;
        RECT 1606.410 200.755 1606.690 201.125 ;
        RECT 1607.790 200.755 1608.070 201.125 ;
        RECT 1703.470 200.755 1703.750 201.125 ;
        RECT 1704.850 200.755 1705.130 201.125 ;
        RECT 1799.610 200.755 1799.890 201.125 ;
        RECT 1800.990 200.755 1801.270 201.125 ;
        RECT 2186.010 200.755 2186.290 201.125 ;
        RECT 1606.420 200.610 1606.680 200.755 ;
        RECT 1607.800 200.610 1608.060 200.755 ;
        RECT 1799.620 200.610 1799.880 200.755 ;
        RECT 1801.000 200.610 1801.260 200.755 ;
        RECT 1193.330 200.075 1193.610 200.445 ;
        RECT 2186.080 199.085 2186.220 200.755 ;
        RECT 2236.220 200.590 2236.360 201.435 ;
        RECT 2221.900 200.445 2222.160 200.590 ;
        RECT 2221.890 200.075 2222.170 200.445 ;
        RECT 2236.160 200.270 2236.420 200.590 ;
        RECT 2359.500 200.445 2359.640 202.115 ;
        RECT 2414.630 201.435 2414.910 201.805 ;
        RECT 2414.700 200.590 2414.840 201.435 ;
        RECT 2380.140 200.445 2380.400 200.590 ;
        RECT 2359.430 200.075 2359.710 200.445 ;
        RECT 2380.130 200.075 2380.410 200.445 ;
        RECT 2414.640 200.270 2414.900 200.590 ;
        RECT 1145.030 198.715 1145.310 199.085 ;
        RECT 2186.010 198.715 2186.290 199.085 ;
      LAYER via2 ;
        RECT 770.130 2722.920 770.410 2723.200 ;
        RECT 1193.330 202.840 1193.610 203.120 ;
        RECT 1200.230 202.840 1200.510 203.120 ;
        RECT 881.910 201.480 882.190 201.760 ;
        RECT 882.830 201.480 883.110 201.760 ;
        RECT 1145.030 201.480 1145.310 201.760 ;
        RECT 1007.490 200.800 1007.770 201.080 ;
        RECT 1096.730 200.120 1097.010 200.400 ;
        RECT 2359.430 202.160 2359.710 202.440 ;
        RECT 1200.230 201.480 1200.510 201.760 ;
        RECT 2236.150 201.480 2236.430 201.760 ;
        RECT 1510.730 200.800 1511.010 201.080 ;
        RECT 1511.650 200.800 1511.930 201.080 ;
        RECT 1606.410 200.800 1606.690 201.080 ;
        RECT 1607.790 200.800 1608.070 201.080 ;
        RECT 1703.470 200.800 1703.750 201.080 ;
        RECT 1704.850 200.800 1705.130 201.080 ;
        RECT 1799.610 200.800 1799.890 201.080 ;
        RECT 1800.990 200.800 1801.270 201.080 ;
        RECT 2186.010 200.800 2186.290 201.080 ;
        RECT 1193.330 200.120 1193.610 200.400 ;
        RECT 2221.890 200.120 2222.170 200.400 ;
        RECT 2414.630 201.480 2414.910 201.760 ;
        RECT 2359.430 200.120 2359.710 200.400 ;
        RECT 2380.130 200.120 2380.410 200.400 ;
        RECT 1145.030 198.760 1145.310 199.040 ;
        RECT 2186.010 198.760 2186.290 199.040 ;
      LAYER met3 ;
        RECT 770.105 2723.220 770.435 2723.225 ;
        RECT 770.105 2723.210 770.690 2723.220 ;
        RECT 770.105 2722.910 770.890 2723.210 ;
        RECT 770.105 2722.900 770.690 2722.910 ;
        RECT 770.105 2722.895 770.435 2722.900 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 1193.305 203.130 1193.635 203.145 ;
        RECT 1200.205 203.130 1200.535 203.145 ;
        RECT 1193.305 202.830 1200.535 203.130 ;
        RECT 1193.305 202.815 1193.635 202.830 ;
        RECT 1200.205 202.815 1200.535 202.830 ;
        RECT 2311.310 202.450 2311.690 202.460 ;
        RECT 2359.405 202.450 2359.735 202.465 ;
        RECT 2311.310 202.150 2359.735 202.450 ;
        RECT 2311.310 202.140 2311.690 202.150 ;
        RECT 2359.405 202.135 2359.735 202.150 ;
        RECT 881.885 201.770 882.215 201.785 ;
        RECT 838.430 201.470 882.215 201.770 ;
        RECT 770.310 200.410 770.690 200.420 ;
        RECT 838.430 200.410 838.730 201.470 ;
        RECT 881.885 201.455 882.215 201.470 ;
        RECT 882.805 201.770 883.135 201.785 ;
        RECT 1145.005 201.770 1145.335 201.785 ;
        RECT 1200.205 201.770 1200.535 201.785 ;
        RECT 1248.710 201.770 1249.090 201.780 ;
        RECT 2236.125 201.770 2236.455 201.785 ;
        RECT 2414.605 201.770 2414.935 201.785 ;
        RECT 882.805 201.470 886.570 201.770 ;
        RECT 882.805 201.455 883.135 201.470 ;
        RECT 886.270 201.090 886.570 201.470 ;
        RECT 1145.005 201.470 1146.010 201.770 ;
        RECT 1145.005 201.455 1145.335 201.470 ;
        RECT 917.510 201.090 917.890 201.100 ;
        RECT 1007.465 201.090 1007.795 201.105 ;
        RECT 886.270 200.790 917.890 201.090 ;
        RECT 917.510 200.780 917.890 200.790 ;
        RECT 976.430 200.790 1007.795 201.090 ;
        RECT 976.430 200.410 976.730 200.790 ;
        RECT 1007.465 200.775 1007.795 200.790 ;
        RECT 770.310 200.110 838.730 200.410 ;
        RECT 918.470 200.110 976.730 200.410 ;
        RECT 1096.705 200.420 1097.035 200.425 ;
        RECT 1096.705 200.410 1097.290 200.420 ;
        RECT 1145.710 200.410 1146.010 201.470 ;
        RECT 1200.205 201.470 1249.090 201.770 ;
        RECT 1200.205 201.455 1200.535 201.470 ;
        RECT 1248.710 201.460 1249.090 201.470 ;
        RECT 1365.590 201.470 1414.650 201.770 ;
        RECT 1193.305 200.410 1193.635 200.425 ;
        RECT 1365.590 200.410 1365.890 201.470 ;
        RECT 1096.705 200.110 1097.670 200.410 ;
        RECT 1145.710 200.110 1193.635 200.410 ;
        RECT 770.310 200.100 770.690 200.110 ;
        RECT 917.510 199.730 917.890 199.740 ;
        RECT 918.470 199.730 918.770 200.110 ;
        RECT 1096.705 200.100 1097.290 200.110 ;
        RECT 1096.705 200.095 1097.035 200.100 ;
        RECT 1193.305 200.095 1193.635 200.110 ;
        RECT 1303.950 200.110 1365.890 200.410 ;
        RECT 1414.350 200.410 1414.650 201.470 ;
        RECT 2236.125 201.470 2294.170 201.770 ;
        RECT 2236.125 201.455 2236.455 201.470 ;
        RECT 1510.705 201.090 1511.035 201.105 ;
        RECT 1463.110 200.790 1511.035 201.090 ;
        RECT 1463.110 200.410 1463.410 200.790 ;
        RECT 1510.705 200.775 1511.035 200.790 ;
        RECT 1511.625 201.090 1511.955 201.105 ;
        RECT 1606.385 201.090 1606.715 201.105 ;
        RECT 1511.625 200.790 1559.090 201.090 ;
        RECT 1511.625 200.775 1511.955 200.790 ;
        RECT 1414.350 200.110 1463.410 200.410 ;
        RECT 1558.790 200.410 1559.090 200.790 ;
        RECT 1559.710 200.790 1606.715 201.090 ;
        RECT 1559.710 200.410 1560.010 200.790 ;
        RECT 1606.385 200.775 1606.715 200.790 ;
        RECT 1607.765 201.090 1608.095 201.105 ;
        RECT 1703.445 201.090 1703.775 201.105 ;
        RECT 1607.765 200.790 1641.890 201.090 ;
        RECT 1607.765 200.775 1608.095 200.790 ;
        RECT 1558.790 200.110 1560.010 200.410 ;
        RECT 1641.590 200.410 1641.890 200.790 ;
        RECT 1656.310 200.790 1703.775 201.090 ;
        RECT 1656.310 200.410 1656.610 200.790 ;
        RECT 1703.445 200.775 1703.775 200.790 ;
        RECT 1704.825 201.090 1705.155 201.105 ;
        RECT 1799.585 201.090 1799.915 201.105 ;
        RECT 1704.825 200.790 1752.290 201.090 ;
        RECT 1704.825 200.775 1705.155 200.790 ;
        RECT 1641.590 200.110 1656.610 200.410 ;
        RECT 1751.990 200.410 1752.290 200.790 ;
        RECT 1752.910 200.790 1799.915 201.090 ;
        RECT 1752.910 200.410 1753.210 200.790 ;
        RECT 1799.585 200.775 1799.915 200.790 ;
        RECT 1800.965 201.090 1801.295 201.105 ;
        RECT 2185.985 201.090 2186.315 201.105 ;
        RECT 1800.965 200.790 1835.090 201.090 ;
        RECT 1800.965 200.775 1801.295 200.790 ;
        RECT 1751.990 200.110 1753.210 200.410 ;
        RECT 1834.790 200.410 1835.090 200.790 ;
        RECT 1849.510 200.790 1945.490 201.090 ;
        RECT 1849.510 200.410 1849.810 200.790 ;
        RECT 1834.790 200.110 1849.810 200.410 ;
        RECT 1945.190 200.410 1945.490 200.790 ;
        RECT 1946.110 200.790 2028.290 201.090 ;
        RECT 1946.110 200.410 1946.410 200.790 ;
        RECT 1945.190 200.110 1946.410 200.410 ;
        RECT 2027.990 200.410 2028.290 200.790 ;
        RECT 2042.710 200.790 2138.690 201.090 ;
        RECT 2042.710 200.410 2043.010 200.790 ;
        RECT 2027.990 200.110 2043.010 200.410 ;
        RECT 2138.390 200.410 2138.690 200.790 ;
        RECT 2139.310 200.790 2186.315 201.090 ;
        RECT 2293.870 201.090 2294.170 201.470 ;
        RECT 2414.605 201.470 2449.650 201.770 ;
        RECT 2414.605 201.455 2414.935 201.470 ;
        RECT 2311.310 201.090 2311.690 201.100 ;
        RECT 2293.870 200.790 2311.690 201.090 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2139.310 200.410 2139.610 200.790 ;
        RECT 2185.985 200.775 2186.315 200.790 ;
        RECT 2311.310 200.780 2311.690 200.790 ;
        RECT 2221.865 200.410 2222.195 200.425 ;
        RECT 2138.390 200.110 2139.610 200.410 ;
        RECT 2221.190 200.110 2222.195 200.410 ;
        RECT 917.510 199.430 918.770 199.730 ;
        RECT 1248.710 199.730 1249.090 199.740 ;
        RECT 1303.950 199.730 1304.250 200.110 ;
        RECT 1248.710 199.430 1304.250 199.730 ;
        RECT 917.510 199.420 917.890 199.430 ;
        RECT 1248.710 199.420 1249.090 199.430 ;
        RECT 1096.910 199.050 1097.290 199.060 ;
        RECT 1145.005 199.050 1145.335 199.065 ;
        RECT 1096.910 198.750 1145.335 199.050 ;
        RECT 1096.910 198.740 1097.290 198.750 ;
        RECT 1145.005 198.735 1145.335 198.750 ;
        RECT 2185.985 199.050 2186.315 199.065 ;
        RECT 2221.190 199.050 2221.490 200.110 ;
        RECT 2221.865 200.095 2222.195 200.110 ;
        RECT 2359.405 200.410 2359.735 200.425 ;
        RECT 2380.105 200.410 2380.435 200.425 ;
        RECT 2359.405 200.110 2380.435 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 2359.405 200.095 2359.735 200.110 ;
        RECT 2380.105 200.095 2380.435 200.110 ;
        RECT 2185.985 198.750 2221.490 199.050 ;
        RECT 2185.985 198.735 2186.315 198.750 ;
      LAYER via3 ;
        RECT 770.340 2722.900 770.660 2723.220 ;
        RECT 2311.340 202.140 2311.660 202.460 ;
        RECT 770.340 200.100 770.660 200.420 ;
        RECT 917.540 200.780 917.860 201.100 ;
        RECT 917.540 199.420 917.860 199.740 ;
        RECT 1096.940 200.100 1097.260 200.420 ;
        RECT 1248.740 201.460 1249.060 201.780 ;
        RECT 2311.340 200.780 2311.660 201.100 ;
        RECT 1248.740 199.420 1249.060 199.740 ;
        RECT 1096.940 198.740 1097.260 199.060 ;
      LAYER met4 ;
        RECT 770.335 2722.895 770.665 2723.225 ;
        RECT 770.350 200.425 770.650 2722.895 ;
        RECT 2311.335 202.135 2311.665 202.465 ;
        RECT 1248.735 201.455 1249.065 201.785 ;
        RECT 917.535 200.775 917.865 201.105 ;
        RECT 770.335 200.095 770.665 200.425 ;
        RECT 917.550 199.745 917.850 200.775 ;
        RECT 1096.935 200.095 1097.265 200.425 ;
        RECT 917.535 199.415 917.865 199.745 ;
        RECT 1096.950 199.065 1097.250 200.095 ;
        RECT 1248.750 199.745 1249.050 201.455 ;
        RECT 2311.350 201.105 2311.650 202.135 ;
        RECT 2311.335 200.775 2311.665 201.105 ;
        RECT 1248.735 199.415 1249.065 199.745 ;
        RECT 1096.935 198.735 1097.265 199.065 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2249.010 2552.960 2249.330 2553.020 ;
        RECT 2899.450 2552.960 2899.770 2553.020 ;
        RECT 2249.010 2552.820 2899.770 2552.960 ;
        RECT 2249.010 2552.760 2249.330 2552.820 ;
        RECT 2899.450 2552.760 2899.770 2552.820 ;
      LAYER via ;
        RECT 2249.040 2552.760 2249.300 2553.020 ;
        RECT 2899.480 2552.760 2899.740 2553.020 ;
      LAYER met2 ;
        RECT 1157.010 2723.130 1157.570 2731.680 ;
        RECT 1157.910 2723.130 1158.190 2723.245 ;
        RECT 1157.010 2722.990 1158.190 2723.130 ;
        RECT 1157.010 2722.680 1157.570 2722.990 ;
        RECT 1157.910 2722.875 1158.190 2722.990 ;
        RECT 2249.030 2714.035 2249.310 2714.405 ;
        RECT 2249.100 2553.050 2249.240 2714.035 ;
        RECT 2249.040 2552.730 2249.300 2553.050 ;
        RECT 2899.480 2552.730 2899.740 2553.050 ;
        RECT 2899.540 2551.885 2899.680 2552.730 ;
        RECT 2899.470 2551.515 2899.750 2551.885 ;
      LAYER via2 ;
        RECT 1157.910 2722.920 1158.190 2723.200 ;
        RECT 2249.030 2714.080 2249.310 2714.360 ;
        RECT 2899.470 2551.560 2899.750 2551.840 ;
      LAYER met3 ;
        RECT 1157.885 2723.220 1158.215 2723.225 ;
        RECT 1157.630 2723.210 1158.215 2723.220 ;
        RECT 1157.430 2722.910 1158.215 2723.210 ;
        RECT 1157.630 2722.900 1158.215 2722.910 ;
        RECT 1157.885 2722.895 1158.215 2722.900 ;
        RECT 1157.630 2716.100 1158.010 2716.420 ;
        RECT 1157.670 2714.370 1157.970 2716.100 ;
        RECT 2249.005 2714.370 2249.335 2714.385 ;
        RECT 1157.670 2714.070 2249.335 2714.370 ;
        RECT 2249.005 2714.055 2249.335 2714.070 ;
        RECT 2899.445 2551.850 2899.775 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2899.445 2551.550 2924.800 2551.850 ;
        RECT 2899.445 2551.535 2899.775 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
      LAYER via3 ;
        RECT 1157.660 2722.900 1157.980 2723.220 ;
        RECT 1157.660 2716.100 1157.980 2716.420 ;
      LAYER met4 ;
        RECT 1157.655 2722.895 1157.985 2723.225 ;
        RECT 1157.670 2716.425 1157.970 2722.895 ;
        RECT 1157.655 2716.095 1157.985 2716.425 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1200.210 2781.100 1200.530 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 1200.210 2780.960 2901.150 2781.100 ;
        RECT 1200.210 2780.900 1200.530 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 1200.240 2780.900 1200.500 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 1200.240 2780.870 1200.500 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 1200.300 2731.970 1200.440 2780.870 ;
        RECT 1198.920 2731.830 1200.440 2731.970 ;
        RECT 1195.650 2731.290 1196.210 2731.680 ;
        RECT 1198.920 2731.290 1199.060 2731.830 ;
        RECT 1195.650 2731.150 1199.060 2731.290 ;
        RECT 1195.650 2722.680 1196.210 2731.150 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.710 3015.700 1235.030 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1234.710 3015.560 2901.150 3015.700 ;
        RECT 1234.710 3015.500 1235.030 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1234.740 3015.500 1235.000 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1234.740 3015.470 1235.000 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1234.800 2731.680 1234.940 3015.470 ;
        RECT 1234.750 2722.680 1235.310 2731.680 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1276.110 3250.300 1276.430 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1276.110 3250.160 2901.150 3250.300 ;
        RECT 1276.110 3250.100 1276.430 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1276.140 3250.100 1276.400 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1276.140 3250.070 1276.400 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1276.200 2731.970 1276.340 3250.070 ;
        RECT 1275.280 2731.830 1276.340 2731.970 ;
        RECT 1273.390 2731.290 1273.950 2731.680 ;
        RECT 1275.280 2731.290 1275.420 2731.830 ;
        RECT 1273.390 2731.150 1275.420 2731.290 ;
        RECT 1273.390 2722.680 1273.950 2731.150 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.510 3484.900 1317.830 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1317.510 3484.760 2901.150 3484.900 ;
        RECT 1317.510 3484.700 1317.830 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1317.540 3484.700 1317.800 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1317.540 3484.670 1317.800 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1317.600 2731.970 1317.740 3484.670 ;
        RECT 1314.380 2731.830 1317.740 2731.970 ;
        RECT 1312.030 2730.610 1312.590 2731.680 ;
        RECT 1314.380 2730.610 1314.520 2731.830 ;
        RECT 1312.030 2730.470 1314.520 2730.610 ;
        RECT 1312.030 2722.680 1312.590 2730.470 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.010 3502.580 1352.330 3502.640 ;
        RECT 2635.870 3502.580 2636.190 3502.640 ;
        RECT 1352.010 3502.440 2636.190 3502.580 ;
        RECT 1352.010 3502.380 1352.330 3502.440 ;
        RECT 2635.870 3502.380 2636.190 3502.440 ;
      LAYER via ;
        RECT 1352.040 3502.380 1352.300 3502.640 ;
        RECT 2635.900 3502.380 2636.160 3502.640 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.670 2636.100 3517.600 ;
        RECT 1352.040 3502.350 1352.300 3502.670 ;
        RECT 2635.900 3502.350 2636.160 3502.670 ;
        RECT 1351.130 2731.290 1351.690 2731.680 ;
        RECT 1352.100 2731.290 1352.240 3502.350 ;
        RECT 1351.130 2731.150 1352.240 2731.290 ;
        RECT 1351.130 2722.680 1351.690 2731.150 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1393.410 3504.280 1393.730 3504.340 ;
        RECT 2311.570 3504.280 2311.890 3504.340 ;
        RECT 1393.410 3504.140 2311.890 3504.280 ;
        RECT 1393.410 3504.080 1393.730 3504.140 ;
        RECT 2311.570 3504.080 2311.890 3504.140 ;
      LAYER via ;
        RECT 1393.440 3504.080 1393.700 3504.340 ;
        RECT 2311.600 3504.080 2311.860 3504.340 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3504.370 2311.800 3517.600 ;
        RECT 1393.440 3504.050 1393.700 3504.370 ;
        RECT 2311.600 3504.050 2311.860 3504.370 ;
        RECT 1389.770 2730.610 1390.330 2731.680 ;
        RECT 1393.500 2730.610 1393.640 3504.050 ;
        RECT 1389.770 2730.470 1393.640 2730.610 ;
        RECT 1389.770 2722.680 1390.330 2730.470 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1434.810 3500.540 1435.130 3500.600 ;
        RECT 1987.270 3500.540 1987.590 3500.600 ;
        RECT 1434.810 3500.400 1987.590 3500.540 ;
        RECT 1434.810 3500.340 1435.130 3500.400 ;
        RECT 1987.270 3500.340 1987.590 3500.400 ;
      LAYER via ;
        RECT 1434.840 3500.340 1435.100 3500.600 ;
        RECT 1987.300 3500.340 1987.560 3500.600 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3500.630 1987.500 3517.600 ;
        RECT 1434.840 3500.310 1435.100 3500.630 ;
        RECT 1987.300 3500.310 1987.560 3500.630 ;
        RECT 1434.900 2731.970 1435.040 3500.310 ;
        RECT 1431.680 2731.830 1435.040 2731.970 ;
        RECT 1428.410 2731.290 1428.970 2731.680 ;
        RECT 1431.680 2731.290 1431.820 2731.830 ;
        RECT 1428.410 2731.150 1431.820 2731.290 ;
        RECT 1428.410 2722.680 1428.970 2731.150 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1469.310 3499.180 1469.630 3499.240 ;
        RECT 1662.510 3499.180 1662.830 3499.240 ;
        RECT 1469.310 3499.040 1662.830 3499.180 ;
        RECT 1469.310 3498.980 1469.630 3499.040 ;
        RECT 1662.510 3498.980 1662.830 3499.040 ;
      LAYER via ;
        RECT 1469.340 3498.980 1469.600 3499.240 ;
        RECT 1662.540 3498.980 1662.800 3499.240 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3499.270 1662.740 3517.600 ;
        RECT 1469.340 3498.950 1469.600 3499.270 ;
        RECT 1662.540 3498.950 1662.800 3499.270 ;
        RECT 1467.510 2731.290 1468.070 2731.680 ;
        RECT 1469.400 2731.290 1469.540 3498.950 ;
        RECT 1467.510 2731.150 1469.540 2731.290 ;
        RECT 1467.510 2722.680 1468.070 2731.150 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3498.840 1338.530 3498.900 ;
        RECT 1504.270 3498.840 1504.590 3498.900 ;
        RECT 1338.210 3498.700 1504.590 3498.840 ;
        RECT 1338.210 3498.640 1338.530 3498.700 ;
        RECT 1504.270 3498.640 1504.590 3498.700 ;
      LAYER via ;
        RECT 1338.240 3498.640 1338.500 3498.900 ;
        RECT 1504.300 3498.640 1504.560 3498.900 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3498.930 1338.440 3517.600 ;
        RECT 1338.240 3498.610 1338.500 3498.930 ;
        RECT 1504.300 3498.610 1504.560 3498.930 ;
        RECT 1504.360 2731.290 1504.500 3498.610 ;
        RECT 1506.150 2731.290 1506.710 2731.680 ;
        RECT 1504.360 2731.150 1506.710 2731.290 ;
        RECT 1506.150 2722.680 1506.710 2731.150 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 809.285 2714.305 809.455 2723.655 ;
        RECT 844.245 2714.305 844.415 2715.155 ;
        RECT 869.085 2714.305 869.255 2715.155 ;
        RECT 869.545 2714.305 869.715 2715.495 ;
        RECT 893.465 2714.305 893.635 2715.495 ;
        RECT 940.845 2714.305 941.015 2715.155 ;
        RECT 965.685 2714.305 965.855 2715.155 ;
        RECT 966.145 2714.305 966.315 2715.495 ;
        RECT 990.065 2714.305 990.235 2715.495 ;
        RECT 1037.445 2714.305 1037.615 2715.155 ;
        RECT 1078.845 2714.305 1079.015 2715.155 ;
        RECT 1318.505 2714.475 1318.675 2714.815 ;
        RECT 1207.645 2714.305 1208.735 2714.475 ;
        RECT 1317.585 2714.305 1318.675 2714.475 ;
        RECT 1352.545 2714.305 1352.715 2715.495 ;
        RECT 1376.465 2714.305 1376.635 2715.495 ;
        RECT 1423.845 2714.305 1424.015 2715.155 ;
        RECT 1448.685 2714.305 1448.855 2715.155 ;
        RECT 1449.145 2714.305 1449.315 2715.495 ;
        RECT 1473.065 2714.305 1473.235 2715.495 ;
        RECT 1497.445 2714.305 1497.615 2715.835 ;
        RECT 1544.365 2714.475 1544.535 2715.835 ;
        RECT 1544.365 2714.305 1545.455 2714.475 ;
        RECT 1545.745 2714.305 1545.915 2715.495 ;
        RECT 1569.665 2714.305 1569.835 2715.495 ;
        RECT 1617.045 2714.305 1617.215 2715.155 ;
        RECT 1642.345 2714.985 1642.975 2715.155 ;
        RECT 1642.805 2714.645 1642.975 2714.985 ;
        RECT 1732.965 2714.645 1733.135 2715.835 ;
        RECT 1779.885 2714.985 1780.055 2715.835 ;
        RECT 1829.105 2714.305 1829.275 2715.155 ;
      LAYER mcon ;
        RECT 809.285 2723.485 809.455 2723.655 ;
        RECT 1497.445 2715.665 1497.615 2715.835 ;
        RECT 869.545 2715.325 869.715 2715.495 ;
        RECT 844.245 2714.985 844.415 2715.155 ;
        RECT 869.085 2714.985 869.255 2715.155 ;
        RECT 893.465 2715.325 893.635 2715.495 ;
        RECT 966.145 2715.325 966.315 2715.495 ;
        RECT 940.845 2714.985 941.015 2715.155 ;
        RECT 965.685 2714.985 965.855 2715.155 ;
        RECT 990.065 2715.325 990.235 2715.495 ;
        RECT 1352.545 2715.325 1352.715 2715.495 ;
        RECT 1037.445 2714.985 1037.615 2715.155 ;
        RECT 1078.845 2714.985 1079.015 2715.155 ;
        RECT 1318.505 2714.645 1318.675 2714.815 ;
        RECT 1208.565 2714.305 1208.735 2714.475 ;
        RECT 1376.465 2715.325 1376.635 2715.495 ;
        RECT 1449.145 2715.325 1449.315 2715.495 ;
        RECT 1423.845 2714.985 1424.015 2715.155 ;
        RECT 1448.685 2714.985 1448.855 2715.155 ;
        RECT 1473.065 2715.325 1473.235 2715.495 ;
        RECT 1544.365 2715.665 1544.535 2715.835 ;
        RECT 1732.965 2715.665 1733.135 2715.835 ;
        RECT 1545.745 2715.325 1545.915 2715.495 ;
        RECT 1545.285 2714.305 1545.455 2714.475 ;
        RECT 1569.665 2715.325 1569.835 2715.495 ;
        RECT 1617.045 2714.985 1617.215 2715.155 ;
        RECT 1779.885 2715.665 1780.055 2715.835 ;
        RECT 1829.105 2714.985 1829.275 2715.155 ;
      LAYER met1 ;
        RECT 809.210 2723.640 809.530 2723.700 ;
        RECT 809.015 2723.500 809.530 2723.640 ;
        RECT 809.210 2723.440 809.530 2723.500 ;
        RECT 1497.385 2715.820 1497.675 2715.865 ;
        RECT 1544.305 2715.820 1544.595 2715.865 ;
        RECT 1497.385 2715.680 1544.595 2715.820 ;
        RECT 1497.385 2715.635 1497.675 2715.680 ;
        RECT 1544.305 2715.635 1544.595 2715.680 ;
        RECT 1732.905 2715.820 1733.195 2715.865 ;
        RECT 1779.825 2715.820 1780.115 2715.865 ;
        RECT 1732.905 2715.680 1780.115 2715.820 ;
        RECT 1732.905 2715.635 1733.195 2715.680 ;
        RECT 1779.825 2715.635 1780.115 2715.680 ;
        RECT 869.485 2715.480 869.775 2715.525 ;
        RECT 893.405 2715.480 893.695 2715.525 ;
        RECT 869.485 2715.340 893.695 2715.480 ;
        RECT 869.485 2715.295 869.775 2715.340 ;
        RECT 893.405 2715.295 893.695 2715.340 ;
        RECT 966.085 2715.480 966.375 2715.525 ;
        RECT 990.005 2715.480 990.295 2715.525 ;
        RECT 966.085 2715.340 990.295 2715.480 ;
        RECT 966.085 2715.295 966.375 2715.340 ;
        RECT 990.005 2715.295 990.295 2715.340 ;
        RECT 1352.485 2715.480 1352.775 2715.525 ;
        RECT 1376.405 2715.480 1376.695 2715.525 ;
        RECT 1352.485 2715.340 1376.695 2715.480 ;
        RECT 1352.485 2715.295 1352.775 2715.340 ;
        RECT 1376.405 2715.295 1376.695 2715.340 ;
        RECT 1449.085 2715.480 1449.375 2715.525 ;
        RECT 1473.005 2715.480 1473.295 2715.525 ;
        RECT 1449.085 2715.340 1473.295 2715.480 ;
        RECT 1449.085 2715.295 1449.375 2715.340 ;
        RECT 1473.005 2715.295 1473.295 2715.340 ;
        RECT 1545.685 2715.480 1545.975 2715.525 ;
        RECT 1569.605 2715.480 1569.895 2715.525 ;
        RECT 1545.685 2715.340 1569.895 2715.480 ;
        RECT 1545.685 2715.295 1545.975 2715.340 ;
        RECT 1569.605 2715.295 1569.895 2715.340 ;
        RECT 844.185 2715.140 844.475 2715.185 ;
        RECT 869.025 2715.140 869.315 2715.185 ;
        RECT 844.185 2715.000 869.315 2715.140 ;
        RECT 844.185 2714.955 844.475 2715.000 ;
        RECT 869.025 2714.955 869.315 2715.000 ;
        RECT 940.785 2715.140 941.075 2715.185 ;
        RECT 965.625 2715.140 965.915 2715.185 ;
        RECT 940.785 2715.000 965.915 2715.140 ;
        RECT 940.785 2714.955 941.075 2715.000 ;
        RECT 965.625 2714.955 965.915 2715.000 ;
        RECT 1037.385 2715.140 1037.675 2715.185 ;
        RECT 1078.785 2715.140 1079.075 2715.185 ;
        RECT 1037.385 2715.000 1079.075 2715.140 ;
        RECT 1037.385 2714.955 1037.675 2715.000 ;
        RECT 1078.785 2714.955 1079.075 2715.000 ;
        RECT 1423.785 2715.140 1424.075 2715.185 ;
        RECT 1448.625 2715.140 1448.915 2715.185 ;
        RECT 1423.785 2715.000 1448.915 2715.140 ;
        RECT 1423.785 2714.955 1424.075 2715.000 ;
        RECT 1448.625 2714.955 1448.915 2715.000 ;
        RECT 1616.985 2715.140 1617.275 2715.185 ;
        RECT 1642.285 2715.140 1642.575 2715.185 ;
        RECT 1616.985 2715.000 1642.575 2715.140 ;
        RECT 1616.985 2714.955 1617.275 2715.000 ;
        RECT 1642.285 2714.955 1642.575 2715.000 ;
        RECT 1779.825 2714.955 1780.115 2715.185 ;
        RECT 1829.045 2715.140 1829.335 2715.185 ;
        RECT 1829.045 2715.000 1849.960 2715.140 ;
        RECT 1829.045 2714.955 1829.335 2715.000 ;
        RECT 1318.445 2714.800 1318.735 2714.845 ;
        RECT 1642.745 2714.800 1643.035 2714.845 ;
        RECT 1318.445 2714.660 1352.240 2714.800 ;
        RECT 1318.445 2714.615 1318.735 2714.660 ;
        RECT 809.225 2714.460 809.515 2714.505 ;
        RECT 844.185 2714.460 844.475 2714.505 ;
        RECT 809.225 2714.320 844.475 2714.460 ;
        RECT 809.225 2714.275 809.515 2714.320 ;
        RECT 844.185 2714.275 844.475 2714.320 ;
        RECT 869.025 2714.460 869.315 2714.505 ;
        RECT 869.485 2714.460 869.775 2714.505 ;
        RECT 869.025 2714.320 869.775 2714.460 ;
        RECT 869.025 2714.275 869.315 2714.320 ;
        RECT 869.485 2714.275 869.775 2714.320 ;
        RECT 893.405 2714.460 893.695 2714.505 ;
        RECT 940.785 2714.460 941.075 2714.505 ;
        RECT 893.405 2714.320 941.075 2714.460 ;
        RECT 893.405 2714.275 893.695 2714.320 ;
        RECT 940.785 2714.275 941.075 2714.320 ;
        RECT 965.625 2714.460 965.915 2714.505 ;
        RECT 966.085 2714.460 966.375 2714.505 ;
        RECT 965.625 2714.320 966.375 2714.460 ;
        RECT 965.625 2714.275 965.915 2714.320 ;
        RECT 966.085 2714.275 966.375 2714.320 ;
        RECT 990.005 2714.460 990.295 2714.505 ;
        RECT 1037.385 2714.460 1037.675 2714.505 ;
        RECT 990.005 2714.320 1037.675 2714.460 ;
        RECT 990.005 2714.275 990.295 2714.320 ;
        RECT 1037.385 2714.275 1037.675 2714.320 ;
        RECT 1078.785 2714.460 1079.075 2714.505 ;
        RECT 1207.585 2714.460 1207.875 2714.505 ;
        RECT 1078.785 2714.320 1207.875 2714.460 ;
        RECT 1078.785 2714.275 1079.075 2714.320 ;
        RECT 1207.585 2714.275 1207.875 2714.320 ;
        RECT 1208.505 2714.460 1208.795 2714.505 ;
        RECT 1317.525 2714.460 1317.815 2714.505 ;
        RECT 1208.505 2714.320 1317.815 2714.460 ;
        RECT 1352.100 2714.460 1352.240 2714.660 ;
        RECT 1642.745 2714.660 1658.600 2714.800 ;
        RECT 1642.745 2714.615 1643.035 2714.660 ;
        RECT 1352.485 2714.460 1352.775 2714.505 ;
        RECT 1352.100 2714.320 1352.775 2714.460 ;
        RECT 1208.505 2714.275 1208.795 2714.320 ;
        RECT 1317.525 2714.275 1317.815 2714.320 ;
        RECT 1352.485 2714.275 1352.775 2714.320 ;
        RECT 1376.405 2714.460 1376.695 2714.505 ;
        RECT 1423.785 2714.460 1424.075 2714.505 ;
        RECT 1376.405 2714.320 1424.075 2714.460 ;
        RECT 1376.405 2714.275 1376.695 2714.320 ;
        RECT 1423.785 2714.275 1424.075 2714.320 ;
        RECT 1448.625 2714.460 1448.915 2714.505 ;
        RECT 1449.085 2714.460 1449.375 2714.505 ;
        RECT 1448.625 2714.320 1449.375 2714.460 ;
        RECT 1448.625 2714.275 1448.915 2714.320 ;
        RECT 1449.085 2714.275 1449.375 2714.320 ;
        RECT 1473.005 2714.460 1473.295 2714.505 ;
        RECT 1497.385 2714.460 1497.675 2714.505 ;
        RECT 1473.005 2714.320 1497.675 2714.460 ;
        RECT 1473.005 2714.275 1473.295 2714.320 ;
        RECT 1497.385 2714.275 1497.675 2714.320 ;
        RECT 1545.225 2714.460 1545.515 2714.505 ;
        RECT 1545.685 2714.460 1545.975 2714.505 ;
        RECT 1545.225 2714.320 1545.975 2714.460 ;
        RECT 1545.225 2714.275 1545.515 2714.320 ;
        RECT 1545.685 2714.275 1545.975 2714.320 ;
        RECT 1569.605 2714.460 1569.895 2714.505 ;
        RECT 1616.985 2714.460 1617.275 2714.505 ;
        RECT 1569.605 2714.320 1617.275 2714.460 ;
        RECT 1658.460 2714.460 1658.600 2714.660 ;
        RECT 1732.905 2714.615 1733.195 2714.845 ;
        RECT 1732.980 2714.460 1733.120 2714.615 ;
        RECT 1658.460 2714.320 1733.120 2714.460 ;
        RECT 1779.900 2714.460 1780.040 2714.955 ;
        RECT 1829.045 2714.460 1829.335 2714.505 ;
        RECT 1779.900 2714.320 1829.335 2714.460 ;
        RECT 1849.820 2714.460 1849.960 2715.000 ;
        RECT 2901.290 2714.460 2901.610 2714.520 ;
        RECT 1849.820 2714.320 2901.610 2714.460 ;
        RECT 1569.605 2714.275 1569.895 2714.320 ;
        RECT 1616.985 2714.275 1617.275 2714.320 ;
        RECT 1829.045 2714.275 1829.335 2714.320 ;
        RECT 2901.290 2714.260 2901.610 2714.320 ;
      LAYER via ;
        RECT 809.240 2723.440 809.500 2723.700 ;
        RECT 2901.320 2714.260 2901.580 2714.520 ;
      LAYER met2 ;
        RECT 807.870 2723.810 808.430 2731.680 ;
        RECT 807.870 2723.730 809.440 2723.810 ;
        RECT 807.870 2723.670 809.500 2723.730 ;
        RECT 807.870 2722.680 808.430 2723.670 ;
        RECT 809.240 2723.410 809.500 2723.670 ;
        RECT 2901.320 2714.230 2901.580 2714.550 ;
        RECT 2901.380 439.805 2901.520 2714.230 ;
        RECT 2901.310 439.435 2901.590 439.805 ;
      LAYER via2 ;
        RECT 2901.310 439.480 2901.590 439.760 ;
      LAYER met3 ;
        RECT 2901.285 439.770 2901.615 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2901.285 439.470 2924.800 439.770 ;
        RECT 2901.285 439.455 2901.615 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3500.200 1014.230 3500.260 ;
        RECT 1538.770 3500.200 1539.090 3500.260 ;
        RECT 1013.910 3500.060 1539.090 3500.200 ;
        RECT 1013.910 3500.000 1014.230 3500.060 ;
        RECT 1538.770 3500.000 1539.090 3500.060 ;
      LAYER via ;
        RECT 1013.940 3500.000 1014.200 3500.260 ;
        RECT 1538.800 3500.000 1539.060 3500.260 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3500.290 1014.140 3517.600 ;
        RECT 1013.940 3499.970 1014.200 3500.290 ;
        RECT 1538.800 3499.970 1539.060 3500.290 ;
        RECT 1538.860 2731.970 1539.000 3499.970 ;
        RECT 1538.860 2731.830 1542.680 2731.970 ;
        RECT 1542.540 2731.290 1542.680 2731.830 ;
        RECT 1544.790 2731.290 1545.350 2731.680 ;
        RECT 1542.540 2731.150 1545.350 2731.290 ;
        RECT 1544.790 2722.680 1545.350 2731.150 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3504.620 689.470 3504.680 ;
        RECT 1580.170 3504.620 1580.490 3504.680 ;
        RECT 689.150 3504.480 1580.490 3504.620 ;
        RECT 689.150 3504.420 689.470 3504.480 ;
        RECT 1580.170 3504.420 1580.490 3504.480 ;
      LAYER via ;
        RECT 689.180 3504.420 689.440 3504.680 ;
        RECT 1580.200 3504.420 1580.460 3504.680 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3504.710 689.380 3517.600 ;
        RECT 689.180 3504.390 689.440 3504.710 ;
        RECT 1580.200 3504.390 1580.460 3504.710 ;
        RECT 1580.260 2731.970 1580.400 3504.390 ;
        RECT 1580.260 2731.830 1581.320 2731.970 ;
        RECT 1581.180 2731.290 1581.320 2731.830 ;
        RECT 1583.890 2731.290 1584.450 2731.680 ;
        RECT 1581.180 2731.150 1584.450 2731.290 ;
        RECT 1583.890 2722.680 1584.450 2731.150 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.920 365.170 3502.980 ;
        RECT 1621.570 3502.920 1621.890 3502.980 ;
        RECT 364.850 3502.780 1621.890 3502.920 ;
        RECT 364.850 3502.720 365.170 3502.780 ;
        RECT 1621.570 3502.720 1621.890 3502.780 ;
      LAYER via ;
        RECT 364.880 3502.720 365.140 3502.980 ;
        RECT 1621.600 3502.720 1621.860 3502.980 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3503.010 365.080 3517.600 ;
        RECT 364.880 3502.690 365.140 3503.010 ;
        RECT 1621.600 3502.690 1621.860 3503.010 ;
        RECT 1621.660 2731.290 1621.800 3502.690 ;
        RECT 1622.530 2731.290 1623.090 2731.680 ;
        RECT 1621.660 2731.150 1623.090 2731.290 ;
        RECT 1622.530 2722.680 1623.090 2731.150 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1656.550 3501.475 1656.830 3501.845 ;
        RECT 1656.620 2731.970 1656.760 3501.475 ;
        RECT 1656.620 2731.830 1659.520 2731.970 ;
        RECT 1659.380 2731.290 1659.520 2731.830 ;
        RECT 1661.170 2731.290 1661.730 2731.680 ;
        RECT 1659.380 2731.150 1661.730 2731.290 ;
        RECT 1661.170 2722.680 1661.730 2731.150 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1656.550 3501.520 1656.830 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1656.525 3501.810 1656.855 3501.825 ;
        RECT 40.545 3501.510 1656.855 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 1656.525 3501.495 1656.855 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1697.470 3263.900 1697.790 3263.960 ;
        RECT 15.250 3263.760 1697.790 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1697.470 3263.700 1697.790 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1697.500 3263.700 1697.760 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1697.500 3263.670 1697.760 3263.990 ;
        RECT 1697.560 2731.970 1697.700 3263.670 ;
        RECT 1697.560 2731.830 1698.160 2731.970 ;
        RECT 1698.020 2731.290 1698.160 2731.830 ;
        RECT 1700.270 2731.290 1700.830 2731.680 ;
        RECT 1698.020 2731.150 1700.830 2731.290 ;
        RECT 1700.270 2722.680 1700.830 2731.150 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 1738.870 2974.220 1739.190 2974.280 ;
        RECT 16.170 2974.080 1739.190 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 1738.870 2974.020 1739.190 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 1738.900 2974.020 1739.160 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 1738.900 2973.990 1739.160 2974.310 ;
        RECT 1738.960 2731.680 1739.100 2973.990 ;
        RECT 1738.910 2722.680 1739.470 2731.680 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2745.060 15.110 2745.120 ;
        RECT 1777.510 2745.060 1777.830 2745.120 ;
        RECT 14.790 2744.920 1777.830 2745.060 ;
        RECT 14.790 2744.860 15.110 2744.920 ;
        RECT 1777.510 2744.860 1777.830 2744.920 ;
      LAYER via ;
        RECT 14.820 2744.860 15.080 2745.120 ;
        RECT 1777.540 2744.860 1777.800 2745.120 ;
      LAYER met2 ;
        RECT 14.820 2744.830 15.080 2745.150 ;
        RECT 1777.540 2744.830 1777.800 2745.150 ;
        RECT 14.880 2693.325 15.020 2744.830 ;
        RECT 1777.600 2731.680 1777.740 2744.830 ;
        RECT 1777.550 2722.680 1778.110 2731.680 ;
        RECT 14.810 2692.955 15.090 2693.325 ;
      LAYER via2 ;
        RECT 14.810 2693.000 15.090 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 14.785 2693.290 15.115 2693.305 ;
        RECT -4.800 2692.990 15.115 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 14.785 2692.975 15.115 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 27.210 2726.360 27.530 2726.420 ;
        RECT 1815.230 2726.360 1815.550 2726.420 ;
        RECT 27.210 2726.220 1815.550 2726.360 ;
        RECT 27.210 2726.160 27.530 2726.220 ;
        RECT 1815.230 2726.160 1815.550 2726.220 ;
        RECT 13.870 2405.740 14.190 2405.800 ;
        RECT 27.210 2405.740 27.530 2405.800 ;
        RECT 13.870 2405.600 27.530 2405.740 ;
        RECT 13.870 2405.540 14.190 2405.600 ;
        RECT 27.210 2405.540 27.530 2405.600 ;
      LAYER via ;
        RECT 27.240 2726.160 27.500 2726.420 ;
        RECT 1815.260 2726.160 1815.520 2726.420 ;
        RECT 13.900 2405.540 14.160 2405.800 ;
        RECT 27.240 2405.540 27.500 2405.800 ;
      LAYER met2 ;
        RECT 1816.650 2726.530 1817.210 2731.680 ;
        RECT 1815.320 2726.450 1817.210 2726.530 ;
        RECT 27.240 2726.130 27.500 2726.450 ;
        RECT 1815.260 2726.390 1817.210 2726.450 ;
        RECT 1815.260 2726.130 1815.520 2726.390 ;
        RECT 27.300 2405.830 27.440 2726.130 ;
        RECT 1816.650 2722.680 1817.210 2726.390 ;
        RECT 13.900 2405.685 14.160 2405.830 ;
        RECT 13.890 2405.315 14.170 2405.685 ;
        RECT 27.240 2405.510 27.500 2405.830 ;
      LAYER via2 ;
        RECT 13.890 2405.360 14.170 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 13.865 2405.650 14.195 2405.665 ;
        RECT -4.800 2405.350 14.195 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 13.865 2405.335 14.195 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.290 2744.380 26.610 2744.440 ;
        RECT 1855.250 2744.380 1855.570 2744.440 ;
        RECT 26.290 2744.240 1855.570 2744.380 ;
        RECT 26.290 2744.180 26.610 2744.240 ;
        RECT 1855.250 2744.180 1855.570 2744.240 ;
        RECT 13.870 2124.220 14.190 2124.280 ;
        RECT 26.290 2124.220 26.610 2124.280 ;
        RECT 13.870 2124.080 26.610 2124.220 ;
        RECT 13.870 2124.020 14.190 2124.080 ;
        RECT 26.290 2124.020 26.610 2124.080 ;
      LAYER via ;
        RECT 26.320 2744.180 26.580 2744.440 ;
        RECT 1855.280 2744.180 1855.540 2744.440 ;
        RECT 13.900 2124.020 14.160 2124.280 ;
        RECT 26.320 2124.020 26.580 2124.280 ;
      LAYER met2 ;
        RECT 26.320 2744.150 26.580 2744.470 ;
        RECT 1855.280 2744.150 1855.540 2744.470 ;
        RECT 26.380 2124.310 26.520 2744.150 ;
        RECT 1855.340 2731.680 1855.480 2744.150 ;
        RECT 1855.290 2722.680 1855.850 2731.680 ;
        RECT 13.900 2123.990 14.160 2124.310 ;
        RECT 26.320 2123.990 26.580 2124.310 ;
        RECT 13.960 2118.725 14.100 2123.990 ;
        RECT 13.890 2118.355 14.170 2118.725 ;
      LAYER via2 ;
        RECT 13.890 2118.400 14.170 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 13.865 2118.690 14.195 2118.705 ;
        RECT -4.800 2118.390 14.195 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 13.865 2118.375 14.195 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.830 2743.020 26.150 2743.080 ;
        RECT 1893.890 2743.020 1894.210 2743.080 ;
        RECT 25.830 2742.880 1894.210 2743.020 ;
        RECT 25.830 2742.820 26.150 2742.880 ;
        RECT 1893.890 2742.820 1894.210 2742.880 ;
        RECT 13.870 1834.880 14.190 1834.940 ;
        RECT 25.830 1834.880 26.150 1834.940 ;
        RECT 13.870 1834.740 26.150 1834.880 ;
        RECT 13.870 1834.680 14.190 1834.740 ;
        RECT 25.830 1834.680 26.150 1834.740 ;
      LAYER via ;
        RECT 25.860 2742.820 26.120 2743.080 ;
        RECT 1893.920 2742.820 1894.180 2743.080 ;
        RECT 13.900 1834.680 14.160 1834.940 ;
        RECT 25.860 1834.680 26.120 1834.940 ;
      LAYER met2 ;
        RECT 25.860 2742.790 26.120 2743.110 ;
        RECT 1893.920 2742.790 1894.180 2743.110 ;
        RECT 25.920 1834.970 26.060 2742.790 ;
        RECT 1893.980 2731.680 1894.120 2742.790 ;
        RECT 1893.930 2722.680 1894.490 2731.680 ;
        RECT 13.900 1834.650 14.160 1834.970 ;
        RECT 25.860 1834.650 26.120 1834.970 ;
        RECT 13.960 1831.085 14.100 1834.650 ;
        RECT 13.890 1830.715 14.170 1831.085 ;
      LAYER via2 ;
        RECT 13.890 1830.760 14.170 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 13.865 1831.050 14.195 1831.065 ;
        RECT -4.800 1830.750 14.195 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 13.865 1830.735 14.195 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 847.925 2720.425 848.095 2723.655 ;
      LAYER mcon ;
        RECT 847.925 2723.485 848.095 2723.655 ;
      LAYER met1 ;
        RECT 847.850 2723.640 848.170 2723.700 ;
        RECT 847.655 2723.500 848.170 2723.640 ;
        RECT 847.850 2723.440 848.170 2723.500 ;
        RECT 847.865 2720.580 848.155 2720.625 ;
        RECT 2889.330 2720.580 2889.650 2720.640 ;
        RECT 847.865 2720.440 2889.650 2720.580 ;
        RECT 847.865 2720.395 848.155 2720.440 ;
        RECT 2889.330 2720.380 2889.650 2720.440 ;
        RECT 2889.330 676.160 2889.650 676.220 ;
        RECT 2903.130 676.160 2903.450 676.220 ;
        RECT 2889.330 676.020 2903.450 676.160 ;
        RECT 2889.330 675.960 2889.650 676.020 ;
        RECT 2903.130 675.960 2903.450 676.020 ;
      LAYER via ;
        RECT 847.880 2723.440 848.140 2723.700 ;
        RECT 2889.360 2720.380 2889.620 2720.640 ;
        RECT 2889.360 675.960 2889.620 676.220 ;
        RECT 2903.160 675.960 2903.420 676.220 ;
      LAYER met2 ;
        RECT 846.510 2723.810 847.070 2731.680 ;
        RECT 846.510 2723.730 848.080 2723.810 ;
        RECT 846.510 2723.670 848.140 2723.730 ;
        RECT 846.510 2722.680 847.070 2723.670 ;
        RECT 847.880 2723.410 848.140 2723.670 ;
        RECT 2889.360 2720.350 2889.620 2720.670 ;
        RECT 2889.420 676.250 2889.560 2720.350 ;
        RECT 2889.360 675.930 2889.620 676.250 ;
        RECT 2903.160 675.930 2903.420 676.250 ;
        RECT 2903.220 674.405 2903.360 675.930 ;
        RECT 2903.150 674.035 2903.430 674.405 ;
      LAYER via2 ;
        RECT 2903.150 674.080 2903.430 674.360 ;
      LAYER met3 ;
        RECT 2903.125 674.370 2903.455 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2903.125 674.070 2924.800 674.370 ;
        RECT 2903.125 674.055 2903.455 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1932.550 2723.130 1932.830 2723.245 ;
        RECT 1933.030 2723.130 1933.590 2731.680 ;
        RECT 1932.550 2722.990 1933.590 2723.130 ;
        RECT 1932.550 2722.875 1932.830 2722.990 ;
        RECT 1933.030 2722.680 1933.590 2722.990 ;
        RECT 16.650 2714.715 16.930 2715.085 ;
        RECT 16.720 1544.125 16.860 2714.715 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 1932.550 2722.920 1932.830 2723.200 ;
        RECT 16.650 2714.760 16.930 2715.040 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 1932.525 2723.220 1932.855 2723.225 ;
        RECT 1932.270 2723.210 1932.855 2723.220 ;
        RECT 1932.070 2722.910 1932.855 2723.210 ;
        RECT 1932.270 2722.900 1932.855 2722.910 ;
        RECT 1932.525 2722.895 1932.855 2722.900 ;
        RECT 16.625 2715.050 16.955 2715.065 ;
        RECT 1156.710 2715.050 1157.090 2715.060 ;
        RECT 16.625 2714.750 1157.090 2715.050 ;
        RECT 16.625 2714.735 16.955 2714.750 ;
        RECT 1156.710 2714.740 1157.090 2714.750 ;
        RECT 1158.550 2715.050 1158.930 2715.060 ;
        RECT 1932.270 2715.050 1932.650 2715.060 ;
        RECT 1158.550 2714.750 1932.650 2715.050 ;
        RECT 1158.550 2714.740 1158.930 2714.750 ;
        RECT 1932.270 2714.740 1932.650 2714.750 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
      LAYER via3 ;
        RECT 1932.300 2722.900 1932.620 2723.220 ;
        RECT 1156.740 2714.740 1157.060 2715.060 ;
        RECT 1158.580 2714.740 1158.900 2715.060 ;
        RECT 1932.300 2714.740 1932.620 2715.060 ;
      LAYER met4 ;
        RECT 1932.295 2722.895 1932.625 2723.225 ;
        RECT 1932.310 2715.065 1932.610 2722.895 ;
        RECT 1156.735 2715.050 1157.065 2715.065 ;
        RECT 1158.575 2715.050 1158.905 2715.065 ;
        RECT 1156.735 2714.750 1158.905 2715.050 ;
        RECT 1156.735 2714.735 1157.065 2714.750 ;
        RECT 1158.575 2714.735 1158.905 2714.750 ;
        RECT 1932.295 2714.735 1932.625 2715.065 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.370 2741.320 25.690 2741.380 ;
        RECT 1971.630 2741.320 1971.950 2741.380 ;
        RECT 25.370 2741.180 1971.950 2741.320 ;
        RECT 25.370 2741.120 25.690 2741.180 ;
        RECT 1971.630 2741.120 1971.950 2741.180 ;
        RECT 13.870 1331.000 14.190 1331.060 ;
        RECT 25.370 1331.000 25.690 1331.060 ;
        RECT 13.870 1330.860 25.690 1331.000 ;
        RECT 13.870 1330.800 14.190 1330.860 ;
        RECT 25.370 1330.800 25.690 1330.860 ;
      LAYER via ;
        RECT 25.400 2741.120 25.660 2741.380 ;
        RECT 1971.660 2741.120 1971.920 2741.380 ;
        RECT 13.900 1330.800 14.160 1331.060 ;
        RECT 25.400 1330.800 25.660 1331.060 ;
      LAYER met2 ;
        RECT 25.400 2741.090 25.660 2741.410 ;
        RECT 1971.660 2741.090 1971.920 2741.410 ;
        RECT 25.460 1331.090 25.600 2741.090 ;
        RECT 1971.720 2731.680 1971.860 2741.090 ;
        RECT 1971.670 2722.680 1972.230 2731.680 ;
        RECT 13.900 1330.770 14.160 1331.090 ;
        RECT 25.400 1330.770 25.660 1331.090 ;
        RECT 13.960 1328.565 14.100 1330.770 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
      LAYER via2 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 748.490 2727.720 748.810 2727.780 ;
        RECT 2008.430 2727.720 2008.750 2727.780 ;
        RECT 748.490 2727.580 2008.750 2727.720 ;
        RECT 748.490 2727.520 748.810 2727.580 ;
        RECT 2008.430 2727.520 2008.750 2727.580 ;
        RECT 16.630 1117.820 16.950 1117.880 ;
        RECT 748.490 1117.820 748.810 1117.880 ;
        RECT 16.630 1117.680 748.810 1117.820 ;
        RECT 16.630 1117.620 16.950 1117.680 ;
        RECT 748.490 1117.620 748.810 1117.680 ;
      LAYER via ;
        RECT 748.520 2727.520 748.780 2727.780 ;
        RECT 2008.460 2727.520 2008.720 2727.780 ;
        RECT 16.660 1117.620 16.920 1117.880 ;
        RECT 748.520 1117.620 748.780 1117.880 ;
      LAYER met2 ;
        RECT 2010.310 2727.890 2010.870 2731.680 ;
        RECT 2008.520 2727.810 2010.870 2727.890 ;
        RECT 748.520 2727.490 748.780 2727.810 ;
        RECT 2008.460 2727.750 2010.870 2727.810 ;
        RECT 2008.460 2727.490 2008.720 2727.750 ;
        RECT 748.580 1117.910 748.720 2727.490 ;
        RECT 2010.310 2722.680 2010.870 2727.750 ;
        RECT 16.660 1117.590 16.920 1117.910 ;
        RECT 748.520 1117.590 748.780 1117.910 ;
        RECT 16.720 1113.005 16.860 1117.590 ;
        RECT 16.650 1112.635 16.930 1113.005 ;
      LAYER via2 ;
        RECT 16.650 1112.680 16.930 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 16.625 1112.970 16.955 1112.985 ;
        RECT -4.800 1112.670 16.955 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 16.625 1112.655 16.955 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.450 2739.620 24.770 2739.680 ;
        RECT 2049.370 2739.620 2049.690 2739.680 ;
        RECT 24.450 2739.480 2049.690 2739.620 ;
        RECT 24.450 2739.420 24.770 2739.480 ;
        RECT 2049.370 2739.420 2049.690 2739.480 ;
        RECT 13.870 897.500 14.190 897.560 ;
        RECT 24.450 897.500 24.770 897.560 ;
        RECT 13.870 897.360 24.770 897.500 ;
        RECT 13.870 897.300 14.190 897.360 ;
        RECT 24.450 897.300 24.770 897.360 ;
      LAYER via ;
        RECT 24.480 2739.420 24.740 2739.680 ;
        RECT 2049.400 2739.420 2049.660 2739.680 ;
        RECT 13.900 897.300 14.160 897.560 ;
        RECT 24.480 897.300 24.740 897.560 ;
      LAYER met2 ;
        RECT 24.480 2739.390 24.740 2739.710 ;
        RECT 2049.400 2739.390 2049.660 2739.710 ;
        RECT 24.540 897.590 24.680 2739.390 ;
        RECT 2049.460 2731.680 2049.600 2739.390 ;
        RECT 2049.410 2722.680 2049.970 2731.680 ;
        RECT 13.900 897.445 14.160 897.590 ;
        RECT 13.890 897.075 14.170 897.445 ;
        RECT 24.480 897.270 24.740 897.590 ;
      LAYER via2 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2086.705 2720.085 2086.875 2723.315 ;
      LAYER mcon ;
        RECT 2086.705 2723.145 2086.875 2723.315 ;
      LAYER met1 ;
        RECT 2086.630 2723.300 2086.950 2723.360 ;
        RECT 2086.435 2723.160 2086.950 2723.300 ;
        RECT 2086.630 2723.100 2086.950 2723.160 ;
        RECT 19.390 2720.240 19.710 2720.300 ;
        RECT 2086.645 2720.240 2086.935 2720.285 ;
        RECT 19.390 2720.100 2086.935 2720.240 ;
        RECT 19.390 2720.040 19.710 2720.100 ;
        RECT 2086.645 2720.055 2086.935 2720.100 ;
      LAYER via ;
        RECT 2086.660 2723.100 2086.920 2723.360 ;
        RECT 19.420 2720.040 19.680 2720.300 ;
      LAYER met2 ;
        RECT 2086.660 2723.130 2086.920 2723.390 ;
        RECT 2088.050 2723.130 2088.610 2731.680 ;
        RECT 2086.660 2723.070 2088.610 2723.130 ;
        RECT 2086.720 2722.990 2088.610 2723.070 ;
        RECT 2088.050 2722.680 2088.610 2722.990 ;
        RECT 19.420 2720.010 19.680 2720.330 ;
        RECT 19.480 681.885 19.620 2720.010 ;
        RECT 19.410 681.515 19.690 681.885 ;
      LAYER via2 ;
        RECT 19.410 681.560 19.690 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 19.385 681.850 19.715 681.865 ;
        RECT -4.800 681.550 19.715 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 19.385 681.535 19.715 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 2739.875 18.770 2740.245 ;
        RECT 2126.670 2739.875 2126.950 2740.245 ;
        RECT 18.560 466.325 18.700 2739.875 ;
        RECT 2126.740 2731.680 2126.880 2739.875 ;
        RECT 2126.690 2722.680 2127.250 2731.680 ;
        RECT 18.490 465.955 18.770 466.325 ;
      LAYER via2 ;
        RECT 18.490 2739.920 18.770 2740.200 ;
        RECT 2126.670 2739.920 2126.950 2740.200 ;
        RECT 18.490 466.000 18.770 466.280 ;
      LAYER met3 ;
        RECT 18.465 2740.210 18.795 2740.225 ;
        RECT 2126.645 2740.210 2126.975 2740.225 ;
        RECT 18.465 2739.910 2126.975 2740.210 ;
        RECT 18.465 2739.895 18.795 2739.910 ;
        RECT 2126.645 2739.895 2126.975 2739.910 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 18.465 466.290 18.795 466.305 ;
        RECT -4.800 465.990 18.795 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 18.465 465.975 18.795 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2163.985 2719.065 2164.155 2723.315 ;
      LAYER mcon ;
        RECT 2163.985 2723.145 2164.155 2723.315 ;
      LAYER met1 ;
        RECT 2163.910 2723.300 2164.230 2723.360 ;
        RECT 2163.715 2723.160 2164.230 2723.300 ;
        RECT 2163.910 2723.100 2164.230 2723.160 ;
        RECT 18.010 2719.220 18.330 2719.280 ;
        RECT 2163.925 2719.220 2164.215 2719.265 ;
        RECT 18.010 2719.080 2164.215 2719.220 ;
        RECT 18.010 2719.020 18.330 2719.080 ;
        RECT 2163.925 2719.035 2164.215 2719.080 ;
      LAYER via ;
        RECT 2163.940 2723.100 2164.200 2723.360 ;
        RECT 18.040 2719.020 18.300 2719.280 ;
      LAYER met2 ;
        RECT 2163.940 2723.130 2164.200 2723.390 ;
        RECT 2165.790 2723.130 2166.350 2731.680 ;
        RECT 2163.940 2723.070 2166.350 2723.130 ;
        RECT 2164.000 2722.990 2166.350 2723.070 ;
        RECT 2165.790 2722.680 2166.350 2722.990 ;
        RECT 18.040 2718.990 18.300 2719.310 ;
        RECT 18.100 250.765 18.240 2718.990 ;
        RECT 18.030 250.395 18.310 250.765 ;
      LAYER via2 ;
        RECT 18.030 250.440 18.310 250.720 ;
      LAYER met3 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 18.005 250.730 18.335 250.745 ;
        RECT -4.800 250.430 18.335 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 18.005 250.415 18.335 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 41.040 14.190 41.100 ;
        RECT 23.990 41.040 24.310 41.100 ;
        RECT 13.870 40.900 24.310 41.040 ;
        RECT 13.870 40.840 14.190 40.900 ;
        RECT 23.990 40.840 24.310 40.900 ;
      LAYER via ;
        RECT 13.900 40.840 14.160 41.100 ;
        RECT 24.020 40.840 24.280 41.100 ;
      LAYER met2 ;
        RECT 24.010 2745.995 24.290 2746.365 ;
        RECT 2204.410 2745.995 2204.690 2746.365 ;
        RECT 24.080 41.130 24.220 2745.995 ;
        RECT 2204.480 2731.680 2204.620 2745.995 ;
        RECT 2204.430 2722.680 2204.990 2731.680 ;
        RECT 13.900 40.810 14.160 41.130 ;
        RECT 24.020 40.810 24.280 41.130 ;
        RECT 13.960 35.885 14.100 40.810 ;
        RECT 13.890 35.515 14.170 35.885 ;
      LAYER via2 ;
        RECT 24.010 2746.040 24.290 2746.320 ;
        RECT 2204.410 2746.040 2204.690 2746.320 ;
        RECT 13.890 35.560 14.170 35.840 ;
      LAYER met3 ;
        RECT 23.985 2746.330 24.315 2746.345 ;
        RECT 2204.385 2746.330 2204.715 2746.345 ;
        RECT 23.985 2746.030 2204.715 2746.330 ;
        RECT 23.985 2746.015 24.315 2746.030 ;
        RECT 2204.385 2746.015 2204.715 2746.030 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 13.865 35.850 14.195 35.865 ;
        RECT -4.800 35.550 14.195 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 13.865 35.535 14.195 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 887.410 2727.040 887.730 2727.100 ;
        RECT 2245.790 2727.040 2246.110 2727.100 ;
        RECT 887.410 2726.900 2246.110 2727.040 ;
        RECT 887.410 2726.840 887.730 2726.900 ;
        RECT 2245.790 2726.840 2246.110 2726.900 ;
        RECT 2245.790 910.760 2246.110 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2245.790 910.620 2901.150 910.760 ;
        RECT 2245.790 910.560 2246.110 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 887.440 2726.840 887.700 2727.100 ;
        RECT 2245.820 2726.840 2246.080 2727.100 ;
        RECT 2245.820 910.560 2246.080 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 885.610 2727.210 886.170 2731.680 ;
        RECT 885.610 2727.130 887.640 2727.210 ;
        RECT 885.610 2727.070 887.700 2727.130 ;
        RECT 885.610 2722.680 886.170 2727.070 ;
        RECT 887.440 2726.810 887.700 2727.070 ;
        RECT 2245.820 2726.810 2246.080 2727.130 ;
        RECT 2245.880 910.850 2246.020 2726.810 ;
        RECT 2245.820 910.530 2246.080 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 923.750 2727.380 924.070 2727.440 ;
        RECT 2246.250 2727.380 2246.570 2727.440 ;
        RECT 923.750 2727.240 2246.570 2727.380 ;
        RECT 923.750 2727.180 924.070 2727.240 ;
        RECT 2246.250 2727.180 2246.570 2727.240 ;
        RECT 2246.250 1145.360 2246.570 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2246.250 1145.220 2901.150 1145.360 ;
        RECT 2246.250 1145.160 2246.570 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 923.780 2727.180 924.040 2727.440 ;
        RECT 2246.280 2727.180 2246.540 2727.440 ;
        RECT 2246.280 1145.160 2246.540 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 923.780 2727.210 924.040 2727.470 ;
        RECT 924.250 2727.210 924.810 2731.680 ;
        RECT 923.780 2727.150 924.810 2727.210 ;
        RECT 2246.280 2727.150 2246.540 2727.470 ;
        RECT 923.840 2727.070 924.810 2727.150 ;
        RECT 924.250 2722.680 924.810 2727.070 ;
        RECT 2246.340 1145.450 2246.480 2727.150 ;
        RECT 2246.280 1145.130 2246.540 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 964.230 2726.020 964.550 2726.080 ;
        RECT 2903.590 2726.020 2903.910 2726.080 ;
        RECT 964.230 2725.880 2903.910 2726.020 ;
        RECT 964.230 2725.820 964.550 2725.880 ;
        RECT 2903.590 2725.820 2903.910 2725.880 ;
      LAYER via ;
        RECT 964.260 2725.820 964.520 2726.080 ;
        RECT 2903.620 2725.820 2903.880 2726.080 ;
      LAYER met2 ;
        RECT 962.890 2725.850 963.450 2731.680 ;
        RECT 964.260 2725.850 964.520 2726.110 ;
        RECT 962.890 2725.790 964.520 2725.850 ;
        RECT 2903.620 2725.790 2903.880 2726.110 ;
        RECT 962.890 2725.710 964.460 2725.790 ;
        RECT 962.890 2722.680 963.450 2725.710 ;
        RECT 2903.680 1378.885 2903.820 2725.790 ;
        RECT 2903.610 1378.515 2903.890 1378.885 ;
      LAYER via2 ;
        RECT 2903.610 1378.560 2903.890 1378.840 ;
      LAYER met3 ;
        RECT 2903.585 1378.850 2903.915 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2903.585 1378.550 2924.800 1378.850 ;
        RECT 2903.585 1378.535 2903.915 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1003.405 2722.805 1003.575 2723.655 ;
      LAYER mcon ;
        RECT 1003.405 2723.485 1003.575 2723.655 ;
      LAYER met1 ;
        RECT 1003.330 2723.640 1003.650 2723.700 ;
        RECT 1003.135 2723.500 1003.650 2723.640 ;
        RECT 1003.330 2723.440 1003.650 2723.500 ;
        RECT 1003.345 2722.960 1003.635 2723.005 ;
        RECT 2904.510 2722.960 2904.830 2723.020 ;
        RECT 1003.345 2722.820 2904.830 2722.960 ;
        RECT 1003.345 2722.775 1003.635 2722.820 ;
        RECT 2904.510 2722.760 2904.830 2722.820 ;
      LAYER via ;
        RECT 1003.360 2723.440 1003.620 2723.700 ;
        RECT 2904.540 2722.760 2904.800 2723.020 ;
      LAYER met2 ;
        RECT 1001.990 2723.810 1002.550 2731.680 ;
        RECT 1001.990 2723.730 1003.560 2723.810 ;
        RECT 1001.990 2723.670 1003.620 2723.730 ;
        RECT 1001.990 2722.680 1002.550 2723.670 ;
        RECT 1003.360 2723.410 1003.620 2723.670 ;
        RECT 2904.540 2722.730 2904.800 2723.050 ;
        RECT 2904.600 1613.485 2904.740 2722.730 ;
        RECT 2904.530 1613.115 2904.810 1613.485 ;
      LAYER via2 ;
        RECT 2904.530 1613.160 2904.810 1613.440 ;
      LAYER met3 ;
        RECT 2904.505 1613.450 2904.835 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2904.505 1613.150 2924.800 1613.450 ;
        RECT 2904.505 1613.135 2904.835 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1040.150 2723.130 1040.430 2723.245 ;
        RECT 1040.630 2723.130 1041.190 2731.680 ;
        RECT 1040.150 2722.990 1041.190 2723.130 ;
        RECT 1040.150 2722.875 1040.430 2722.990 ;
        RECT 1040.630 2722.680 1041.190 2722.990 ;
        RECT 2899.930 2716.755 2900.210 2717.125 ;
        RECT 2900.000 1848.085 2900.140 2716.755 ;
        RECT 2899.930 1847.715 2900.210 1848.085 ;
      LAYER via2 ;
        RECT 1040.150 2722.920 1040.430 2723.200 ;
        RECT 2899.930 2716.800 2900.210 2717.080 ;
        RECT 2899.930 1847.760 2900.210 1848.040 ;
      LAYER met3 ;
        RECT 1040.125 2723.210 1040.455 2723.225 ;
        RECT 1040.790 2723.210 1041.170 2723.220 ;
        RECT 1040.125 2722.910 1041.170 2723.210 ;
        RECT 1040.125 2722.895 1040.455 2722.910 ;
        RECT 1040.790 2722.900 1041.170 2722.910 ;
        RECT 1040.790 2717.090 1041.170 2717.100 ;
        RECT 2899.905 2717.090 2900.235 2717.105 ;
        RECT 1040.790 2716.790 2900.235 2717.090 ;
        RECT 1040.790 2716.780 1041.170 2716.790 ;
        RECT 2899.905 2716.775 2900.235 2716.790 ;
        RECT 2899.905 1848.050 2900.235 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2899.905 1847.750 2924.800 1848.050 ;
        RECT 2899.905 1847.735 2900.235 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
      LAYER via3 ;
        RECT 1040.820 2722.900 1041.140 2723.220 ;
        RECT 1040.820 2716.780 1041.140 2717.100 ;
      LAYER met4 ;
        RECT 1040.815 2722.895 1041.145 2723.225 ;
        RECT 1040.830 2717.105 1041.130 2722.895 ;
        RECT 1040.815 2716.775 1041.145 2717.105 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1080.610 2723.980 1080.930 2724.040 ;
        RECT 2247.170 2723.980 2247.490 2724.040 ;
        RECT 1080.610 2723.840 2247.490 2723.980 ;
        RECT 1080.610 2723.780 1080.930 2723.840 ;
        RECT 2247.170 2723.780 2247.490 2723.840 ;
        RECT 2247.170 2083.760 2247.490 2083.820 ;
        RECT 2900.370 2083.760 2900.690 2083.820 ;
        RECT 2247.170 2083.620 2900.690 2083.760 ;
        RECT 2247.170 2083.560 2247.490 2083.620 ;
        RECT 2900.370 2083.560 2900.690 2083.620 ;
      LAYER via ;
        RECT 1080.640 2723.780 1080.900 2724.040 ;
        RECT 2247.200 2723.780 2247.460 2724.040 ;
        RECT 2247.200 2083.560 2247.460 2083.820 ;
        RECT 2900.400 2083.560 2900.660 2083.820 ;
      LAYER met2 ;
        RECT 1079.270 2723.810 1079.830 2731.680 ;
        RECT 1080.640 2723.810 1080.900 2724.070 ;
        RECT 1079.270 2723.750 1080.900 2723.810 ;
        RECT 2247.200 2723.750 2247.460 2724.070 ;
        RECT 1079.270 2723.670 1080.840 2723.750 ;
        RECT 1079.270 2722.680 1079.830 2723.670 ;
        RECT 2247.260 2083.850 2247.400 2723.750 ;
        RECT 2247.200 2083.530 2247.460 2083.850 ;
        RECT 2900.400 2083.530 2900.660 2083.850 ;
        RECT 2900.460 2082.685 2900.600 2083.530 ;
        RECT 2900.390 2082.315 2900.670 2082.685 ;
      LAYER via2 ;
        RECT 2900.390 2082.360 2900.670 2082.640 ;
      LAYER met3 ;
        RECT 2900.365 2082.650 2900.695 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.365 2082.350 2924.800 2082.650 ;
        RECT 2900.365 2082.335 2900.695 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1118.330 2745.740 1118.650 2745.800 ;
        RECT 2248.090 2745.740 2248.410 2745.800 ;
        RECT 1118.330 2745.600 2248.410 2745.740 ;
        RECT 1118.330 2745.540 1118.650 2745.600 ;
        RECT 2248.090 2745.540 2248.410 2745.600 ;
        RECT 2248.090 2318.360 2248.410 2318.420 ;
        RECT 2900.370 2318.360 2900.690 2318.420 ;
        RECT 2248.090 2318.220 2900.690 2318.360 ;
        RECT 2248.090 2318.160 2248.410 2318.220 ;
        RECT 2900.370 2318.160 2900.690 2318.220 ;
      LAYER via ;
        RECT 1118.360 2745.540 1118.620 2745.800 ;
        RECT 2248.120 2745.540 2248.380 2745.800 ;
        RECT 2248.120 2318.160 2248.380 2318.420 ;
        RECT 2900.400 2318.160 2900.660 2318.420 ;
      LAYER met2 ;
        RECT 1118.360 2745.510 1118.620 2745.830 ;
        RECT 2248.120 2745.510 2248.380 2745.830 ;
        RECT 1118.420 2731.680 1118.560 2745.510 ;
        RECT 1118.370 2722.680 1118.930 2731.680 ;
        RECT 2248.180 2318.450 2248.320 2745.510 ;
        RECT 2248.120 2318.130 2248.380 2318.450 ;
        RECT 2900.400 2318.130 2900.660 2318.450 ;
        RECT 2900.460 2317.285 2900.600 2318.130 ;
        RECT 2900.390 2316.915 2900.670 2317.285 ;
      LAYER via2 ;
        RECT 2900.390 2316.960 2900.670 2317.240 ;
      LAYER met3 ;
        RECT 2900.365 2317.250 2900.695 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.365 2316.950 2924.800 2317.250 ;
        RECT 2900.365 2316.935 2900.695 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 782.070 2760.360 782.390 2760.420 ;
        RECT 2887.490 2760.360 2887.810 2760.420 ;
        RECT 782.070 2760.220 2887.810 2760.360 ;
        RECT 782.070 2760.160 782.390 2760.220 ;
        RECT 2887.490 2760.160 2887.810 2760.220 ;
        RECT 2887.490 151.540 2887.810 151.600 ;
        RECT 2898.070 151.540 2898.390 151.600 ;
        RECT 2887.490 151.400 2898.390 151.540 ;
        RECT 2887.490 151.340 2887.810 151.400 ;
        RECT 2898.070 151.340 2898.390 151.400 ;
      LAYER via ;
        RECT 782.100 2760.160 782.360 2760.420 ;
        RECT 2887.520 2760.160 2887.780 2760.420 ;
        RECT 2887.520 151.340 2887.780 151.600 ;
        RECT 2898.100 151.340 2898.360 151.600 ;
      LAYER met2 ;
        RECT 782.100 2760.130 782.360 2760.450 ;
        RECT 2887.520 2760.130 2887.780 2760.450 ;
        RECT 782.160 2731.680 782.300 2760.130 ;
        RECT 782.110 2722.680 782.670 2731.680 ;
        RECT 2887.580 151.630 2887.720 2760.130 ;
        RECT 2887.520 151.310 2887.780 151.630 ;
        RECT 2898.100 151.310 2898.360 151.630 ;
        RECT 2898.160 146.725 2898.300 151.310 ;
        RECT 2898.090 146.355 2898.370 146.725 ;
      LAYER via2 ;
        RECT 2898.090 146.400 2898.370 146.680 ;
      LAYER met3 ;
        RECT 2898.065 146.690 2898.395 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2898.065 146.390 2924.800 146.690 ;
        RECT 2898.065 146.375 2898.395 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1171.690 2723.640 1172.010 2723.700 ;
        RECT 2900.370 2723.640 2900.690 2723.700 ;
        RECT 1171.690 2723.500 2900.690 2723.640 ;
        RECT 1171.690 2723.440 1172.010 2723.500 ;
        RECT 2900.370 2723.440 2900.690 2723.500 ;
      LAYER via ;
        RECT 1171.720 2723.440 1171.980 2723.700 ;
        RECT 2900.400 2723.440 2900.660 2723.700 ;
      LAYER met2 ;
        RECT 1169.890 2723.810 1170.450 2731.680 ;
        RECT 1169.890 2723.730 1171.920 2723.810 ;
        RECT 1169.890 2723.670 1171.980 2723.730 ;
        RECT 1169.890 2722.680 1170.450 2723.670 ;
        RECT 1171.720 2723.410 1171.980 2723.670 ;
        RECT 2900.400 2723.410 2900.660 2723.730 ;
        RECT 2900.460 2493.405 2900.600 2723.410 ;
        RECT 2900.390 2493.035 2900.670 2493.405 ;
      LAYER via2 ;
        RECT 2900.390 2493.080 2900.670 2493.360 ;
      LAYER met3 ;
        RECT 2900.365 2493.370 2900.695 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.365 2493.070 2924.800 2493.370 ;
        RECT 2900.365 2493.055 2900.695 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.330 2726.700 1210.650 2726.760 ;
        RECT 2900.830 2726.700 2901.150 2726.760 ;
        RECT 1210.330 2726.560 2901.150 2726.700 ;
        RECT 1210.330 2726.500 1210.650 2726.560 ;
        RECT 2900.830 2726.500 2901.150 2726.560 ;
      LAYER via ;
        RECT 1210.360 2726.500 1210.620 2726.760 ;
        RECT 2900.860 2726.500 2901.120 2726.760 ;
      LAYER met2 ;
        RECT 1208.530 2726.530 1209.090 2731.680 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2726.790 2901.060 2727.635 ;
        RECT 1210.360 2726.530 1210.620 2726.790 ;
        RECT 1208.530 2726.470 1210.620 2726.530 ;
        RECT 2900.860 2726.470 2901.120 2726.790 ;
        RECT 1208.530 2726.390 1210.560 2726.470 ;
        RECT 1208.530 2722.680 1209.090 2726.390 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 2960.280 1248.830 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1248.510 2960.140 2901.150 2960.280 ;
        RECT 1248.510 2960.080 1248.830 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 1248.540 2960.080 1248.800 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1248.540 2960.050 1248.800 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1247.630 2731.290 1248.190 2731.680 ;
        RECT 1248.600 2731.290 1248.740 2960.050 ;
        RECT 1247.630 2731.150 1248.740 2731.290 ;
        RECT 1247.630 2722.680 1248.190 2731.150 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1289.910 3194.880 1290.230 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1289.910 3194.740 2901.150 3194.880 ;
        RECT 1289.910 3194.680 1290.230 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 1289.940 3194.680 1290.200 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1289.940 3194.650 1290.200 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 1290.000 2731.970 1290.140 3194.650 ;
        RECT 1288.160 2731.830 1290.140 2731.970 ;
        RECT 1286.270 2731.290 1286.830 2731.680 ;
        RECT 1288.160 2731.290 1288.300 2731.830 ;
        RECT 1286.270 2731.150 1288.300 2731.290 ;
        RECT 1286.270 2722.680 1286.830 2731.150 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 1331.310 3429.480 1331.630 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 1331.310 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1506.200 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2149.740 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1331.310 3429.280 1331.630 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1331.340 3429.280 1331.600 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1331.340 3429.250 1331.600 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1331.400 2731.970 1331.540 3429.250 ;
        RECT 1327.260 2731.830 1331.540 2731.970 ;
        RECT 1324.910 2730.610 1325.470 2731.680 ;
        RECT 1327.260 2730.610 1327.400 2731.830 ;
        RECT 1324.910 2730.470 1327.400 2730.610 ;
        RECT 1324.910 2722.680 1325.470 2730.470 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1365.810 3502.240 1366.130 3502.300 ;
        RECT 2717.290 3502.240 2717.610 3502.300 ;
        RECT 1365.810 3502.100 2717.610 3502.240 ;
        RECT 1365.810 3502.040 1366.130 3502.100 ;
        RECT 2717.290 3502.040 2717.610 3502.100 ;
      LAYER via ;
        RECT 1365.840 3502.040 1366.100 3502.300 ;
        RECT 2717.320 3502.040 2717.580 3502.300 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3502.330 2717.520 3517.600 ;
        RECT 1365.840 3502.010 1366.100 3502.330 ;
        RECT 2717.320 3502.010 2717.580 3502.330 ;
        RECT 1364.010 2731.290 1364.570 2731.680 ;
        RECT 1365.900 2731.290 1366.040 3502.010 ;
        RECT 1364.010 2731.150 1366.040 2731.290 ;
        RECT 1364.010 2722.680 1364.570 2731.150 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 3503.940 1407.530 3504.000 ;
        RECT 2392.530 3503.940 2392.850 3504.000 ;
        RECT 1407.210 3503.800 2392.850 3503.940 ;
        RECT 1407.210 3503.740 1407.530 3503.800 ;
        RECT 2392.530 3503.740 2392.850 3503.800 ;
      LAYER via ;
        RECT 1407.240 3503.740 1407.500 3504.000 ;
        RECT 2392.560 3503.740 2392.820 3504.000 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3504.030 2392.760 3517.600 ;
        RECT 1407.240 3503.710 1407.500 3504.030 ;
        RECT 2392.560 3503.710 2392.820 3504.030 ;
        RECT 1407.300 2731.970 1407.440 3503.710 ;
        RECT 1405.920 2731.830 1407.440 2731.970 ;
        RECT 1402.650 2731.290 1403.210 2731.680 ;
        RECT 1405.920 2731.290 1406.060 2731.830 ;
        RECT 1402.650 2731.150 1406.060 2731.290 ;
        RECT 1402.650 2722.680 1403.210 2731.150 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 3500.880 1442.030 3500.940 ;
        RECT 2068.230 3500.880 2068.550 3500.940 ;
        RECT 1441.710 3500.740 2068.550 3500.880 ;
        RECT 1441.710 3500.680 1442.030 3500.740 ;
        RECT 2068.230 3500.680 2068.550 3500.740 ;
      LAYER via ;
        RECT 1441.740 3500.680 1442.000 3500.940 ;
        RECT 2068.260 3500.680 2068.520 3500.940 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3500.970 2068.460 3517.600 ;
        RECT 1441.740 3500.650 1442.000 3500.970 ;
        RECT 2068.260 3500.650 2068.520 3500.970 ;
        RECT 1441.800 2731.680 1441.940 3500.650 ;
        RECT 1441.290 2731.150 1441.940 2731.680 ;
        RECT 1441.290 2722.680 1441.850 2731.150 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1483.110 3499.520 1483.430 3499.580 ;
        RECT 1743.930 3499.520 1744.250 3499.580 ;
        RECT 1483.110 3499.380 1744.250 3499.520 ;
        RECT 1483.110 3499.320 1483.430 3499.380 ;
        RECT 1743.930 3499.320 1744.250 3499.380 ;
      LAYER via ;
        RECT 1483.140 3499.320 1483.400 3499.580 ;
        RECT 1743.960 3499.320 1744.220 3499.580 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3499.610 1744.160 3517.600 ;
        RECT 1483.140 3499.290 1483.400 3499.610 ;
        RECT 1743.960 3499.290 1744.220 3499.610 ;
        RECT 1480.390 2730.610 1480.950 2731.680 ;
        RECT 1483.200 2730.610 1483.340 3499.290 ;
        RECT 1480.390 2730.470 1483.340 2730.610 ;
        RECT 1480.390 2722.680 1480.950 2730.470 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3498.500 1419.490 3498.560 ;
        RECT 1518.070 3498.500 1518.390 3498.560 ;
        RECT 1419.170 3498.360 1518.390 3498.500 ;
        RECT 1419.170 3498.300 1419.490 3498.360 ;
        RECT 1518.070 3498.300 1518.390 3498.360 ;
      LAYER via ;
        RECT 1419.200 3498.300 1419.460 3498.560 ;
        RECT 1518.100 3498.300 1518.360 3498.560 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3498.590 1419.400 3517.600 ;
        RECT 1419.200 3498.270 1419.460 3498.590 ;
        RECT 1518.100 3498.270 1518.360 3498.590 ;
        RECT 1518.160 2731.290 1518.300 3498.270 ;
        RECT 1519.030 2731.290 1519.590 2731.680 ;
        RECT 1518.160 2731.150 1519.590 2731.290 ;
        RECT 1519.030 2722.680 1519.590 2731.150 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 820.325 2719.745 820.495 2723.655 ;
      LAYER mcon ;
        RECT 820.325 2723.485 820.495 2723.655 ;
      LAYER met1 ;
        RECT 820.250 2723.640 820.570 2723.700 ;
        RECT 820.055 2723.500 820.570 2723.640 ;
        RECT 820.250 2723.440 820.570 2723.500 ;
        RECT 820.265 2719.900 820.555 2719.945 ;
        RECT 2888.410 2719.900 2888.730 2719.960 ;
        RECT 820.265 2719.760 2888.730 2719.900 ;
        RECT 820.265 2719.715 820.555 2719.760 ;
        RECT 2888.410 2719.700 2888.730 2719.760 ;
        RECT 2888.410 386.140 2888.730 386.200 ;
        RECT 2898.070 386.140 2898.390 386.200 ;
        RECT 2888.410 386.000 2898.390 386.140 ;
        RECT 2888.410 385.940 2888.730 386.000 ;
        RECT 2898.070 385.940 2898.390 386.000 ;
      LAYER via ;
        RECT 820.280 2723.440 820.540 2723.700 ;
        RECT 2888.440 2719.700 2888.700 2719.960 ;
        RECT 2888.440 385.940 2888.700 386.200 ;
        RECT 2898.100 385.940 2898.360 386.200 ;
      LAYER met2 ;
        RECT 820.750 2723.810 821.310 2731.680 ;
        RECT 820.340 2723.730 821.310 2723.810 ;
        RECT 820.280 2723.670 821.310 2723.730 ;
        RECT 820.280 2723.410 820.540 2723.670 ;
        RECT 820.750 2722.680 821.310 2723.670 ;
        RECT 2888.440 2719.670 2888.700 2719.990 ;
        RECT 2888.500 386.230 2888.640 2719.670 ;
        RECT 2888.440 385.910 2888.700 386.230 ;
        RECT 2898.100 385.910 2898.360 386.230 ;
        RECT 2898.160 381.325 2898.300 385.910 ;
        RECT 2898.090 380.955 2898.370 381.325 ;
      LAYER via2 ;
        RECT 2898.090 381.000 2898.370 381.280 ;
      LAYER met3 ;
        RECT 2898.065 381.290 2898.395 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2898.065 380.990 2924.800 381.290 ;
        RECT 2898.065 380.975 2898.395 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3499.860 1095.190 3499.920 ;
        RECT 1552.570 3499.860 1552.890 3499.920 ;
        RECT 1094.870 3499.720 1552.890 3499.860 ;
        RECT 1094.870 3499.660 1095.190 3499.720 ;
        RECT 1552.570 3499.660 1552.890 3499.720 ;
      LAYER via ;
        RECT 1094.900 3499.660 1095.160 3499.920 ;
        RECT 1552.600 3499.660 1552.860 3499.920 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3499.950 1095.100 3517.600 ;
        RECT 1094.900 3499.630 1095.160 3499.950 ;
        RECT 1552.600 3499.630 1552.860 3499.950 ;
        RECT 1552.660 2731.970 1552.800 3499.630 ;
        RECT 1552.660 2731.830 1555.560 2731.970 ;
        RECT 1555.420 2731.290 1555.560 2731.830 ;
        RECT 1557.670 2731.290 1558.230 2731.680 ;
        RECT 1555.420 2731.150 1558.230 2731.290 ;
        RECT 1557.670 2722.680 1558.230 2731.150 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.960 770.890 3505.020 ;
        RECT 1593.970 3504.960 1594.290 3505.020 ;
        RECT 770.570 3504.820 1594.290 3504.960 ;
        RECT 770.570 3504.760 770.890 3504.820 ;
        RECT 1593.970 3504.760 1594.290 3504.820 ;
      LAYER via ;
        RECT 770.600 3504.760 770.860 3505.020 ;
        RECT 1594.000 3504.760 1594.260 3505.020 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3505.050 770.800 3517.600 ;
        RECT 770.600 3504.730 770.860 3505.050 ;
        RECT 1594.000 3504.730 1594.260 3505.050 ;
        RECT 1594.060 2731.290 1594.200 3504.730 ;
        RECT 1596.770 2731.290 1597.330 2731.680 ;
        RECT 1594.060 2731.150 1597.330 2731.290 ;
        RECT 1596.770 2722.680 1597.330 2731.150 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3503.260 446.130 3503.320 ;
        RECT 1635.370 3503.260 1635.690 3503.320 ;
        RECT 445.810 3503.120 1635.690 3503.260 ;
        RECT 445.810 3503.060 446.130 3503.120 ;
        RECT 1635.370 3503.060 1635.690 3503.120 ;
      LAYER via ;
        RECT 445.840 3503.060 446.100 3503.320 ;
        RECT 1635.400 3503.060 1635.660 3503.320 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.350 446.040 3517.600 ;
        RECT 445.840 3503.030 446.100 3503.350 ;
        RECT 1635.400 3503.030 1635.660 3503.350 ;
        RECT 1635.460 2731.680 1635.600 3503.030 ;
        RECT 1635.410 2722.680 1635.970 2731.680 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1669.870 3501.560 1670.190 3501.620 ;
        RECT 121.510 3501.420 1670.190 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1669.870 3501.360 1670.190 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1669.900 3501.360 1670.160 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1669.900 3501.330 1670.160 3501.650 ;
        RECT 1669.960 2731.970 1670.100 3501.330 ;
        RECT 1669.960 2731.830 1672.400 2731.970 ;
        RECT 1672.260 2731.290 1672.400 2731.830 ;
        RECT 1674.050 2731.290 1674.610 2731.680 ;
        RECT 1672.260 2731.150 1674.610 2731.290 ;
        RECT 1674.050 2722.680 1674.610 2731.150 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1711.270 3339.720 1711.590 3339.780 ;
        RECT 17.090 3339.580 1711.590 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1711.270 3339.520 1711.590 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1711.300 3339.520 1711.560 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1711.300 3339.490 1711.560 3339.810 ;
        RECT 1711.360 2731.290 1711.500 3339.490 ;
        RECT 1713.150 2731.290 1713.710 2731.680 ;
        RECT 1711.360 2731.150 1713.710 2731.290 ;
        RECT 1713.150 2722.680 1713.710 2731.150 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 1745.770 3050.040 1746.090 3050.100 ;
        RECT 17.090 3049.900 1746.090 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 1745.770 3049.840 1746.090 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 1745.800 3049.840 1746.060 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 1745.800 3049.810 1746.060 3050.130 ;
        RECT 1745.860 2731.970 1746.000 3049.810 ;
        RECT 1745.860 2731.830 1748.760 2731.970 ;
        RECT 1748.620 2731.290 1748.760 2731.830 ;
        RECT 1751.790 2731.290 1752.350 2731.680 ;
        RECT 1748.620 2731.150 1752.350 2731.290 ;
        RECT 1751.790 2722.680 1752.350 2731.150 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2760.700 17.410 2760.760 ;
        RECT 1787.170 2760.700 1787.490 2760.760 ;
        RECT 17.090 2760.560 1787.490 2760.700 ;
        RECT 17.090 2760.500 17.410 2760.560 ;
        RECT 1787.170 2760.500 1787.490 2760.560 ;
      LAYER via ;
        RECT 17.120 2760.500 17.380 2760.760 ;
        RECT 1787.200 2760.500 1787.460 2760.760 ;
      LAYER met2 ;
        RECT 17.110 2765.035 17.390 2765.405 ;
        RECT 17.180 2760.790 17.320 2765.035 ;
        RECT 17.120 2760.470 17.380 2760.790 ;
        RECT 1787.200 2760.470 1787.460 2760.790 ;
        RECT 1787.260 2731.290 1787.400 2760.470 ;
        RECT 1790.430 2731.290 1790.990 2731.680 ;
        RECT 1787.260 2731.150 1790.990 2731.290 ;
        RECT 1790.430 2722.680 1790.990 2731.150 ;
      LAYER via2 ;
        RECT 17.110 2765.080 17.390 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 17.085 2765.370 17.415 2765.385 ;
        RECT -4.800 2765.070 17.415 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 17.085 2765.055 17.415 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.530 2744.720 23.850 2744.780 ;
        RECT 1829.490 2744.720 1829.810 2744.780 ;
        RECT 23.530 2744.580 1829.810 2744.720 ;
        RECT 23.530 2744.520 23.850 2744.580 ;
        RECT 1829.490 2744.520 1829.810 2744.580 ;
        RECT 13.870 2477.820 14.190 2477.880 ;
        RECT 23.530 2477.820 23.850 2477.880 ;
        RECT 13.870 2477.680 23.850 2477.820 ;
        RECT 13.870 2477.620 14.190 2477.680 ;
        RECT 23.530 2477.620 23.850 2477.680 ;
      LAYER via ;
        RECT 23.560 2744.520 23.820 2744.780 ;
        RECT 1829.520 2744.520 1829.780 2744.780 ;
        RECT 13.900 2477.620 14.160 2477.880 ;
        RECT 23.560 2477.620 23.820 2477.880 ;
      LAYER met2 ;
        RECT 23.560 2744.490 23.820 2744.810 ;
        RECT 1829.520 2744.490 1829.780 2744.810 ;
        RECT 23.620 2477.910 23.760 2744.490 ;
        RECT 1829.580 2731.680 1829.720 2744.490 ;
        RECT 1829.530 2722.680 1830.090 2731.680 ;
        RECT 13.900 2477.765 14.160 2477.910 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
        RECT 23.560 2477.590 23.820 2477.910 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 2743.700 27.070 2743.760 ;
        RECT 1868.130 2743.700 1868.450 2743.760 ;
        RECT 26.750 2743.560 1868.450 2743.700 ;
        RECT 26.750 2743.500 27.070 2743.560 ;
        RECT 1868.130 2743.500 1868.450 2743.560 ;
        RECT 13.870 2192.900 14.190 2192.960 ;
        RECT 26.750 2192.900 27.070 2192.960 ;
        RECT 13.870 2192.760 27.070 2192.900 ;
        RECT 13.870 2192.700 14.190 2192.760 ;
        RECT 26.750 2192.700 27.070 2192.760 ;
      LAYER via ;
        RECT 26.780 2743.500 27.040 2743.760 ;
        RECT 1868.160 2743.500 1868.420 2743.760 ;
        RECT 13.900 2192.700 14.160 2192.960 ;
        RECT 26.780 2192.700 27.040 2192.960 ;
      LAYER met2 ;
        RECT 26.780 2743.470 27.040 2743.790 ;
        RECT 1868.160 2743.470 1868.420 2743.790 ;
        RECT 26.840 2192.990 26.980 2743.470 ;
        RECT 1868.220 2731.680 1868.360 2743.470 ;
        RECT 1868.170 2722.680 1868.730 2731.680 ;
        RECT 13.900 2192.670 14.160 2192.990 ;
        RECT 26.780 2192.670 27.040 2192.990 ;
        RECT 13.960 2190.125 14.100 2192.670 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
      LAYER via2 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.810 2742.680 32.130 2742.740 ;
        RECT 1906.770 2742.680 1907.090 2742.740 ;
        RECT 31.810 2742.540 1907.090 2742.680 ;
        RECT 31.810 2742.480 32.130 2742.540 ;
        RECT 1906.770 2742.480 1907.090 2742.540 ;
        RECT 14.790 1903.220 15.110 1903.280 ;
        RECT 31.810 1903.220 32.130 1903.280 ;
        RECT 14.790 1903.080 32.130 1903.220 ;
        RECT 14.790 1903.020 15.110 1903.080 ;
        RECT 31.810 1903.020 32.130 1903.080 ;
      LAYER via ;
        RECT 31.840 2742.480 32.100 2742.740 ;
        RECT 1906.800 2742.480 1907.060 2742.740 ;
        RECT 14.820 1903.020 15.080 1903.280 ;
        RECT 31.840 1903.020 32.100 1903.280 ;
      LAYER met2 ;
        RECT 31.840 2742.450 32.100 2742.770 ;
        RECT 1906.800 2742.450 1907.060 2742.770 ;
        RECT 31.900 1903.310 32.040 2742.450 ;
        RECT 1906.860 2731.680 1907.000 2742.450 ;
        RECT 1906.810 2722.680 1907.370 2731.680 ;
        RECT 14.820 1903.165 15.080 1903.310 ;
        RECT 14.810 1902.795 15.090 1903.165 ;
        RECT 31.840 1902.990 32.100 1903.310 ;
      LAYER via2 ;
        RECT 14.810 1902.840 15.090 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 14.785 1903.130 15.115 1903.145 ;
        RECT -4.800 1902.830 15.115 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 14.785 1902.815 15.115 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 860.805 2720.765 860.975 2723.655 ;
      LAYER mcon ;
        RECT 860.805 2723.485 860.975 2723.655 ;
      LAYER met1 ;
        RECT 860.730 2723.640 861.050 2723.700 ;
        RECT 860.535 2723.500 861.050 2723.640 ;
        RECT 860.730 2723.440 861.050 2723.500 ;
        RECT 860.745 2720.920 861.035 2720.965 ;
        RECT 2901.750 2720.920 2902.070 2720.980 ;
        RECT 860.745 2720.780 2902.070 2720.920 ;
        RECT 860.745 2720.735 861.035 2720.780 ;
        RECT 2901.750 2720.720 2902.070 2720.780 ;
      LAYER via ;
        RECT 860.760 2723.440 861.020 2723.700 ;
        RECT 2901.780 2720.720 2902.040 2720.980 ;
      LAYER met2 ;
        RECT 859.390 2723.810 859.950 2731.680 ;
        RECT 859.390 2723.730 860.960 2723.810 ;
        RECT 859.390 2723.670 861.020 2723.730 ;
        RECT 859.390 2722.680 859.950 2723.670 ;
        RECT 860.760 2723.410 861.020 2723.670 ;
        RECT 2901.780 2720.690 2902.040 2721.010 ;
        RECT 2901.840 615.925 2901.980 2720.690 ;
        RECT 2901.770 615.555 2902.050 615.925 ;
      LAYER via2 ;
        RECT 2901.770 615.600 2902.050 615.880 ;
      LAYER met3 ;
        RECT 2901.745 615.890 2902.075 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2901.745 615.590 2924.800 615.890 ;
        RECT 2901.745 615.575 2902.075 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.350 2742.000 31.670 2742.060 ;
        RECT 1945.870 2742.000 1946.190 2742.060 ;
        RECT 31.350 2741.860 1946.190 2742.000 ;
        RECT 31.350 2741.800 31.670 2741.860 ;
        RECT 1945.870 2741.800 1946.190 2741.860 ;
        RECT 15.710 1620.680 16.030 1620.740 ;
        RECT 31.350 1620.680 31.670 1620.740 ;
        RECT 15.710 1620.540 31.670 1620.680 ;
        RECT 15.710 1620.480 16.030 1620.540 ;
        RECT 31.350 1620.480 31.670 1620.540 ;
      LAYER via ;
        RECT 31.380 2741.800 31.640 2742.060 ;
        RECT 1945.900 2741.800 1946.160 2742.060 ;
        RECT 15.740 1620.480 16.000 1620.740 ;
        RECT 31.380 1620.480 31.640 1620.740 ;
      LAYER met2 ;
        RECT 31.380 2741.770 31.640 2742.090 ;
        RECT 1945.900 2741.770 1946.160 2742.090 ;
        RECT 31.440 1620.770 31.580 2741.770 ;
        RECT 1945.960 2731.680 1946.100 2741.770 ;
        RECT 1945.910 2722.680 1946.470 2731.680 ;
        RECT 15.740 1620.450 16.000 1620.770 ;
        RECT 31.380 1620.450 31.640 1620.770 ;
        RECT 15.800 1615.525 15.940 1620.450 ;
        RECT 15.730 1615.155 16.010 1615.525 ;
      LAYER via2 ;
        RECT 15.730 1615.200 16.010 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 15.705 1615.490 16.035 1615.505 ;
        RECT -4.800 1615.190 16.035 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 15.705 1615.175 16.035 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 30.890 2740.980 31.210 2741.040 ;
        RECT 1984.510 2740.980 1984.830 2741.040 ;
        RECT 30.890 2740.840 1984.830 2740.980 ;
        RECT 30.890 2740.780 31.210 2740.840 ;
        RECT 1984.510 2740.780 1984.830 2740.840 ;
        RECT 15.710 1400.700 16.030 1400.760 ;
        RECT 30.890 1400.700 31.210 1400.760 ;
        RECT 15.710 1400.560 31.210 1400.700 ;
        RECT 15.710 1400.500 16.030 1400.560 ;
        RECT 30.890 1400.500 31.210 1400.560 ;
      LAYER via ;
        RECT 30.920 2740.780 31.180 2741.040 ;
        RECT 1984.540 2740.780 1984.800 2741.040 ;
        RECT 15.740 1400.500 16.000 1400.760 ;
        RECT 30.920 1400.500 31.180 1400.760 ;
      LAYER met2 ;
        RECT 30.920 2740.750 31.180 2741.070 ;
        RECT 1984.540 2740.750 1984.800 2741.070 ;
        RECT 30.980 1400.790 31.120 2740.750 ;
        RECT 1984.600 2731.680 1984.740 2740.750 ;
        RECT 1984.550 2722.680 1985.110 2731.680 ;
        RECT 15.740 1400.645 16.000 1400.790 ;
        RECT 15.730 1400.275 16.010 1400.645 ;
        RECT 30.920 1400.470 31.180 1400.790 ;
      LAYER via2 ;
        RECT 15.730 1400.320 16.010 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 15.705 1400.610 16.035 1400.625 ;
        RECT -4.800 1400.310 16.035 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 15.705 1400.295 16.035 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 51.590 2740.640 51.910 2740.700 ;
        RECT 2023.150 2740.640 2023.470 2740.700 ;
        RECT 51.590 2740.500 2023.470 2740.640 ;
        RECT 51.590 2740.440 51.910 2740.500 ;
        RECT 2023.150 2740.440 2023.470 2740.500 ;
        RECT 15.250 1186.840 15.570 1186.900 ;
        RECT 51.590 1186.840 51.910 1186.900 ;
        RECT 15.250 1186.700 51.910 1186.840 ;
        RECT 15.250 1186.640 15.570 1186.700 ;
        RECT 51.590 1186.640 51.910 1186.700 ;
      LAYER via ;
        RECT 51.620 2740.440 51.880 2740.700 ;
        RECT 2023.180 2740.440 2023.440 2740.700 ;
        RECT 15.280 1186.640 15.540 1186.900 ;
        RECT 51.620 1186.640 51.880 1186.900 ;
      LAYER met2 ;
        RECT 51.620 2740.410 51.880 2740.730 ;
        RECT 2023.180 2740.410 2023.440 2740.730 ;
        RECT 51.680 1186.930 51.820 2740.410 ;
        RECT 2023.240 2731.680 2023.380 2740.410 ;
        RECT 2023.190 2722.680 2023.750 2731.680 ;
        RECT 15.280 1186.610 15.540 1186.930 ;
        RECT 51.620 1186.610 51.880 1186.930 ;
        RECT 15.340 1185.085 15.480 1186.610 ;
        RECT 15.270 1184.715 15.550 1185.085 ;
      LAYER via2 ;
        RECT 15.270 1184.760 15.550 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 15.245 1185.050 15.575 1185.065 ;
        RECT -4.800 1184.750 15.575 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 15.245 1184.735 15.575 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2060.945 2721.105 2061.115 2723.315 ;
      LAYER mcon ;
        RECT 2060.945 2723.145 2061.115 2723.315 ;
      LAYER met1 ;
        RECT 2060.870 2723.300 2061.190 2723.360 ;
        RECT 2060.675 2723.160 2061.190 2723.300 ;
        RECT 2060.870 2723.100 2061.190 2723.160 ;
        RECT 24.910 2721.260 25.230 2721.320 ;
        RECT 2060.885 2721.260 2061.175 2721.305 ;
        RECT 24.910 2721.120 2061.175 2721.260 ;
        RECT 24.910 2721.060 25.230 2721.120 ;
        RECT 2060.885 2721.075 2061.175 2721.120 ;
        RECT 13.870 969.580 14.190 969.640 ;
        RECT 24.910 969.580 25.230 969.640 ;
        RECT 13.870 969.440 25.230 969.580 ;
        RECT 13.870 969.380 14.190 969.440 ;
        RECT 24.910 969.380 25.230 969.440 ;
      LAYER via ;
        RECT 2060.900 2723.100 2061.160 2723.360 ;
        RECT 24.940 2721.060 25.200 2721.320 ;
        RECT 13.900 969.380 14.160 969.640 ;
        RECT 24.940 969.380 25.200 969.640 ;
      LAYER met2 ;
        RECT 2060.900 2723.130 2061.160 2723.390 ;
        RECT 2062.290 2723.130 2062.850 2731.680 ;
        RECT 2060.900 2723.070 2062.850 2723.130 ;
        RECT 2060.960 2722.990 2062.850 2723.070 ;
        RECT 2062.290 2722.680 2062.850 2722.990 ;
        RECT 24.940 2721.030 25.200 2721.350 ;
        RECT 25.000 969.670 25.140 2721.030 ;
        RECT 13.900 969.525 14.160 969.670 ;
        RECT 13.890 969.155 14.170 969.525 ;
        RECT 24.940 969.350 25.200 969.670 ;
      LAYER via2 ;
        RECT 13.890 969.200 14.170 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 13.865 969.490 14.195 969.505 ;
        RECT -4.800 969.190 14.195 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 13.865 969.175 14.195 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 99.890 2739.960 100.210 2740.020 ;
        RECT 2100.890 2739.960 2101.210 2740.020 ;
        RECT 99.890 2739.820 2101.210 2739.960 ;
        RECT 99.890 2739.760 100.210 2739.820 ;
        RECT 2100.890 2739.760 2101.210 2739.820 ;
        RECT 16.630 758.780 16.950 758.840 ;
        RECT 99.890 758.780 100.210 758.840 ;
        RECT 16.630 758.640 100.210 758.780 ;
        RECT 16.630 758.580 16.950 758.640 ;
        RECT 99.890 758.580 100.210 758.640 ;
      LAYER via ;
        RECT 99.920 2739.760 100.180 2740.020 ;
        RECT 2100.920 2739.760 2101.180 2740.020 ;
        RECT 16.660 758.580 16.920 758.840 ;
        RECT 99.920 758.580 100.180 758.840 ;
      LAYER met2 ;
        RECT 99.920 2739.730 100.180 2740.050 ;
        RECT 2100.920 2739.730 2101.180 2740.050 ;
        RECT 99.980 758.870 100.120 2739.730 ;
        RECT 2100.980 2731.680 2101.120 2739.730 ;
        RECT 2100.930 2722.680 2101.490 2731.680 ;
        RECT 16.660 758.550 16.920 758.870 ;
        RECT 99.920 758.550 100.180 758.870 ;
        RECT 16.720 753.965 16.860 758.550 ;
        RECT 16.650 753.595 16.930 753.965 ;
      LAYER via2 ;
        RECT 16.650 753.640 16.930 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 16.625 753.930 16.955 753.945 ;
        RECT -4.800 753.630 16.955 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 16.625 753.615 16.955 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2139.145 2719.405 2139.315 2723.315 ;
      LAYER mcon ;
        RECT 2139.145 2723.145 2139.315 2723.315 ;
      LAYER met1 ;
        RECT 2139.070 2723.300 2139.390 2723.360 ;
        RECT 2139.070 2723.160 2139.585 2723.300 ;
        RECT 2139.070 2723.100 2139.390 2723.160 ;
        RECT 18.930 2719.560 19.250 2719.620 ;
        RECT 2139.085 2719.560 2139.375 2719.605 ;
        RECT 18.930 2719.420 2139.375 2719.560 ;
        RECT 18.930 2719.360 19.250 2719.420 ;
        RECT 2139.085 2719.375 2139.375 2719.420 ;
      LAYER via ;
        RECT 2139.100 2723.100 2139.360 2723.360 ;
        RECT 18.960 2719.360 19.220 2719.620 ;
      LAYER met2 ;
        RECT 2139.100 2723.130 2139.360 2723.390 ;
        RECT 2139.570 2723.130 2140.130 2731.680 ;
        RECT 2139.100 2723.070 2140.130 2723.130 ;
        RECT 2139.160 2722.990 2140.130 2723.070 ;
        RECT 2139.570 2722.680 2140.130 2722.990 ;
        RECT 18.960 2719.330 19.220 2719.650 ;
        RECT 19.020 538.405 19.160 2719.330 ;
        RECT 18.950 538.035 19.230 538.405 ;
      LAYER via2 ;
        RECT 18.950 538.080 19.230 538.360 ;
      LAYER met3 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 18.925 538.370 19.255 538.385 ;
        RECT -4.800 538.070 19.255 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 18.925 538.055 19.255 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 106.790 324.260 107.110 324.320 ;
        RECT 16.630 324.120 107.110 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 106.790 324.060 107.110 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 106.820 324.060 107.080 324.320 ;
      LAYER met2 ;
        RECT 106.810 2741.235 107.090 2741.605 ;
        RECT 2178.650 2741.235 2178.930 2741.605 ;
        RECT 106.880 324.350 107.020 2741.235 ;
        RECT 2178.720 2731.680 2178.860 2741.235 ;
        RECT 2178.670 2722.680 2179.230 2731.680 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 106.820 324.030 107.080 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 106.810 2741.280 107.090 2741.560 ;
        RECT 2178.650 2741.280 2178.930 2741.560 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 106.785 2741.570 107.115 2741.585 ;
        RECT 2178.625 2741.570 2178.955 2741.585 ;
        RECT 106.785 2741.270 2178.955 2741.570 ;
        RECT 106.785 2741.255 107.115 2741.270 ;
        RECT 2178.625 2741.255 2178.955 2741.270 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2215.505 2718.725 2215.675 2723.315 ;
      LAYER mcon ;
        RECT 2215.505 2723.145 2215.675 2723.315 ;
      LAYER met1 ;
        RECT 2215.430 2723.300 2215.750 2723.360 ;
        RECT 2215.235 2723.160 2215.750 2723.300 ;
        RECT 2215.430 2723.100 2215.750 2723.160 ;
        RECT 17.090 2718.880 17.410 2718.940 ;
        RECT 2215.445 2718.880 2215.735 2718.925 ;
        RECT 17.090 2718.740 2215.735 2718.880 ;
        RECT 17.090 2718.680 17.410 2718.740 ;
        RECT 2215.445 2718.695 2215.735 2718.740 ;
      LAYER via ;
        RECT 2215.460 2723.100 2215.720 2723.360 ;
        RECT 17.120 2718.680 17.380 2718.940 ;
      LAYER met2 ;
        RECT 2215.460 2723.130 2215.720 2723.390 ;
        RECT 2217.310 2723.130 2217.870 2731.680 ;
        RECT 2215.460 2723.070 2217.870 2723.130 ;
        RECT 2215.520 2722.990 2217.870 2723.070 ;
        RECT 2217.310 2722.680 2217.870 2722.990 ;
        RECT 17.120 2718.650 17.380 2718.970 ;
        RECT 17.180 107.285 17.320 2718.650 ;
        RECT 17.110 106.915 17.390 107.285 ;
      LAYER via2 ;
        RECT 17.110 106.960 17.390 107.240 ;
      LAYER met3 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 17.085 107.250 17.415 107.265 ;
        RECT -4.800 106.950 17.415 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 17.085 106.935 17.415 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 900.365 2721.785 900.535 2723.655 ;
      LAYER mcon ;
        RECT 900.365 2723.485 900.535 2723.655 ;
      LAYER met1 ;
        RECT 900.290 2723.640 900.610 2723.700 ;
        RECT 900.095 2723.500 900.610 2723.640 ;
        RECT 900.290 2723.440 900.610 2723.500 ;
        RECT 900.305 2721.940 900.595 2721.985 ;
        RECT 2902.210 2721.940 2902.530 2722.000 ;
        RECT 900.305 2721.800 2902.530 2721.940 ;
        RECT 900.305 2721.755 900.595 2721.800 ;
        RECT 2902.210 2721.740 2902.530 2721.800 ;
      LAYER via ;
        RECT 900.320 2723.440 900.580 2723.700 ;
        RECT 2902.240 2721.740 2902.500 2722.000 ;
      LAYER met2 ;
        RECT 898.490 2723.810 899.050 2731.680 ;
        RECT 898.490 2723.730 900.520 2723.810 ;
        RECT 898.490 2723.670 900.580 2723.730 ;
        RECT 898.490 2722.680 899.050 2723.670 ;
        RECT 900.320 2723.410 900.580 2723.670 ;
        RECT 2902.240 2721.710 2902.500 2722.030 ;
        RECT 2902.300 850.525 2902.440 2721.710 ;
        RECT 2902.230 850.155 2902.510 850.525 ;
      LAYER via2 ;
        RECT 2902.230 850.200 2902.510 850.480 ;
      LAYER met3 ;
        RECT 2902.205 850.490 2902.535 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2902.205 850.190 2924.800 850.490 ;
        RECT 2902.205 850.175 2902.535 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 938.010 2725.680 938.330 2725.740 ;
        RECT 2902.670 2725.680 2902.990 2725.740 ;
        RECT 938.010 2725.540 2902.990 2725.680 ;
        RECT 938.010 2725.480 938.330 2725.540 ;
        RECT 2902.670 2725.480 2902.990 2725.540 ;
      LAYER via ;
        RECT 938.040 2725.480 938.300 2725.740 ;
        RECT 2902.700 2725.480 2902.960 2725.740 ;
      LAYER met2 ;
        RECT 937.130 2725.850 937.690 2731.680 ;
        RECT 937.130 2725.770 938.240 2725.850 ;
        RECT 937.130 2725.710 938.300 2725.770 ;
        RECT 937.130 2722.680 937.690 2725.710 ;
        RECT 938.040 2725.450 938.300 2725.710 ;
        RECT 2902.700 2725.450 2902.960 2725.770 ;
        RECT 2902.760 1085.125 2902.900 2725.450 ;
        RECT 2902.690 1084.755 2902.970 1085.125 ;
      LAYER via2 ;
        RECT 2902.690 1084.800 2902.970 1085.080 ;
      LAYER met3 ;
        RECT 2902.665 1085.090 2902.995 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2902.665 1084.790 2924.800 1085.090 ;
        RECT 2902.665 1084.775 2902.995 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 977.645 2722.465 977.815 2723.655 ;
      LAYER mcon ;
        RECT 977.645 2723.485 977.815 2723.655 ;
      LAYER met1 ;
        RECT 977.570 2723.640 977.890 2723.700 ;
        RECT 977.375 2723.500 977.890 2723.640 ;
        RECT 977.570 2723.440 977.890 2723.500 ;
        RECT 977.585 2722.620 977.875 2722.665 ;
        RECT 2903.130 2722.620 2903.450 2722.680 ;
        RECT 977.585 2722.480 2903.450 2722.620 ;
        RECT 977.585 2722.435 977.875 2722.480 ;
        RECT 2903.130 2722.420 2903.450 2722.480 ;
      LAYER via ;
        RECT 977.600 2723.440 977.860 2723.700 ;
        RECT 2903.160 2722.420 2903.420 2722.680 ;
      LAYER met2 ;
        RECT 975.770 2723.810 976.330 2731.680 ;
        RECT 975.770 2723.730 977.800 2723.810 ;
        RECT 975.770 2723.670 977.860 2723.730 ;
        RECT 975.770 2722.680 976.330 2723.670 ;
        RECT 977.600 2723.410 977.860 2723.670 ;
        RECT 2903.160 2722.390 2903.420 2722.710 ;
        RECT 2903.220 1319.725 2903.360 2722.390 ;
        RECT 2903.150 1319.355 2903.430 1319.725 ;
      LAYER via2 ;
        RECT 2903.150 1319.400 2903.430 1319.680 ;
      LAYER met3 ;
        RECT 2903.125 1319.690 2903.455 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2903.125 1319.390 2924.800 1319.690 ;
        RECT 2903.125 1319.375 2903.455 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1014.870 2723.130 1015.430 2731.680 ;
        RECT 1015.770 2723.130 1016.050 2723.245 ;
        RECT 1014.870 2722.990 1016.050 2723.130 ;
        RECT 1014.870 2722.680 1015.430 2722.990 ;
        RECT 1015.770 2722.875 1016.050 2722.990 ;
        RECT 2904.070 2715.395 2904.350 2715.765 ;
        RECT 2904.140 1554.325 2904.280 2715.395 ;
        RECT 2904.070 1553.955 2904.350 1554.325 ;
      LAYER via2 ;
        RECT 1015.770 2722.920 1016.050 2723.200 ;
        RECT 2904.070 2715.440 2904.350 2715.720 ;
        RECT 2904.070 1554.000 2904.350 1554.280 ;
      LAYER met3 ;
        RECT 1015.745 2723.220 1016.075 2723.225 ;
        RECT 1015.745 2723.210 1016.330 2723.220 ;
        RECT 1015.745 2722.910 1016.530 2723.210 ;
        RECT 1015.745 2722.900 1016.330 2722.910 ;
        RECT 1015.745 2722.895 1016.075 2722.900 ;
        RECT 1015.950 2715.730 1016.330 2715.740 ;
        RECT 1155.790 2715.730 1156.170 2715.740 ;
        RECT 1015.950 2715.430 1156.170 2715.730 ;
        RECT 1015.950 2715.420 1016.330 2715.430 ;
        RECT 1155.790 2715.420 1156.170 2715.430 ;
        RECT 1159.470 2715.730 1159.850 2715.740 ;
        RECT 2904.045 2715.730 2904.375 2715.745 ;
        RECT 1159.470 2715.430 2904.375 2715.730 ;
        RECT 1159.470 2715.420 1159.850 2715.430 ;
        RECT 2904.045 2715.415 2904.375 2715.430 ;
        RECT 2904.045 1554.290 2904.375 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2904.045 1553.990 2924.800 1554.290 ;
        RECT 2904.045 1553.975 2904.375 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
      LAYER via3 ;
        RECT 1015.980 2722.900 1016.300 2723.220 ;
        RECT 1015.980 2715.420 1016.300 2715.740 ;
        RECT 1155.820 2715.420 1156.140 2715.740 ;
        RECT 1159.500 2715.420 1159.820 2715.740 ;
      LAYER met4 ;
        RECT 1015.975 2722.895 1016.305 2723.225 ;
        RECT 1015.990 2715.745 1016.290 2722.895 ;
        RECT 1015.975 2715.415 1016.305 2715.745 ;
        RECT 1155.815 2715.415 1156.145 2715.745 ;
        RECT 1159.495 2715.415 1159.825 2715.745 ;
        RECT 1155.830 2714.370 1156.130 2715.415 ;
        RECT 1159.510 2714.370 1159.810 2715.415 ;
        RECT 1155.830 2714.070 1159.810 2714.370 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1053.490 2745.315 1053.770 2745.685 ;
        RECT 1053.560 2731.680 1053.700 2745.315 ;
        RECT 1053.510 2722.680 1054.070 2731.680 ;
      LAYER via2 ;
        RECT 1053.490 2745.360 1053.770 2745.640 ;
      LAYER met3 ;
        RECT 1053.465 2745.650 1053.795 2745.665 ;
        RECT 2238.630 2745.650 2239.010 2745.660 ;
        RECT 1053.465 2745.350 2239.010 2745.650 ;
        RECT 1053.465 2745.335 1053.795 2745.350 ;
        RECT 2238.630 2745.340 2239.010 2745.350 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2916.710 1789.270 2924.800 1789.570 ;
        RECT 2238.630 1788.890 2239.010 1788.900 ;
        RECT 2238.630 1788.590 2256.450 1788.890 ;
        RECT 2238.630 1788.580 2239.010 1788.590 ;
        RECT 2256.150 1788.210 2256.450 1788.590 ;
        RECT 2304.910 1788.590 2353.050 1788.890 ;
        RECT 2256.150 1787.910 2304.290 1788.210 ;
        RECT 2303.990 1787.530 2304.290 1787.910 ;
        RECT 2304.910 1787.530 2305.210 1788.590 ;
        RECT 2352.750 1788.210 2353.050 1788.590 ;
        RECT 2401.510 1788.590 2449.650 1788.890 ;
        RECT 2352.750 1787.910 2400.890 1788.210 ;
        RECT 2303.990 1787.230 2305.210 1787.530 ;
        RECT 2400.590 1787.530 2400.890 1787.910 ;
        RECT 2401.510 1787.530 2401.810 1788.590 ;
        RECT 2449.350 1788.210 2449.650 1788.590 ;
        RECT 2498.110 1788.590 2546.250 1788.890 ;
        RECT 2449.350 1787.910 2497.490 1788.210 ;
        RECT 2400.590 1787.230 2401.810 1787.530 ;
        RECT 2497.190 1787.530 2497.490 1787.910 ;
        RECT 2498.110 1787.530 2498.410 1788.590 ;
        RECT 2545.950 1788.210 2546.250 1788.590 ;
        RECT 2594.710 1788.590 2642.850 1788.890 ;
        RECT 2545.950 1787.910 2594.090 1788.210 ;
        RECT 2497.190 1787.230 2498.410 1787.530 ;
        RECT 2593.790 1787.530 2594.090 1787.910 ;
        RECT 2594.710 1787.530 2595.010 1788.590 ;
        RECT 2642.550 1788.210 2642.850 1788.590 ;
        RECT 2691.310 1788.590 2739.450 1788.890 ;
        RECT 2642.550 1787.910 2690.690 1788.210 ;
        RECT 2593.790 1787.230 2595.010 1787.530 ;
        RECT 2690.390 1787.530 2690.690 1787.910 ;
        RECT 2691.310 1787.530 2691.610 1788.590 ;
        RECT 2739.150 1788.210 2739.450 1788.590 ;
        RECT 2787.910 1788.590 2836.050 1788.890 ;
        RECT 2739.150 1787.910 2787.290 1788.210 ;
        RECT 2690.390 1787.230 2691.610 1787.530 ;
        RECT 2786.990 1787.530 2787.290 1787.910 ;
        RECT 2787.910 1787.530 2788.210 1788.590 ;
        RECT 2835.750 1788.210 2836.050 1788.590 ;
        RECT 2916.710 1788.210 2917.010 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2835.750 1787.910 2883.890 1788.210 ;
        RECT 2786.990 1787.230 2788.210 1787.530 ;
        RECT 2883.590 1787.530 2883.890 1787.910 ;
        RECT 2884.510 1787.910 2917.010 1788.210 ;
        RECT 2884.510 1787.530 2884.810 1787.910 ;
        RECT 2883.590 1787.230 2884.810 1787.530 ;
      LAYER via3 ;
        RECT 2238.660 2745.340 2238.980 2745.660 ;
        RECT 2238.660 1788.580 2238.980 1788.900 ;
      LAYER met4 ;
        RECT 2238.655 2745.335 2238.985 2745.665 ;
        RECT 2238.670 1788.905 2238.970 2745.335 ;
        RECT 2238.655 1788.575 2238.985 1788.905 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1092.110 2745.400 1092.430 2745.460 ;
        RECT 2246.710 2745.400 2247.030 2745.460 ;
        RECT 1092.110 2745.260 2247.030 2745.400 ;
        RECT 1092.110 2745.200 1092.430 2745.260 ;
        RECT 2246.710 2745.200 2247.030 2745.260 ;
        RECT 2246.710 2028.340 2247.030 2028.400 ;
        RECT 2900.370 2028.340 2900.690 2028.400 ;
        RECT 2246.710 2028.200 2900.690 2028.340 ;
        RECT 2246.710 2028.140 2247.030 2028.200 ;
        RECT 2900.370 2028.140 2900.690 2028.200 ;
      LAYER via ;
        RECT 1092.140 2745.200 1092.400 2745.460 ;
        RECT 2246.740 2745.200 2247.000 2745.460 ;
        RECT 2246.740 2028.140 2247.000 2028.400 ;
        RECT 2900.400 2028.140 2900.660 2028.400 ;
      LAYER met2 ;
        RECT 1092.140 2745.170 1092.400 2745.490 ;
        RECT 2246.740 2745.170 2247.000 2745.490 ;
        RECT 1092.200 2731.680 1092.340 2745.170 ;
        RECT 1092.150 2722.680 1092.710 2731.680 ;
        RECT 2246.800 2028.430 2246.940 2745.170 ;
        RECT 2246.740 2028.110 2247.000 2028.430 ;
        RECT 2900.400 2028.110 2900.660 2028.430 ;
        RECT 2900.460 2024.205 2900.600 2028.110 ;
        RECT 2900.390 2023.835 2900.670 2024.205 ;
      LAYER via2 ;
        RECT 2900.390 2023.880 2900.670 2024.160 ;
      LAYER met3 ;
        RECT 2900.365 2024.170 2900.695 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.365 2023.870 2924.800 2024.170 ;
        RECT 2900.365 2023.855 2900.695 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1131.210 2746.080 1131.530 2746.140 ;
        RECT 2247.630 2746.080 2247.950 2746.140 ;
        RECT 1131.210 2745.940 2247.950 2746.080 ;
        RECT 1131.210 2745.880 1131.530 2745.940 ;
        RECT 2247.630 2745.880 2247.950 2745.940 ;
        RECT 2247.630 2262.940 2247.950 2263.000 ;
        RECT 2900.370 2262.940 2900.690 2263.000 ;
        RECT 2247.630 2262.800 2900.690 2262.940 ;
        RECT 2247.630 2262.740 2247.950 2262.800 ;
        RECT 2900.370 2262.740 2900.690 2262.800 ;
      LAYER via ;
        RECT 1131.240 2745.880 1131.500 2746.140 ;
        RECT 2247.660 2745.880 2247.920 2746.140 ;
        RECT 2247.660 2262.740 2247.920 2263.000 ;
        RECT 2900.400 2262.740 2900.660 2263.000 ;
      LAYER met2 ;
        RECT 1131.240 2745.850 1131.500 2746.170 ;
        RECT 2247.660 2745.850 2247.920 2746.170 ;
        RECT 1131.300 2731.680 1131.440 2745.850 ;
        RECT 1131.250 2722.680 1131.810 2731.680 ;
        RECT 2247.720 2263.030 2247.860 2745.850 ;
        RECT 2247.660 2262.710 2247.920 2263.030 ;
        RECT 2900.400 2262.710 2900.660 2263.030 ;
        RECT 2900.460 2258.805 2900.600 2262.710 ;
        RECT 2900.390 2258.435 2900.670 2258.805 ;
      LAYER via2 ;
        RECT 2900.390 2258.480 2900.670 2258.760 ;
      LAYER met3 ;
        RECT 2900.365 2258.770 2900.695 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.365 2258.470 2924.800 2258.770 ;
        RECT 2900.365 2258.455 2900.695 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1070.105 1014.305 1070.275 1049.155 ;
        RECT 1070.565 161.925 1070.735 234.515 ;
      LAYER mcon ;
        RECT 1070.105 1048.985 1070.275 1049.155 ;
        RECT 1070.565 234.345 1070.735 234.515 ;
      LAYER met1 ;
        RECT 1070.030 1049.140 1070.350 1049.200 ;
        RECT 1069.835 1049.000 1070.350 1049.140 ;
        RECT 1070.030 1048.940 1070.350 1049.000 ;
        RECT 1070.030 1014.460 1070.350 1014.520 ;
        RECT 1069.835 1014.320 1070.350 1014.460 ;
        RECT 1070.030 1014.260 1070.350 1014.320 ;
        RECT 1070.030 966.180 1070.350 966.240 ;
        RECT 1070.490 966.180 1070.810 966.240 ;
        RECT 1070.030 966.040 1070.810 966.180 ;
        RECT 1070.030 965.980 1070.350 966.040 ;
        RECT 1070.490 965.980 1070.810 966.040 ;
        RECT 1070.490 497.120 1070.810 497.380 ;
        RECT 1070.580 496.700 1070.720 497.120 ;
        RECT 1070.490 496.440 1070.810 496.700 ;
        RECT 1070.490 289.920 1070.810 289.980 ;
        RECT 1070.950 289.920 1071.270 289.980 ;
        RECT 1070.490 289.780 1071.270 289.920 ;
        RECT 1070.490 289.720 1070.810 289.780 ;
        RECT 1070.950 289.720 1071.270 289.780 ;
        RECT 1070.030 234.500 1070.350 234.560 ;
        RECT 1070.505 234.500 1070.795 234.545 ;
        RECT 1070.030 234.360 1070.795 234.500 ;
        RECT 1070.030 234.300 1070.350 234.360 ;
        RECT 1070.505 234.315 1070.795 234.360 ;
        RECT 1069.570 162.080 1069.890 162.140 ;
        RECT 1070.505 162.080 1070.795 162.125 ;
        RECT 1069.570 161.940 1070.795 162.080 ;
        RECT 1069.570 161.880 1069.890 161.940 ;
        RECT 1070.505 161.895 1070.795 161.940 ;
        RECT 633.030 36.960 633.350 37.020 ;
        RECT 1070.490 36.960 1070.810 37.020 ;
        RECT 633.030 36.820 1070.810 36.960 ;
        RECT 633.030 36.760 633.350 36.820 ;
        RECT 1070.490 36.760 1070.810 36.820 ;
      LAYER via ;
        RECT 1070.060 1048.940 1070.320 1049.200 ;
        RECT 1070.060 1014.260 1070.320 1014.520 ;
        RECT 1070.060 965.980 1070.320 966.240 ;
        RECT 1070.520 965.980 1070.780 966.240 ;
        RECT 1070.520 497.120 1070.780 497.380 ;
        RECT 1070.520 496.440 1070.780 496.700 ;
        RECT 1070.520 289.720 1070.780 289.980 ;
        RECT 1070.980 289.720 1071.240 289.980 ;
        RECT 1070.060 234.300 1070.320 234.560 ;
        RECT 1069.600 161.880 1069.860 162.140 ;
        RECT 633.060 36.760 633.320 37.020 ;
        RECT 1070.520 36.760 1070.780 37.020 ;
      LAYER met2 ;
        RECT 1075.130 1220.330 1075.690 1228.680 ;
        RECT 1073.340 1220.190 1075.690 1220.330 ;
        RECT 1073.340 1196.530 1073.480 1220.190 ;
        RECT 1075.130 1219.680 1075.690 1220.190 ;
        RECT 1070.580 1196.390 1073.480 1196.530 ;
        RECT 1070.580 1097.250 1070.720 1196.390 ;
        RECT 1070.120 1097.110 1070.720 1097.250 ;
        RECT 1070.120 1049.230 1070.260 1097.110 ;
        RECT 1070.060 1048.910 1070.320 1049.230 ;
        RECT 1070.060 1014.230 1070.320 1014.550 ;
        RECT 1070.120 966.270 1070.260 1014.230 ;
        RECT 1070.060 965.950 1070.320 966.270 ;
        RECT 1070.520 965.950 1070.780 966.270 ;
        RECT 1070.580 883.050 1070.720 965.950 ;
        RECT 1070.120 882.910 1070.720 883.050 ;
        RECT 1070.120 881.690 1070.260 882.910 ;
        RECT 1070.120 881.550 1070.720 881.690 ;
        RECT 1070.580 787.170 1070.720 881.550 ;
        RECT 1070.120 787.030 1070.720 787.170 ;
        RECT 1070.120 786.490 1070.260 787.030 ;
        RECT 1070.120 786.350 1070.720 786.490 ;
        RECT 1070.580 497.410 1070.720 786.350 ;
        RECT 1070.520 497.090 1070.780 497.410 ;
        RECT 1070.520 496.410 1070.780 496.730 ;
        RECT 1070.580 403.650 1070.720 496.410 ;
        RECT 1070.580 403.510 1071.180 403.650 ;
        RECT 1071.040 290.010 1071.180 403.510 ;
        RECT 1070.520 289.690 1070.780 290.010 ;
        RECT 1070.980 289.690 1071.240 290.010 ;
        RECT 1070.580 241.810 1070.720 289.690 ;
        RECT 1070.120 241.670 1070.720 241.810 ;
        RECT 1070.120 234.590 1070.260 241.670 ;
        RECT 1070.060 234.270 1070.320 234.590 ;
        RECT 1069.600 161.850 1069.860 162.170 ;
        RECT 1069.660 96.970 1069.800 161.850 ;
        RECT 1069.660 96.830 1070.260 96.970 ;
        RECT 1070.120 75.890 1070.260 96.830 ;
        RECT 1070.120 75.750 1070.720 75.890 ;
        RECT 1070.580 37.050 1070.720 75.750 ;
        RECT 633.060 36.730 633.320 37.050 ;
        RECT 1070.520 36.730 1070.780 37.050 ;
        RECT 633.120 2.400 633.260 36.730 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 34.240 1994.030 34.300 ;
        RECT 2417.370 34.240 2417.690 34.300 ;
        RECT 1993.710 34.100 2417.690 34.240 ;
        RECT 1993.710 34.040 1994.030 34.100 ;
        RECT 2417.370 34.040 2417.690 34.100 ;
      LAYER via ;
        RECT 1993.740 34.040 1994.000 34.300 ;
        RECT 2417.400 34.040 2417.660 34.300 ;
      LAYER met2 ;
        RECT 1991.450 1220.330 1992.010 1228.680 ;
        RECT 1991.450 1220.190 1993.940 1220.330 ;
        RECT 1991.450 1219.680 1992.010 1220.190 ;
        RECT 1993.800 34.330 1993.940 1220.190 ;
        RECT 1993.740 34.010 1994.000 34.330 ;
        RECT 2417.400 34.010 2417.660 34.330 ;
        RECT 2417.460 2.400 2417.600 34.010 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.150 35.260 2000.470 35.320 ;
        RECT 2434.850 35.260 2435.170 35.320 ;
        RECT 2000.150 35.120 2435.170 35.260 ;
        RECT 2000.150 35.060 2000.470 35.120 ;
        RECT 2434.850 35.060 2435.170 35.120 ;
      LAYER via ;
        RECT 2000.180 35.060 2000.440 35.320 ;
        RECT 2434.880 35.060 2435.140 35.320 ;
      LAYER met2 ;
        RECT 2000.650 1220.330 2001.210 1228.680 ;
        RECT 2000.240 1220.190 2001.210 1220.330 ;
        RECT 2000.240 35.350 2000.380 1220.190 ;
        RECT 2000.650 1219.680 2001.210 1220.190 ;
        RECT 2000.180 35.030 2000.440 35.350 ;
        RECT 2434.880 35.030 2435.140 35.350 ;
        RECT 2434.940 2.400 2435.080 35.030 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2009.810 1207.580 2010.130 1207.640 ;
        RECT 2013.950 1207.580 2014.270 1207.640 ;
        RECT 2009.810 1207.440 2014.270 1207.580 ;
        RECT 2009.810 1207.380 2010.130 1207.440 ;
        RECT 2013.950 1207.380 2014.270 1207.440 ;
        RECT 2013.950 35.600 2014.270 35.660 ;
        RECT 2452.790 35.600 2453.110 35.660 ;
        RECT 2013.950 35.460 2453.110 35.600 ;
        RECT 2013.950 35.400 2014.270 35.460 ;
        RECT 2452.790 35.400 2453.110 35.460 ;
      LAYER via ;
        RECT 2009.840 1207.380 2010.100 1207.640 ;
        RECT 2013.980 1207.380 2014.240 1207.640 ;
        RECT 2013.980 35.400 2014.240 35.660 ;
        RECT 2452.820 35.400 2453.080 35.660 ;
      LAYER met2 ;
        RECT 2009.850 1219.680 2010.410 1228.680 ;
        RECT 2009.900 1207.670 2010.040 1219.680 ;
        RECT 2009.840 1207.350 2010.100 1207.670 ;
        RECT 2013.980 1207.350 2014.240 1207.670 ;
        RECT 2014.040 35.690 2014.180 1207.350 ;
        RECT 2013.980 35.370 2014.240 35.690 ;
        RECT 2452.820 35.370 2453.080 35.690 ;
        RECT 2452.880 2.400 2453.020 35.370 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 35.940 2021.630 36.000 ;
        RECT 2470.730 35.940 2471.050 36.000 ;
        RECT 2021.310 35.800 2471.050 35.940 ;
        RECT 2021.310 35.740 2021.630 35.800 ;
        RECT 2470.730 35.740 2471.050 35.800 ;
      LAYER via ;
        RECT 2021.340 35.740 2021.600 36.000 ;
        RECT 2470.760 35.740 2471.020 36.000 ;
      LAYER met2 ;
        RECT 2019.050 1220.330 2019.610 1228.680 ;
        RECT 2019.050 1220.190 2021.540 1220.330 ;
        RECT 2019.050 1219.680 2019.610 1220.190 ;
        RECT 2021.400 36.030 2021.540 1220.190 ;
        RECT 2021.340 35.710 2021.600 36.030 ;
        RECT 2470.760 35.710 2471.020 36.030 ;
        RECT 2470.820 2.400 2470.960 35.710 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2027.750 36.280 2028.070 36.340 ;
        RECT 2488.670 36.280 2488.990 36.340 ;
        RECT 2027.750 36.140 2488.990 36.280 ;
        RECT 2027.750 36.080 2028.070 36.140 ;
        RECT 2488.670 36.080 2488.990 36.140 ;
      LAYER via ;
        RECT 2027.780 36.080 2028.040 36.340 ;
        RECT 2488.700 36.080 2488.960 36.340 ;
      LAYER met2 ;
        RECT 2028.250 1220.330 2028.810 1228.680 ;
        RECT 2027.840 1220.190 2028.810 1220.330 ;
        RECT 2027.840 36.370 2027.980 1220.190 ;
        RECT 2028.250 1219.680 2028.810 1220.190 ;
        RECT 2027.780 36.050 2028.040 36.370 ;
        RECT 2488.700 36.050 2488.960 36.370 ;
        RECT 2488.760 2.400 2488.900 36.050 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2037.410 1207.580 2037.730 1207.640 ;
        RECT 2041.550 1207.580 2041.870 1207.640 ;
        RECT 2037.410 1207.440 2041.870 1207.580 ;
        RECT 2037.410 1207.380 2037.730 1207.440 ;
        RECT 2041.550 1207.380 2041.870 1207.440 ;
        RECT 2041.550 36.620 2041.870 36.680 ;
        RECT 2506.150 36.620 2506.470 36.680 ;
        RECT 2041.550 36.480 2506.470 36.620 ;
        RECT 2041.550 36.420 2041.870 36.480 ;
        RECT 2506.150 36.420 2506.470 36.480 ;
      LAYER via ;
        RECT 2037.440 1207.380 2037.700 1207.640 ;
        RECT 2041.580 1207.380 2041.840 1207.640 ;
        RECT 2041.580 36.420 2041.840 36.680 ;
        RECT 2506.180 36.420 2506.440 36.680 ;
      LAYER met2 ;
        RECT 2037.450 1219.680 2038.010 1228.680 ;
        RECT 2037.500 1207.670 2037.640 1219.680 ;
        RECT 2037.440 1207.350 2037.700 1207.670 ;
        RECT 2041.580 1207.350 2041.840 1207.670 ;
        RECT 2041.640 36.710 2041.780 1207.350 ;
        RECT 2041.580 36.390 2041.840 36.710 ;
        RECT 2506.180 36.390 2506.440 36.710 ;
        RECT 2506.240 2.400 2506.380 36.390 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 36.960 2049.230 37.020 ;
        RECT 2524.090 36.960 2524.410 37.020 ;
        RECT 2048.910 36.820 2524.410 36.960 ;
        RECT 2048.910 36.760 2049.230 36.820 ;
        RECT 2524.090 36.760 2524.410 36.820 ;
      LAYER via ;
        RECT 2048.940 36.760 2049.200 37.020 ;
        RECT 2524.120 36.760 2524.380 37.020 ;
      LAYER met2 ;
        RECT 2046.650 1220.330 2047.210 1228.680 ;
        RECT 2046.650 1220.190 2049.140 1220.330 ;
        RECT 2046.650 1219.680 2047.210 1220.190 ;
        RECT 2049.000 37.050 2049.140 1220.190 ;
        RECT 2048.940 36.730 2049.200 37.050 ;
        RECT 2524.120 36.730 2524.380 37.050 ;
        RECT 2524.180 2.400 2524.320 36.730 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.350 37.300 2055.670 37.360 ;
        RECT 2542.030 37.300 2542.350 37.360 ;
        RECT 2055.350 37.160 2542.350 37.300 ;
        RECT 2055.350 37.100 2055.670 37.160 ;
        RECT 2542.030 37.100 2542.350 37.160 ;
      LAYER via ;
        RECT 2055.380 37.100 2055.640 37.360 ;
        RECT 2542.060 37.100 2542.320 37.360 ;
      LAYER met2 ;
        RECT 2055.390 1219.680 2055.950 1228.680 ;
        RECT 2055.440 37.390 2055.580 1219.680 ;
        RECT 2055.380 37.070 2055.640 37.390 ;
        RECT 2542.060 37.070 2542.320 37.390 ;
        RECT 2542.120 2.400 2542.260 37.070 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2064.550 1210.640 2064.870 1210.700 ;
        RECT 2069.610 1210.640 2069.930 1210.700 ;
        RECT 2064.550 1210.500 2069.930 1210.640 ;
        RECT 2064.550 1210.440 2064.870 1210.500 ;
        RECT 2069.610 1210.440 2069.930 1210.500 ;
        RECT 2069.610 21.320 2069.930 21.380 ;
        RECT 2559.970 21.320 2560.290 21.380 ;
        RECT 2069.610 21.180 2560.290 21.320 ;
        RECT 2069.610 21.120 2069.930 21.180 ;
        RECT 2559.970 21.120 2560.290 21.180 ;
      LAYER via ;
        RECT 2064.580 1210.440 2064.840 1210.700 ;
        RECT 2069.640 1210.440 2069.900 1210.700 ;
        RECT 2069.640 21.120 2069.900 21.380 ;
        RECT 2560.000 21.120 2560.260 21.380 ;
      LAYER met2 ;
        RECT 2064.590 1219.680 2065.150 1228.680 ;
        RECT 2064.640 1210.730 2064.780 1219.680 ;
        RECT 2064.580 1210.410 2064.840 1210.730 ;
        RECT 2069.640 1210.410 2069.900 1210.730 ;
        RECT 2069.700 21.410 2069.840 1210.410 ;
        RECT 2069.640 21.090 2069.900 21.410 ;
        RECT 2560.000 21.090 2560.260 21.410 ;
        RECT 2560.060 2.400 2560.200 21.090 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.510 21.660 2076.830 21.720 ;
        RECT 2577.910 21.660 2578.230 21.720 ;
        RECT 2076.510 21.520 2578.230 21.660 ;
        RECT 2076.510 21.460 2076.830 21.520 ;
        RECT 2577.910 21.460 2578.230 21.520 ;
      LAYER via ;
        RECT 2076.540 21.460 2076.800 21.720 ;
        RECT 2577.940 21.460 2578.200 21.720 ;
      LAYER met2 ;
        RECT 2073.790 1220.330 2074.350 1228.680 ;
        RECT 2073.790 1220.190 2076.740 1220.330 ;
        RECT 2073.790 1219.680 2074.350 1220.190 ;
        RECT 2076.600 21.750 2076.740 1220.190 ;
        RECT 2076.540 21.430 2076.800 21.750 ;
        RECT 2577.940 21.430 2578.200 21.750 ;
        RECT 2578.000 2.400 2578.140 21.430 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 811.510 37.980 811.830 38.040 ;
        RECT 1167.090 37.980 1167.410 38.040 ;
        RECT 811.510 37.840 1167.410 37.980 ;
        RECT 811.510 37.780 811.830 37.840 ;
        RECT 1167.090 37.780 1167.410 37.840 ;
      LAYER via ;
        RECT 811.540 37.780 811.800 38.040 ;
        RECT 1167.120 37.780 1167.380 38.040 ;
      LAYER met2 ;
        RECT 1166.670 1220.330 1167.230 1228.680 ;
        RECT 1166.670 1219.680 1167.320 1220.330 ;
        RECT 1167.180 38.070 1167.320 1219.680 ;
        RECT 811.540 37.750 811.800 38.070 ;
        RECT 1167.120 37.750 1167.380 38.070 ;
        RECT 811.600 2.400 811.740 37.750 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2120.285 22.185 2120.455 27.115 ;
      LAYER mcon ;
        RECT 2120.285 26.945 2120.455 27.115 ;
      LAYER met1 ;
        RECT 2082.950 27.440 2083.270 27.500 ;
        RECT 2082.950 27.300 2096.980 27.440 ;
        RECT 2082.950 27.240 2083.270 27.300 ;
        RECT 2096.840 27.100 2096.980 27.300 ;
        RECT 2120.225 27.100 2120.515 27.145 ;
        RECT 2096.840 26.960 2120.515 27.100 ;
        RECT 2120.225 26.915 2120.515 26.960 ;
        RECT 2120.225 22.340 2120.515 22.385 ;
        RECT 2595.390 22.340 2595.710 22.400 ;
        RECT 2120.225 22.200 2595.710 22.340 ;
        RECT 2120.225 22.155 2120.515 22.200 ;
        RECT 2595.390 22.140 2595.710 22.200 ;
      LAYER via ;
        RECT 2082.980 27.240 2083.240 27.500 ;
        RECT 2595.420 22.140 2595.680 22.400 ;
      LAYER met2 ;
        RECT 2082.990 1219.680 2083.550 1228.680 ;
        RECT 2083.040 27.530 2083.180 1219.680 ;
        RECT 2082.980 27.210 2083.240 27.530 ;
        RECT 2595.420 22.110 2595.680 22.430 ;
        RECT 2595.480 2.400 2595.620 22.110 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2114.305 27.625 2115.395 27.795 ;
        RECT 2114.305 27.285 2114.475 27.625 ;
        RECT 2115.225 25.415 2115.395 27.625 ;
        RECT 2115.225 25.245 2116.775 25.415 ;
        RECT 2116.605 23.885 2116.775 25.245 ;
      LAYER met1 ;
        RECT 2092.150 1207.580 2092.470 1207.640 ;
        RECT 2097.210 1207.580 2097.530 1207.640 ;
        RECT 2092.150 1207.440 2097.530 1207.580 ;
        RECT 2092.150 1207.380 2092.470 1207.440 ;
        RECT 2097.210 1207.380 2097.530 1207.440 ;
        RECT 2097.210 27.440 2097.530 27.500 ;
        RECT 2114.245 27.440 2114.535 27.485 ;
        RECT 2097.210 27.300 2114.535 27.440 ;
        RECT 2097.210 27.240 2097.530 27.300 ;
        RECT 2114.245 27.255 2114.535 27.300 ;
        RECT 2116.545 24.040 2116.835 24.085 ;
        RECT 2138.150 24.040 2138.470 24.100 ;
        RECT 2116.545 23.900 2138.470 24.040 ;
        RECT 2116.545 23.855 2116.835 23.900 ;
        RECT 2138.150 23.840 2138.470 23.900 ;
        RECT 2139.530 22.000 2139.850 22.060 ;
        RECT 2613.330 22.000 2613.650 22.060 ;
        RECT 2139.530 21.860 2613.650 22.000 ;
        RECT 2139.530 21.800 2139.850 21.860 ;
        RECT 2613.330 21.800 2613.650 21.860 ;
      LAYER via ;
        RECT 2092.180 1207.380 2092.440 1207.640 ;
        RECT 2097.240 1207.380 2097.500 1207.640 ;
        RECT 2097.240 27.240 2097.500 27.500 ;
        RECT 2138.180 23.840 2138.440 24.100 ;
        RECT 2139.560 21.800 2139.820 22.060 ;
        RECT 2613.360 21.800 2613.620 22.060 ;
      LAYER met2 ;
        RECT 2092.190 1219.680 2092.750 1228.680 ;
        RECT 2092.240 1207.670 2092.380 1219.680 ;
        RECT 2092.180 1207.350 2092.440 1207.670 ;
        RECT 2097.240 1207.350 2097.500 1207.670 ;
        RECT 2097.300 27.530 2097.440 1207.350 ;
        RECT 2097.240 27.210 2097.500 27.530 ;
        RECT 2138.180 23.810 2138.440 24.130 ;
        RECT 2138.240 22.285 2138.380 23.810 ;
        RECT 2138.170 21.915 2138.450 22.285 ;
        RECT 2139.550 21.915 2139.830 22.285 ;
        RECT 2139.560 21.770 2139.820 21.915 ;
        RECT 2613.360 21.770 2613.620 22.090 ;
        RECT 2613.420 2.400 2613.560 21.770 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
      LAYER via2 ;
        RECT 2138.170 21.960 2138.450 22.240 ;
        RECT 2139.550 21.960 2139.830 22.240 ;
      LAYER met3 ;
        RECT 2138.145 22.250 2138.475 22.265 ;
        RECT 2139.525 22.250 2139.855 22.265 ;
        RECT 2138.145 21.950 2139.855 22.250 ;
        RECT 2138.145 21.935 2138.475 21.950 ;
        RECT 2139.525 21.935 2139.855 21.950 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2116.605 25.585 2116.775 40.715 ;
        RECT 2132.245 22.525 2132.415 25.755 ;
      LAYER mcon ;
        RECT 2116.605 40.545 2116.775 40.715 ;
        RECT 2132.245 25.585 2132.415 25.755 ;
      LAYER met1 ;
        RECT 2104.110 40.700 2104.430 40.760 ;
        RECT 2116.545 40.700 2116.835 40.745 ;
        RECT 2104.110 40.560 2116.835 40.700 ;
        RECT 2104.110 40.500 2104.430 40.560 ;
        RECT 2116.545 40.515 2116.835 40.560 ;
        RECT 2116.545 25.740 2116.835 25.785 ;
        RECT 2132.185 25.740 2132.475 25.785 ;
        RECT 2116.545 25.600 2132.475 25.740 ;
        RECT 2116.545 25.555 2116.835 25.600 ;
        RECT 2132.185 25.555 2132.475 25.600 ;
        RECT 2132.185 22.680 2132.475 22.725 ;
        RECT 2631.270 22.680 2631.590 22.740 ;
        RECT 2132.185 22.540 2631.590 22.680 ;
        RECT 2132.185 22.495 2132.475 22.540 ;
        RECT 2631.270 22.480 2631.590 22.540 ;
      LAYER via ;
        RECT 2104.140 40.500 2104.400 40.760 ;
        RECT 2631.300 22.480 2631.560 22.740 ;
      LAYER met2 ;
        RECT 2101.390 1220.330 2101.950 1228.680 ;
        RECT 2101.390 1220.190 2104.340 1220.330 ;
        RECT 2101.390 1219.680 2101.950 1220.190 ;
        RECT 2104.200 40.790 2104.340 1220.190 ;
        RECT 2104.140 40.470 2104.400 40.790 ;
        RECT 2631.300 22.450 2631.560 22.770 ;
        RECT 2631.360 2.400 2631.500 22.450 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2114.305 23.035 2114.475 23.715 ;
        RECT 2114.305 22.865 2115.395 23.035 ;
      LAYER mcon ;
        RECT 2114.305 23.545 2114.475 23.715 ;
        RECT 2115.225 22.865 2115.395 23.035 ;
      LAYER met1 ;
        RECT 2111.010 23.700 2111.330 23.760 ;
        RECT 2114.245 23.700 2114.535 23.745 ;
        RECT 2111.010 23.560 2114.535 23.700 ;
        RECT 2111.010 23.500 2111.330 23.560 ;
        RECT 2114.245 23.515 2114.535 23.560 ;
        RECT 2115.165 23.020 2115.455 23.065 ;
        RECT 2649.210 23.020 2649.530 23.080 ;
        RECT 2115.165 22.880 2649.530 23.020 ;
        RECT 2115.165 22.835 2115.455 22.880 ;
        RECT 2649.210 22.820 2649.530 22.880 ;
      LAYER via ;
        RECT 2111.040 23.500 2111.300 23.760 ;
        RECT 2649.240 22.820 2649.500 23.080 ;
      LAYER met2 ;
        RECT 2110.590 1220.330 2111.150 1228.680 ;
        RECT 2110.590 1219.680 2111.240 1220.330 ;
        RECT 2111.100 23.790 2111.240 1219.680 ;
        RECT 2111.040 23.470 2111.300 23.790 ;
        RECT 2649.240 22.790 2649.500 23.110 ;
        RECT 2649.300 2.400 2649.440 22.790 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2123.505 1062.585 2123.675 1110.695 ;
        RECT 2122.585 869.125 2122.755 910.775 ;
        RECT 2123.505 786.505 2123.675 814.215 ;
        RECT 2123.505 689.605 2123.675 717.655 ;
        RECT 2123.505 621.265 2123.675 669.375 ;
        RECT 2123.505 572.645 2123.675 620.755 ;
        RECT 2123.505 496.485 2123.675 535.415 ;
        RECT 2123.505 386.325 2123.675 434.775 ;
        RECT 2123.505 289.765 2123.675 337.875 ;
        RECT 2123.505 193.205 2123.675 241.315 ;
      LAYER mcon ;
        RECT 2123.505 1110.525 2123.675 1110.695 ;
        RECT 2122.585 910.605 2122.755 910.775 ;
        RECT 2123.505 814.045 2123.675 814.215 ;
        RECT 2123.505 717.485 2123.675 717.655 ;
        RECT 2123.505 669.205 2123.675 669.375 ;
        RECT 2123.505 620.585 2123.675 620.755 ;
        RECT 2123.505 535.245 2123.675 535.415 ;
        RECT 2123.505 434.605 2123.675 434.775 ;
        RECT 2123.505 337.705 2123.675 337.875 ;
        RECT 2123.505 241.145 2123.675 241.315 ;
      LAYER met1 ;
        RECT 2119.750 1207.580 2120.070 1207.640 ;
        RECT 2123.890 1207.580 2124.210 1207.640 ;
        RECT 2119.750 1207.440 2124.210 1207.580 ;
        RECT 2119.750 1207.380 2120.070 1207.440 ;
        RECT 2123.890 1207.380 2124.210 1207.440 ;
        RECT 2123.430 1111.360 2123.750 1111.420 ;
        RECT 2123.890 1111.360 2124.210 1111.420 ;
        RECT 2123.430 1111.220 2124.210 1111.360 ;
        RECT 2123.430 1111.160 2123.750 1111.220 ;
        RECT 2123.890 1111.160 2124.210 1111.220 ;
        RECT 2123.430 1110.680 2123.750 1110.740 ;
        RECT 2123.235 1110.540 2123.750 1110.680 ;
        RECT 2123.430 1110.480 2123.750 1110.540 ;
        RECT 2123.445 1062.740 2123.735 1062.785 ;
        RECT 2123.890 1062.740 2124.210 1062.800 ;
        RECT 2123.445 1062.600 2124.210 1062.740 ;
        RECT 2123.445 1062.555 2123.735 1062.600 ;
        RECT 2123.890 1062.540 2124.210 1062.600 ;
        RECT 2122.970 1014.460 2123.290 1014.520 ;
        RECT 2123.430 1014.460 2123.750 1014.520 ;
        RECT 2122.970 1014.320 2123.750 1014.460 ;
        RECT 2122.970 1014.260 2123.290 1014.320 ;
        RECT 2123.430 1014.260 2123.750 1014.320 ;
        RECT 2122.510 966.180 2122.830 966.240 ;
        RECT 2123.890 966.180 2124.210 966.240 ;
        RECT 2122.510 966.040 2124.210 966.180 ;
        RECT 2122.510 965.980 2122.830 966.040 ;
        RECT 2123.890 965.980 2124.210 966.040 ;
        RECT 2122.970 917.900 2123.290 917.960 ;
        RECT 2123.430 917.900 2123.750 917.960 ;
        RECT 2122.970 917.760 2123.750 917.900 ;
        RECT 2122.970 917.700 2123.290 917.760 ;
        RECT 2123.430 917.700 2123.750 917.760 ;
        RECT 2122.510 910.760 2122.830 910.820 ;
        RECT 2122.315 910.620 2122.830 910.760 ;
        RECT 2122.510 910.560 2122.830 910.620 ;
        RECT 2122.525 869.280 2122.815 869.325 ;
        RECT 2123.430 869.280 2123.750 869.340 ;
        RECT 2122.525 869.140 2123.750 869.280 ;
        RECT 2122.525 869.095 2122.815 869.140 ;
        RECT 2123.430 869.080 2123.750 869.140 ;
        RECT 2123.430 862.480 2123.750 862.540 ;
        RECT 2124.810 862.480 2125.130 862.540 ;
        RECT 2123.430 862.340 2125.130 862.480 ;
        RECT 2123.430 862.280 2123.750 862.340 ;
        RECT 2124.810 862.280 2125.130 862.340 ;
        RECT 2123.430 814.200 2123.750 814.260 ;
        RECT 2123.235 814.060 2123.750 814.200 ;
        RECT 2123.430 814.000 2123.750 814.060 ;
        RECT 2123.430 786.660 2123.750 786.720 ;
        RECT 2123.235 786.520 2123.750 786.660 ;
        RECT 2123.430 786.460 2123.750 786.520 ;
        RECT 2123.430 765.920 2123.750 765.980 ;
        RECT 2123.890 765.920 2124.210 765.980 ;
        RECT 2123.430 765.780 2124.210 765.920 ;
        RECT 2123.430 765.720 2123.750 765.780 ;
        RECT 2123.890 765.720 2124.210 765.780 ;
        RECT 2123.430 717.640 2123.750 717.700 ;
        RECT 2123.235 717.500 2123.750 717.640 ;
        RECT 2123.430 717.440 2123.750 717.500 ;
        RECT 2123.430 689.760 2123.750 689.820 ;
        RECT 2123.235 689.620 2123.750 689.760 ;
        RECT 2123.430 689.560 2123.750 689.620 ;
        RECT 2123.445 669.360 2123.735 669.405 ;
        RECT 2123.890 669.360 2124.210 669.420 ;
        RECT 2123.445 669.220 2124.210 669.360 ;
        RECT 2123.445 669.175 2123.735 669.220 ;
        RECT 2123.890 669.160 2124.210 669.220 ;
        RECT 2123.430 621.420 2123.750 621.480 ;
        RECT 2123.235 621.280 2123.750 621.420 ;
        RECT 2123.430 621.220 2123.750 621.280 ;
        RECT 2123.430 620.740 2123.750 620.800 ;
        RECT 2123.235 620.600 2123.750 620.740 ;
        RECT 2123.430 620.540 2123.750 620.600 ;
        RECT 2123.445 572.800 2123.735 572.845 ;
        RECT 2123.890 572.800 2124.210 572.860 ;
        RECT 2123.445 572.660 2124.210 572.800 ;
        RECT 2123.445 572.615 2123.735 572.660 ;
        RECT 2123.890 572.600 2124.210 572.660 ;
        RECT 2123.445 535.400 2123.735 535.445 ;
        RECT 2123.890 535.400 2124.210 535.460 ;
        RECT 2123.445 535.260 2124.210 535.400 ;
        RECT 2123.445 535.215 2123.735 535.260 ;
        RECT 2123.890 535.200 2124.210 535.260 ;
        RECT 2123.430 496.640 2123.750 496.700 ;
        RECT 2123.235 496.500 2123.750 496.640 ;
        RECT 2123.430 496.440 2123.750 496.500 ;
        RECT 2123.430 434.760 2123.750 434.820 ;
        RECT 2123.235 434.620 2123.750 434.760 ;
        RECT 2123.430 434.560 2123.750 434.620 ;
        RECT 2123.445 386.480 2123.735 386.525 ;
        RECT 2123.890 386.480 2124.210 386.540 ;
        RECT 2123.445 386.340 2124.210 386.480 ;
        RECT 2123.445 386.295 2123.735 386.340 ;
        RECT 2123.890 386.280 2124.210 386.340 ;
        RECT 2123.430 337.860 2123.750 337.920 ;
        RECT 2123.235 337.720 2123.750 337.860 ;
        RECT 2123.430 337.660 2123.750 337.720 ;
        RECT 2123.445 289.920 2123.735 289.965 ;
        RECT 2123.890 289.920 2124.210 289.980 ;
        RECT 2123.445 289.780 2124.210 289.920 ;
        RECT 2123.445 289.735 2123.735 289.780 ;
        RECT 2123.890 289.720 2124.210 289.780 ;
        RECT 2123.430 241.300 2123.750 241.360 ;
        RECT 2123.235 241.160 2123.750 241.300 ;
        RECT 2123.430 241.100 2123.750 241.160 ;
        RECT 2123.445 193.360 2123.735 193.405 ;
        RECT 2123.890 193.360 2124.210 193.420 ;
        RECT 2123.445 193.220 2124.210 193.360 ;
        RECT 2123.445 193.175 2123.735 193.220 ;
        RECT 2123.890 193.160 2124.210 193.220 ;
        RECT 2123.890 159.020 2124.210 159.080 ;
        RECT 2124.810 159.020 2125.130 159.080 ;
        RECT 2123.890 158.880 2125.130 159.020 ;
        RECT 2123.890 158.820 2124.210 158.880 ;
        RECT 2124.810 158.820 2125.130 158.880 ;
        RECT 2123.890 62.460 2124.210 62.520 ;
        RECT 2124.810 62.460 2125.130 62.520 ;
        RECT 2123.890 62.320 2125.130 62.460 ;
        RECT 2123.890 62.260 2124.210 62.320 ;
        RECT 2124.810 62.260 2125.130 62.320 ;
        RECT 2123.890 23.360 2124.210 23.420 ;
        RECT 2667.150 23.360 2667.470 23.420 ;
        RECT 2123.890 23.220 2667.470 23.360 ;
        RECT 2123.890 23.160 2124.210 23.220 ;
        RECT 2667.150 23.160 2667.470 23.220 ;
      LAYER via ;
        RECT 2119.780 1207.380 2120.040 1207.640 ;
        RECT 2123.920 1207.380 2124.180 1207.640 ;
        RECT 2123.460 1111.160 2123.720 1111.420 ;
        RECT 2123.920 1111.160 2124.180 1111.420 ;
        RECT 2123.460 1110.480 2123.720 1110.740 ;
        RECT 2123.920 1062.540 2124.180 1062.800 ;
        RECT 2123.000 1014.260 2123.260 1014.520 ;
        RECT 2123.460 1014.260 2123.720 1014.520 ;
        RECT 2122.540 965.980 2122.800 966.240 ;
        RECT 2123.920 965.980 2124.180 966.240 ;
        RECT 2123.000 917.700 2123.260 917.960 ;
        RECT 2123.460 917.700 2123.720 917.960 ;
        RECT 2122.540 910.560 2122.800 910.820 ;
        RECT 2123.460 869.080 2123.720 869.340 ;
        RECT 2123.460 862.280 2123.720 862.540 ;
        RECT 2124.840 862.280 2125.100 862.540 ;
        RECT 2123.460 814.000 2123.720 814.260 ;
        RECT 2123.460 786.460 2123.720 786.720 ;
        RECT 2123.460 765.720 2123.720 765.980 ;
        RECT 2123.920 765.720 2124.180 765.980 ;
        RECT 2123.460 717.440 2123.720 717.700 ;
        RECT 2123.460 689.560 2123.720 689.820 ;
        RECT 2123.920 669.160 2124.180 669.420 ;
        RECT 2123.460 621.220 2123.720 621.480 ;
        RECT 2123.460 620.540 2123.720 620.800 ;
        RECT 2123.920 572.600 2124.180 572.860 ;
        RECT 2123.920 535.200 2124.180 535.460 ;
        RECT 2123.460 496.440 2123.720 496.700 ;
        RECT 2123.460 434.560 2123.720 434.820 ;
        RECT 2123.920 386.280 2124.180 386.540 ;
        RECT 2123.460 337.660 2123.720 337.920 ;
        RECT 2123.920 289.720 2124.180 289.980 ;
        RECT 2123.460 241.100 2123.720 241.360 ;
        RECT 2123.920 193.160 2124.180 193.420 ;
        RECT 2123.920 158.820 2124.180 159.080 ;
        RECT 2124.840 158.820 2125.100 159.080 ;
        RECT 2123.920 62.260 2124.180 62.520 ;
        RECT 2124.840 62.260 2125.100 62.520 ;
        RECT 2123.920 23.160 2124.180 23.420 ;
        RECT 2667.180 23.160 2667.440 23.420 ;
      LAYER met2 ;
        RECT 2119.790 1219.680 2120.350 1228.680 ;
        RECT 2119.840 1207.670 2119.980 1219.680 ;
        RECT 2119.780 1207.350 2120.040 1207.670 ;
        RECT 2123.920 1207.350 2124.180 1207.670 ;
        RECT 2123.980 1111.450 2124.120 1207.350 ;
        RECT 2123.460 1111.130 2123.720 1111.450 ;
        RECT 2123.920 1111.130 2124.180 1111.450 ;
        RECT 2123.520 1110.770 2123.660 1111.130 ;
        RECT 2123.460 1110.450 2123.720 1110.770 ;
        RECT 2123.920 1062.685 2124.180 1062.830 ;
        RECT 2122.990 1062.315 2123.270 1062.685 ;
        RECT 2123.910 1062.315 2124.190 1062.685 ;
        RECT 2123.060 1014.550 2123.200 1062.315 ;
        RECT 2122.530 1014.035 2122.810 1014.405 ;
        RECT 2123.000 1014.230 2123.260 1014.550 ;
        RECT 2123.460 1014.405 2123.720 1014.550 ;
        RECT 2123.450 1014.035 2123.730 1014.405 ;
        RECT 2122.600 966.270 2122.740 1014.035 ;
        RECT 2122.540 965.950 2122.800 966.270 ;
        RECT 2123.920 966.125 2124.180 966.270 ;
        RECT 2122.990 965.755 2123.270 966.125 ;
        RECT 2123.910 965.755 2124.190 966.125 ;
        RECT 2123.060 917.990 2123.200 965.755 ;
        RECT 2122.530 917.475 2122.810 917.845 ;
        RECT 2123.000 917.670 2123.260 917.990 ;
        RECT 2123.460 917.845 2123.720 917.990 ;
        RECT 2123.450 917.475 2123.730 917.845 ;
        RECT 2122.600 910.850 2122.740 917.475 ;
        RECT 2122.540 910.530 2122.800 910.850 ;
        RECT 2123.460 869.050 2123.720 869.370 ;
        RECT 2123.520 862.570 2123.660 869.050 ;
        RECT 2123.460 862.250 2123.720 862.570 ;
        RECT 2124.840 862.250 2125.100 862.570 ;
        RECT 2124.900 814.485 2125.040 862.250 ;
        RECT 2123.910 814.370 2124.190 814.485 ;
        RECT 2123.520 814.290 2124.190 814.370 ;
        RECT 2123.460 814.230 2124.190 814.290 ;
        RECT 2123.460 813.970 2123.720 814.230 ;
        RECT 2123.910 814.115 2124.190 814.230 ;
        RECT 2124.830 814.115 2125.110 814.485 ;
        RECT 2123.460 786.430 2123.720 786.750 ;
        RECT 2123.520 766.090 2123.660 786.430 ;
        RECT 2123.520 766.010 2124.120 766.090 ;
        RECT 2123.460 765.950 2124.180 766.010 ;
        RECT 2123.460 765.690 2123.720 765.950 ;
        RECT 2123.920 765.690 2124.180 765.950 ;
        RECT 2123.520 717.730 2123.660 765.690 ;
        RECT 2123.980 765.535 2124.120 765.690 ;
        RECT 2123.460 717.410 2123.720 717.730 ;
        RECT 2123.460 689.530 2123.720 689.850 ;
        RECT 2123.520 669.530 2123.660 689.530 ;
        RECT 2123.520 669.450 2124.120 669.530 ;
        RECT 2123.520 669.390 2124.180 669.450 ;
        RECT 2123.920 669.130 2124.180 669.390 ;
        RECT 2123.980 668.975 2124.120 669.130 ;
        RECT 2123.460 621.190 2123.720 621.510 ;
        RECT 2123.520 620.830 2123.660 621.190 ;
        RECT 2123.460 620.510 2123.720 620.830 ;
        RECT 2123.920 572.570 2124.180 572.890 ;
        RECT 2123.980 535.490 2124.120 572.570 ;
        RECT 2123.920 535.170 2124.180 535.490 ;
        RECT 2123.460 496.410 2123.720 496.730 ;
        RECT 2123.520 483.210 2123.660 496.410 ;
        RECT 2123.520 483.070 2124.120 483.210 ;
        RECT 2123.980 434.930 2124.120 483.070 ;
        RECT 2123.520 434.850 2124.120 434.930 ;
        RECT 2123.460 434.790 2124.120 434.850 ;
        RECT 2123.460 434.530 2123.720 434.790 ;
        RECT 2123.920 386.250 2124.180 386.570 ;
        RECT 2123.980 339.165 2124.120 386.250 ;
        RECT 2123.910 338.795 2124.190 339.165 ;
        RECT 2123.450 338.115 2123.730 338.485 ;
        RECT 2123.520 337.950 2123.660 338.115 ;
        RECT 2123.460 337.630 2123.720 337.950 ;
        RECT 2123.920 289.690 2124.180 290.010 ;
        RECT 2123.980 265.610 2124.120 289.690 ;
        RECT 2123.520 265.470 2124.120 265.610 ;
        RECT 2123.520 241.390 2123.660 265.470 ;
        RECT 2123.460 241.070 2123.720 241.390 ;
        RECT 2123.920 193.130 2124.180 193.450 ;
        RECT 2123.980 159.110 2124.120 193.130 ;
        RECT 2123.920 158.790 2124.180 159.110 ;
        RECT 2124.840 158.790 2125.100 159.110 ;
        RECT 2124.900 62.550 2125.040 158.790 ;
        RECT 2123.920 62.230 2124.180 62.550 ;
        RECT 2124.840 62.230 2125.100 62.550 ;
        RECT 2123.980 23.450 2124.120 62.230 ;
        RECT 2123.920 23.130 2124.180 23.450 ;
        RECT 2667.180 23.130 2667.440 23.450 ;
        RECT 2667.240 2.400 2667.380 23.130 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
      LAYER via2 ;
        RECT 2122.990 1062.360 2123.270 1062.640 ;
        RECT 2123.910 1062.360 2124.190 1062.640 ;
        RECT 2122.530 1014.080 2122.810 1014.360 ;
        RECT 2123.450 1014.080 2123.730 1014.360 ;
        RECT 2122.990 965.800 2123.270 966.080 ;
        RECT 2123.910 965.800 2124.190 966.080 ;
        RECT 2122.530 917.520 2122.810 917.800 ;
        RECT 2123.450 917.520 2123.730 917.800 ;
        RECT 2123.910 814.160 2124.190 814.440 ;
        RECT 2124.830 814.160 2125.110 814.440 ;
        RECT 2123.910 338.840 2124.190 339.120 ;
        RECT 2123.450 338.160 2123.730 338.440 ;
      LAYER met3 ;
        RECT 2122.965 1062.650 2123.295 1062.665 ;
        RECT 2123.885 1062.650 2124.215 1062.665 ;
        RECT 2122.965 1062.350 2124.215 1062.650 ;
        RECT 2122.965 1062.335 2123.295 1062.350 ;
        RECT 2123.885 1062.335 2124.215 1062.350 ;
        RECT 2122.505 1014.370 2122.835 1014.385 ;
        RECT 2123.425 1014.370 2123.755 1014.385 ;
        RECT 2122.505 1014.070 2123.755 1014.370 ;
        RECT 2122.505 1014.055 2122.835 1014.070 ;
        RECT 2123.425 1014.055 2123.755 1014.070 ;
        RECT 2122.965 966.090 2123.295 966.105 ;
        RECT 2123.885 966.090 2124.215 966.105 ;
        RECT 2122.965 965.790 2124.215 966.090 ;
        RECT 2122.965 965.775 2123.295 965.790 ;
        RECT 2123.885 965.775 2124.215 965.790 ;
        RECT 2122.505 917.810 2122.835 917.825 ;
        RECT 2123.425 917.810 2123.755 917.825 ;
        RECT 2122.505 917.510 2123.755 917.810 ;
        RECT 2122.505 917.495 2122.835 917.510 ;
        RECT 2123.425 917.495 2123.755 917.510 ;
        RECT 2123.885 814.450 2124.215 814.465 ;
        RECT 2124.805 814.450 2125.135 814.465 ;
        RECT 2123.885 814.150 2125.135 814.450 ;
        RECT 2123.885 814.135 2124.215 814.150 ;
        RECT 2124.805 814.135 2125.135 814.150 ;
        RECT 2123.885 339.130 2124.215 339.145 ;
        RECT 2122.750 338.830 2124.215 339.130 ;
        RECT 2122.750 338.450 2123.050 338.830 ;
        RECT 2123.885 338.815 2124.215 338.830 ;
        RECT 2123.425 338.450 2123.755 338.465 ;
        RECT 2122.750 338.150 2123.755 338.450 ;
        RECT 2123.425 338.135 2123.755 338.150 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2162.605 23.715 2162.775 26.095 ;
        RECT 2162.605 23.545 2163.695 23.715 ;
      LAYER mcon ;
        RECT 2162.605 25.925 2162.775 26.095 ;
        RECT 2163.525 23.545 2163.695 23.715 ;
      LAYER met1 ;
        RECT 2128.950 1207.580 2129.270 1207.640 ;
        RECT 2131.710 1207.580 2132.030 1207.640 ;
        RECT 2128.950 1207.440 2132.030 1207.580 ;
        RECT 2128.950 1207.380 2129.270 1207.440 ;
        RECT 2131.710 1207.380 2132.030 1207.440 ;
        RECT 2131.710 26.080 2132.030 26.140 ;
        RECT 2162.545 26.080 2162.835 26.125 ;
        RECT 2131.710 25.940 2162.835 26.080 ;
        RECT 2131.710 25.880 2132.030 25.940 ;
        RECT 2162.545 25.895 2162.835 25.940 ;
        RECT 2163.465 23.700 2163.755 23.745 ;
        RECT 2684.630 23.700 2684.950 23.760 ;
        RECT 2163.465 23.560 2684.950 23.700 ;
        RECT 2163.465 23.515 2163.755 23.560 ;
        RECT 2684.630 23.500 2684.950 23.560 ;
      LAYER via ;
        RECT 2128.980 1207.380 2129.240 1207.640 ;
        RECT 2131.740 1207.380 2132.000 1207.640 ;
        RECT 2131.740 25.880 2132.000 26.140 ;
        RECT 2684.660 23.500 2684.920 23.760 ;
      LAYER met2 ;
        RECT 2128.990 1219.680 2129.550 1228.680 ;
        RECT 2129.040 1207.670 2129.180 1219.680 ;
        RECT 2128.980 1207.350 2129.240 1207.670 ;
        RECT 2131.740 1207.350 2132.000 1207.670 ;
        RECT 2131.800 26.170 2131.940 1207.350 ;
        RECT 2131.740 25.850 2132.000 26.170 ;
        RECT 2684.660 23.470 2684.920 23.790 ;
        RECT 2684.720 2.400 2684.860 23.470 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2162.990 27.440 2163.310 27.500 ;
        RECT 2702.570 27.440 2702.890 27.500 ;
        RECT 2162.990 27.300 2702.890 27.440 ;
        RECT 2162.990 27.240 2163.310 27.300 ;
        RECT 2702.570 27.240 2702.890 27.300 ;
        RECT 2138.150 25.740 2138.470 25.800 ;
        RECT 2162.990 25.740 2163.310 25.800 ;
        RECT 2138.150 25.600 2163.310 25.740 ;
        RECT 2138.150 25.540 2138.470 25.600 ;
        RECT 2162.990 25.540 2163.310 25.600 ;
      LAYER via ;
        RECT 2163.020 27.240 2163.280 27.500 ;
        RECT 2702.600 27.240 2702.860 27.500 ;
        RECT 2138.180 25.540 2138.440 25.800 ;
        RECT 2163.020 25.540 2163.280 25.800 ;
      LAYER met2 ;
        RECT 2138.190 1219.680 2138.750 1228.680 ;
        RECT 2138.240 25.830 2138.380 1219.680 ;
        RECT 2163.020 27.210 2163.280 27.530 ;
        RECT 2702.600 27.210 2702.860 27.530 ;
        RECT 2163.080 25.830 2163.220 27.210 ;
        RECT 2138.180 25.510 2138.440 25.830 ;
        RECT 2163.020 25.510 2163.280 25.830 ;
        RECT 2702.660 2.400 2702.800 27.210 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2147.350 1207.580 2147.670 1207.640 ;
        RECT 2152.410 1207.580 2152.730 1207.640 ;
        RECT 2147.350 1207.440 2152.730 1207.580 ;
        RECT 2147.350 1207.380 2147.670 1207.440 ;
        RECT 2152.410 1207.380 2152.730 1207.440 ;
        RECT 2720.510 27.100 2720.830 27.160 ;
        RECT 2164.460 26.960 2720.830 27.100 ;
        RECT 2152.410 26.760 2152.730 26.820 ;
        RECT 2164.460 26.760 2164.600 26.960 ;
        RECT 2720.510 26.900 2720.830 26.960 ;
        RECT 2152.410 26.620 2164.600 26.760 ;
        RECT 2152.410 26.560 2152.730 26.620 ;
      LAYER via ;
        RECT 2147.380 1207.380 2147.640 1207.640 ;
        RECT 2152.440 1207.380 2152.700 1207.640 ;
        RECT 2152.440 26.560 2152.700 26.820 ;
        RECT 2720.540 26.900 2720.800 27.160 ;
      LAYER met2 ;
        RECT 2147.390 1219.680 2147.950 1228.680 ;
        RECT 2147.440 1207.670 2147.580 1219.680 ;
        RECT 2147.380 1207.350 2147.640 1207.670 ;
        RECT 2152.440 1207.350 2152.700 1207.670 ;
        RECT 2152.500 26.850 2152.640 1207.350 ;
        RECT 2720.540 26.870 2720.800 27.190 ;
        RECT 2152.440 26.530 2152.700 26.850 ;
        RECT 2720.600 2.400 2720.740 26.870 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2162.145 26.945 2163.235 27.115 ;
        RECT 2163.065 26.095 2163.235 26.945 ;
        RECT 2163.065 25.925 2164.615 26.095 ;
        RECT 2185.605 24.905 2185.775 26.095 ;
        RECT 2191.585 24.225 2191.755 25.075 ;
        RECT 2207.685 24.225 2207.855 26.775 ;
      LAYER mcon ;
        RECT 2207.685 26.605 2207.855 26.775 ;
        RECT 2164.445 25.925 2164.615 26.095 ;
        RECT 2185.605 25.925 2185.775 26.095 ;
        RECT 2191.585 24.905 2191.755 25.075 ;
      LAYER met1 ;
        RECT 2158.850 27.100 2159.170 27.160 ;
        RECT 2162.085 27.100 2162.375 27.145 ;
        RECT 2158.850 26.960 2162.375 27.100 ;
        RECT 2158.850 26.900 2159.170 26.960 ;
        RECT 2162.085 26.915 2162.375 26.960 ;
        RECT 2207.625 26.760 2207.915 26.805 ;
        RECT 2738.450 26.760 2738.770 26.820 ;
        RECT 2207.625 26.620 2738.770 26.760 ;
        RECT 2207.625 26.575 2207.915 26.620 ;
        RECT 2738.450 26.560 2738.770 26.620 ;
        RECT 2164.385 26.080 2164.675 26.125 ;
        RECT 2185.545 26.080 2185.835 26.125 ;
        RECT 2164.385 25.940 2185.835 26.080 ;
        RECT 2164.385 25.895 2164.675 25.940 ;
        RECT 2185.545 25.895 2185.835 25.940 ;
        RECT 2185.545 25.060 2185.835 25.105 ;
        RECT 2191.525 25.060 2191.815 25.105 ;
        RECT 2185.545 24.920 2191.815 25.060 ;
        RECT 2185.545 24.875 2185.835 24.920 ;
        RECT 2191.525 24.875 2191.815 24.920 ;
        RECT 2191.525 24.380 2191.815 24.425 ;
        RECT 2207.625 24.380 2207.915 24.425 ;
        RECT 2191.525 24.240 2207.915 24.380 ;
        RECT 2191.525 24.195 2191.815 24.240 ;
        RECT 2207.625 24.195 2207.915 24.240 ;
      LAYER via ;
        RECT 2158.880 26.900 2159.140 27.160 ;
        RECT 2738.480 26.560 2738.740 26.820 ;
      LAYER met2 ;
        RECT 2156.590 1220.330 2157.150 1228.680 ;
        RECT 2156.590 1220.190 2159.080 1220.330 ;
        RECT 2156.590 1219.680 2157.150 1220.190 ;
        RECT 2158.940 27.190 2159.080 1220.190 ;
        RECT 2158.880 26.870 2159.140 27.190 ;
        RECT 2738.480 26.530 2738.740 26.850 ;
        RECT 2738.540 2.400 2738.680 26.530 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 26.760 2166.530 26.820 ;
        RECT 2166.210 26.620 2168.740 26.760 ;
        RECT 2166.210 26.560 2166.530 26.620 ;
        RECT 2168.600 26.420 2168.740 26.620 ;
        RECT 2755.930 26.420 2756.250 26.480 ;
        RECT 2168.600 26.280 2756.250 26.420 ;
        RECT 2755.930 26.220 2756.250 26.280 ;
      LAYER via ;
        RECT 2166.240 26.560 2166.500 26.820 ;
        RECT 2755.960 26.220 2756.220 26.480 ;
      LAYER met2 ;
        RECT 2165.790 1220.330 2166.350 1228.680 ;
        RECT 2165.790 1219.680 2166.440 1220.330 ;
        RECT 2166.300 26.850 2166.440 1219.680 ;
        RECT 2166.240 26.530 2166.500 26.850 ;
        RECT 2755.960 26.190 2756.220 26.510 ;
        RECT 2756.020 2.400 2756.160 26.190 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 829.450 17.240 829.770 17.300 ;
        RECT 1173.070 17.240 1173.390 17.300 ;
        RECT 829.450 17.100 1173.390 17.240 ;
        RECT 829.450 17.040 829.770 17.100 ;
        RECT 1173.070 17.040 1173.390 17.100 ;
      LAYER via ;
        RECT 829.480 17.040 829.740 17.300 ;
        RECT 1173.100 17.040 1173.360 17.300 ;
      LAYER met2 ;
        RECT 1175.870 1221.010 1176.430 1228.680 ;
        RECT 1173.620 1220.870 1176.430 1221.010 ;
        RECT 1173.620 1196.700 1173.760 1220.870 ;
        RECT 1175.870 1219.680 1176.430 1220.870 ;
        RECT 1173.160 1196.560 1173.760 1196.700 ;
        RECT 1173.160 17.330 1173.300 1196.560 ;
        RECT 829.480 17.010 829.740 17.330 ;
        RECT 1173.100 17.010 1173.360 17.330 ;
        RECT 829.540 2.400 829.680 17.010 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2203.545 24.565 2203.715 25.755 ;
        RECT 2232.525 24.565 2232.695 26.095 ;
      LAYER mcon ;
        RECT 2232.525 25.925 2232.695 26.095 ;
        RECT 2203.545 25.585 2203.715 25.755 ;
      LAYER met1 ;
        RECT 2174.490 1207.580 2174.810 1207.640 ;
        RECT 2180.010 1207.580 2180.330 1207.640 ;
        RECT 2174.490 1207.440 2180.330 1207.580 ;
        RECT 2174.490 1207.380 2174.810 1207.440 ;
        RECT 2180.010 1207.380 2180.330 1207.440 ;
        RECT 2232.465 26.080 2232.755 26.125 ;
        RECT 2773.870 26.080 2774.190 26.140 ;
        RECT 2232.465 25.940 2774.190 26.080 ;
        RECT 2232.465 25.895 2232.755 25.940 ;
        RECT 2773.870 25.880 2774.190 25.940 ;
        RECT 2180.010 25.740 2180.330 25.800 ;
        RECT 2203.485 25.740 2203.775 25.785 ;
        RECT 2180.010 25.600 2203.775 25.740 ;
        RECT 2180.010 25.540 2180.330 25.600 ;
        RECT 2203.485 25.555 2203.775 25.600 ;
        RECT 2203.485 24.720 2203.775 24.765 ;
        RECT 2232.465 24.720 2232.755 24.765 ;
        RECT 2203.485 24.580 2232.755 24.720 ;
        RECT 2203.485 24.535 2203.775 24.580 ;
        RECT 2232.465 24.535 2232.755 24.580 ;
      LAYER via ;
        RECT 2174.520 1207.380 2174.780 1207.640 ;
        RECT 2180.040 1207.380 2180.300 1207.640 ;
        RECT 2773.900 25.880 2774.160 26.140 ;
        RECT 2180.040 25.540 2180.300 25.800 ;
      LAYER met2 ;
        RECT 2174.530 1219.680 2175.090 1228.680 ;
        RECT 2174.580 1207.670 2174.720 1219.680 ;
        RECT 2174.520 1207.350 2174.780 1207.670 ;
        RECT 2180.040 1207.350 2180.300 1207.670 ;
        RECT 2180.100 25.830 2180.240 1207.350 ;
        RECT 2773.900 25.850 2774.160 26.170 ;
        RECT 2180.040 25.510 2180.300 25.830 ;
        RECT 2773.960 2.400 2774.100 25.850 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2183.690 1207.580 2184.010 1207.640 ;
        RECT 2186.910 1207.580 2187.230 1207.640 ;
        RECT 2183.690 1207.440 2187.230 1207.580 ;
        RECT 2183.690 1207.380 2184.010 1207.440 ;
        RECT 2186.910 1207.380 2187.230 1207.440 ;
        RECT 2186.910 26.080 2187.230 26.140 ;
        RECT 2186.910 25.940 2232.220 26.080 ;
        RECT 2186.910 25.880 2187.230 25.940 ;
        RECT 2232.080 25.740 2232.220 25.940 ;
        RECT 2791.810 25.740 2792.130 25.800 ;
        RECT 2232.080 25.600 2792.130 25.740 ;
        RECT 2791.810 25.540 2792.130 25.600 ;
      LAYER via ;
        RECT 2183.720 1207.380 2183.980 1207.640 ;
        RECT 2186.940 1207.380 2187.200 1207.640 ;
        RECT 2186.940 25.880 2187.200 26.140 ;
        RECT 2791.840 25.540 2792.100 25.800 ;
      LAYER met2 ;
        RECT 2183.730 1219.680 2184.290 1228.680 ;
        RECT 2183.780 1207.670 2183.920 1219.680 ;
        RECT 2183.720 1207.350 2183.980 1207.670 ;
        RECT 2186.940 1207.350 2187.200 1207.670 ;
        RECT 2187.000 26.170 2187.140 1207.350 ;
        RECT 2186.940 25.850 2187.200 26.170 ;
        RECT 2791.840 25.510 2792.100 25.830 ;
        RECT 2791.900 2.400 2792.040 25.510 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2193.350 25.060 2193.670 25.120 ;
        RECT 2809.750 25.060 2810.070 25.120 ;
        RECT 2193.350 24.920 2810.070 25.060 ;
        RECT 2193.350 24.860 2193.670 24.920 ;
        RECT 2809.750 24.860 2810.070 24.920 ;
      LAYER via ;
        RECT 2193.380 24.860 2193.640 25.120 ;
        RECT 2809.780 24.860 2810.040 25.120 ;
      LAYER met2 ;
        RECT 2192.930 1220.330 2193.490 1228.680 ;
        RECT 2192.930 1219.680 2193.580 1220.330 ;
        RECT 2193.440 25.150 2193.580 1219.680 ;
        RECT 2193.380 24.830 2193.640 25.150 ;
        RECT 2809.780 24.830 2810.040 25.150 ;
        RECT 2809.840 2.400 2809.980 24.830 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2202.090 1210.640 2202.410 1210.700 ;
        RECT 2207.610 1210.640 2207.930 1210.700 ;
        RECT 2202.090 1210.500 2207.930 1210.640 ;
        RECT 2202.090 1210.440 2202.410 1210.500 ;
        RECT 2207.610 1210.440 2207.930 1210.500 ;
        RECT 2207.610 25.740 2207.930 25.800 ;
        RECT 2207.610 25.600 2231.760 25.740 ;
        RECT 2207.610 25.540 2207.930 25.600 ;
        RECT 2231.620 25.400 2231.760 25.600 ;
        RECT 2827.690 25.400 2828.010 25.460 ;
        RECT 2231.620 25.260 2828.010 25.400 ;
        RECT 2827.690 25.200 2828.010 25.260 ;
      LAYER via ;
        RECT 2202.120 1210.440 2202.380 1210.700 ;
        RECT 2207.640 1210.440 2207.900 1210.700 ;
        RECT 2207.640 25.540 2207.900 25.800 ;
        RECT 2827.720 25.200 2827.980 25.460 ;
      LAYER met2 ;
        RECT 2202.130 1219.680 2202.690 1228.680 ;
        RECT 2202.180 1210.730 2202.320 1219.680 ;
        RECT 2202.120 1210.410 2202.380 1210.730 ;
        RECT 2207.640 1210.410 2207.900 1210.730 ;
        RECT 2207.700 25.830 2207.840 1210.410 ;
        RECT 2207.640 25.510 2207.900 25.830 ;
        RECT 2827.720 25.170 2827.980 25.490 ;
        RECT 2827.780 2.400 2827.920 25.170 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2232.985 23.885 2233.155 24.735 ;
      LAYER mcon ;
        RECT 2232.985 24.565 2233.155 24.735 ;
      LAYER met1 ;
        RECT 2232.925 24.720 2233.215 24.765 ;
        RECT 2845.170 24.720 2845.490 24.780 ;
        RECT 2232.925 24.580 2845.490 24.720 ;
        RECT 2232.925 24.535 2233.215 24.580 ;
        RECT 2845.170 24.520 2845.490 24.580 ;
        RECT 2214.050 24.040 2214.370 24.100 ;
        RECT 2232.925 24.040 2233.215 24.085 ;
        RECT 2214.050 23.900 2233.215 24.040 ;
        RECT 2214.050 23.840 2214.370 23.900 ;
        RECT 2232.925 23.855 2233.215 23.900 ;
      LAYER via ;
        RECT 2845.200 24.520 2845.460 24.780 ;
        RECT 2214.080 23.840 2214.340 24.100 ;
      LAYER met2 ;
        RECT 2211.330 1220.330 2211.890 1228.680 ;
        RECT 2211.330 1220.190 2214.280 1220.330 ;
        RECT 2211.330 1219.680 2211.890 1220.190 ;
        RECT 2214.140 24.130 2214.280 1220.190 ;
        RECT 2845.200 24.490 2845.460 24.810 ;
        RECT 2214.080 23.810 2214.340 24.130 ;
        RECT 2845.260 2.400 2845.400 24.490 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2221.410 24.380 2221.730 24.440 ;
        RECT 2863.110 24.380 2863.430 24.440 ;
        RECT 2221.410 24.240 2863.430 24.380 ;
        RECT 2221.410 24.180 2221.730 24.240 ;
        RECT 2863.110 24.180 2863.430 24.240 ;
      LAYER via ;
        RECT 2221.440 24.180 2221.700 24.440 ;
        RECT 2863.140 24.180 2863.400 24.440 ;
      LAYER met2 ;
        RECT 2220.530 1220.330 2221.090 1228.680 ;
        RECT 2220.530 1220.190 2221.640 1220.330 ;
        RECT 2220.530 1219.680 2221.090 1220.190 ;
        RECT 2221.500 24.470 2221.640 1220.190 ;
        RECT 2221.440 24.150 2221.700 24.470 ;
        RECT 2863.140 24.150 2863.400 24.470 ;
        RECT 2863.200 2.400 2863.340 24.150 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2229.690 1210.300 2230.010 1210.360 ;
        RECT 2235.210 1210.300 2235.530 1210.360 ;
        RECT 2229.690 1210.160 2235.530 1210.300 ;
        RECT 2229.690 1210.100 2230.010 1210.160 ;
        RECT 2235.210 1210.100 2235.530 1210.160 ;
        RECT 2235.210 24.040 2235.530 24.100 ;
        RECT 2881.050 24.040 2881.370 24.100 ;
        RECT 2235.210 23.900 2881.370 24.040 ;
        RECT 2235.210 23.840 2235.530 23.900 ;
        RECT 2881.050 23.840 2881.370 23.900 ;
      LAYER via ;
        RECT 2229.720 1210.100 2229.980 1210.360 ;
        RECT 2235.240 1210.100 2235.500 1210.360 ;
        RECT 2235.240 23.840 2235.500 24.100 ;
        RECT 2881.080 23.840 2881.340 24.100 ;
      LAYER met2 ;
        RECT 2229.730 1219.680 2230.290 1228.680 ;
        RECT 2229.780 1210.390 2229.920 1219.680 ;
        RECT 2229.720 1210.070 2229.980 1210.390 ;
        RECT 2235.240 1210.070 2235.500 1210.390 ;
        RECT 2235.300 24.130 2235.440 1210.070 ;
        RECT 2235.240 23.810 2235.500 24.130 ;
        RECT 2881.080 23.810 2881.340 24.130 ;
        RECT 2881.140 2.400 2881.280 23.810 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2238.890 1210.300 2239.210 1210.360 ;
        RECT 2242.110 1210.300 2242.430 1210.360 ;
        RECT 2238.890 1210.160 2242.430 1210.300 ;
        RECT 2238.890 1210.100 2239.210 1210.160 ;
        RECT 2242.110 1210.100 2242.430 1210.160 ;
      LAYER via ;
        RECT 2238.920 1210.100 2239.180 1210.360 ;
        RECT 2242.140 1210.100 2242.400 1210.360 ;
      LAYER met2 ;
        RECT 2238.930 1219.680 2239.490 1228.680 ;
        RECT 2238.980 1210.390 2239.120 1219.680 ;
        RECT 2238.920 1210.070 2239.180 1210.390 ;
        RECT 2242.140 1210.070 2242.400 1210.390 ;
        RECT 2242.200 24.325 2242.340 1210.070 ;
        RECT 2242.130 23.955 2242.410 24.325 ;
        RECT 2899.010 23.955 2899.290 24.325 ;
        RECT 2899.080 2.400 2899.220 23.955 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 2242.130 24.000 2242.410 24.280 ;
        RECT 2899.010 24.000 2899.290 24.280 ;
      LAYER met3 ;
        RECT 2242.105 24.290 2242.435 24.305 ;
        RECT 2898.985 24.290 2899.315 24.305 ;
        RECT 2242.105 23.990 2899.315 24.290 ;
        RECT 2242.105 23.975 2242.435 23.990 ;
        RECT 2898.985 23.975 2899.315 23.990 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1181.425 786.165 1181.595 821.015 ;
        RECT 1131.745 17.425 1131.915 18.275 ;
      LAYER mcon ;
        RECT 1181.425 820.845 1181.595 821.015 ;
        RECT 1131.745 18.105 1131.915 18.275 ;
      LAYER met1 ;
        RECT 1181.810 1159.300 1182.130 1159.360 ;
        RECT 1182.730 1159.300 1183.050 1159.360 ;
        RECT 1181.810 1159.160 1183.050 1159.300 ;
        RECT 1181.810 1159.100 1182.130 1159.160 ;
        RECT 1182.730 1159.100 1183.050 1159.160 ;
        RECT 1181.350 966.180 1181.670 966.240 ;
        RECT 1182.270 966.180 1182.590 966.240 ;
        RECT 1181.350 966.040 1182.590 966.180 ;
        RECT 1181.350 965.980 1181.670 966.040 ;
        RECT 1182.270 965.980 1182.590 966.040 ;
        RECT 1181.350 869.620 1181.670 869.680 ;
        RECT 1182.270 869.620 1182.590 869.680 ;
        RECT 1181.350 869.480 1182.590 869.620 ;
        RECT 1181.350 869.420 1181.670 869.480 ;
        RECT 1182.270 869.420 1182.590 869.480 ;
        RECT 1181.350 821.000 1181.670 821.060 ;
        RECT 1181.155 820.860 1181.670 821.000 ;
        RECT 1181.350 820.800 1181.670 820.860 ;
        RECT 1181.350 786.320 1181.670 786.380 ;
        RECT 1181.155 786.180 1181.670 786.320 ;
        RECT 1181.350 786.120 1181.670 786.180 ;
        RECT 1181.350 724.440 1181.670 724.500 ;
        RECT 1181.810 724.440 1182.130 724.500 ;
        RECT 1181.350 724.300 1182.130 724.440 ;
        RECT 1181.350 724.240 1181.670 724.300 ;
        RECT 1181.810 724.240 1182.130 724.300 ;
        RECT 1181.350 579.400 1181.670 579.660 ;
        RECT 1181.440 579.260 1181.580 579.400 ;
        RECT 1181.810 579.260 1182.130 579.320 ;
        RECT 1181.440 579.120 1182.130 579.260 ;
        RECT 1181.810 579.060 1182.130 579.120 ;
        RECT 1180.890 435.100 1181.210 435.160 ;
        RECT 1181.350 435.100 1181.670 435.160 ;
        RECT 1180.890 434.960 1181.670 435.100 ;
        RECT 1180.890 434.900 1181.210 434.960 ;
        RECT 1181.350 434.900 1181.670 434.960 ;
        RECT 1180.890 386.480 1181.210 386.540 ;
        RECT 1181.350 386.480 1181.670 386.540 ;
        RECT 1180.890 386.340 1181.670 386.480 ;
        RECT 1180.890 386.280 1181.210 386.340 ;
        RECT 1181.350 386.280 1181.670 386.340 ;
        RECT 1181.350 337.860 1181.670 337.920 ;
        RECT 1181.810 337.860 1182.130 337.920 ;
        RECT 1181.350 337.720 1182.130 337.860 ;
        RECT 1181.350 337.660 1181.670 337.720 ;
        RECT 1181.810 337.660 1182.130 337.720 ;
        RECT 1181.350 241.300 1181.670 241.360 ;
        RECT 1181.810 241.300 1182.130 241.360 ;
        RECT 1181.350 241.160 1182.130 241.300 ;
        RECT 1181.350 241.100 1181.670 241.160 ;
        RECT 1181.810 241.100 1182.130 241.160 ;
        RECT 1181.350 145.420 1181.670 145.480 ;
        RECT 1180.980 145.280 1181.670 145.420 ;
        RECT 1180.980 145.140 1181.120 145.280 ;
        RECT 1181.350 145.220 1181.670 145.280 ;
        RECT 1180.890 144.880 1181.210 145.140 ;
        RECT 1180.890 96.800 1181.210 96.860 ;
        RECT 1181.350 96.800 1181.670 96.860 ;
        RECT 1180.890 96.660 1181.670 96.800 ;
        RECT 1180.890 96.600 1181.210 96.660 ;
        RECT 1181.350 96.600 1181.670 96.660 ;
        RECT 1131.685 18.260 1131.975 18.305 ;
        RECT 1131.685 18.120 1132.820 18.260 ;
        RECT 1131.685 18.075 1131.975 18.120 ;
        RECT 1132.680 17.920 1132.820 18.120 ;
        RECT 1181.350 17.920 1181.670 17.980 ;
        RECT 1132.680 17.780 1181.670 17.920 ;
        RECT 1181.350 17.720 1181.670 17.780 ;
        RECT 846.930 17.580 847.250 17.640 ;
        RECT 1131.685 17.580 1131.975 17.625 ;
        RECT 846.930 17.440 1131.975 17.580 ;
        RECT 846.930 17.380 847.250 17.440 ;
        RECT 1131.685 17.395 1131.975 17.440 ;
      LAYER via ;
        RECT 1181.840 1159.100 1182.100 1159.360 ;
        RECT 1182.760 1159.100 1183.020 1159.360 ;
        RECT 1181.380 965.980 1181.640 966.240 ;
        RECT 1182.300 965.980 1182.560 966.240 ;
        RECT 1181.380 869.420 1181.640 869.680 ;
        RECT 1182.300 869.420 1182.560 869.680 ;
        RECT 1181.380 820.800 1181.640 821.060 ;
        RECT 1181.380 786.120 1181.640 786.380 ;
        RECT 1181.380 724.240 1181.640 724.500 ;
        RECT 1181.840 724.240 1182.100 724.500 ;
        RECT 1181.380 579.400 1181.640 579.660 ;
        RECT 1181.840 579.060 1182.100 579.320 ;
        RECT 1180.920 434.900 1181.180 435.160 ;
        RECT 1181.380 434.900 1181.640 435.160 ;
        RECT 1180.920 386.280 1181.180 386.540 ;
        RECT 1181.380 386.280 1181.640 386.540 ;
        RECT 1181.380 337.660 1181.640 337.920 ;
        RECT 1181.840 337.660 1182.100 337.920 ;
        RECT 1181.380 241.100 1181.640 241.360 ;
        RECT 1181.840 241.100 1182.100 241.360 ;
        RECT 1181.380 145.220 1181.640 145.480 ;
        RECT 1180.920 144.880 1181.180 145.140 ;
        RECT 1180.920 96.600 1181.180 96.860 ;
        RECT 1181.380 96.600 1181.640 96.860 ;
        RECT 1181.380 17.720 1181.640 17.980 ;
        RECT 846.960 17.380 847.220 17.640 ;
      LAYER met2 ;
        RECT 1185.070 1221.010 1185.630 1228.680 ;
        RECT 1182.820 1220.870 1185.630 1221.010 ;
        RECT 1182.820 1159.390 1182.960 1220.870 ;
        RECT 1185.070 1219.680 1185.630 1220.870 ;
        RECT 1181.840 1159.070 1182.100 1159.390 ;
        RECT 1182.760 1159.070 1183.020 1159.390 ;
        RECT 1181.900 1076.850 1182.040 1159.070 ;
        RECT 1181.440 1076.710 1182.040 1076.850 ;
        RECT 1181.440 1027.890 1181.580 1076.710 ;
        RECT 1181.440 1027.750 1182.040 1027.890 ;
        RECT 1181.900 990.490 1182.040 1027.750 ;
        RECT 1181.900 990.350 1182.500 990.490 ;
        RECT 1182.360 966.270 1182.500 990.350 ;
        RECT 1181.380 965.950 1181.640 966.270 ;
        RECT 1182.300 965.950 1182.560 966.270 ;
        RECT 1181.440 942.210 1181.580 965.950 ;
        RECT 1181.440 942.070 1182.040 942.210 ;
        RECT 1181.900 893.930 1182.040 942.070 ;
        RECT 1181.900 893.790 1182.500 893.930 ;
        RECT 1182.360 869.710 1182.500 893.790 ;
        RECT 1181.380 869.390 1181.640 869.710 ;
        RECT 1182.300 869.390 1182.560 869.710 ;
        RECT 1181.440 821.090 1181.580 869.390 ;
        RECT 1181.380 820.770 1181.640 821.090 ;
        RECT 1181.380 786.090 1181.640 786.410 ;
        RECT 1181.440 748.410 1181.580 786.090 ;
        RECT 1181.440 748.270 1182.040 748.410 ;
        RECT 1181.900 724.530 1182.040 748.270 ;
        RECT 1181.380 724.210 1181.640 724.530 ;
        RECT 1181.840 724.210 1182.100 724.530 ;
        RECT 1181.440 651.850 1181.580 724.210 ;
        RECT 1181.440 651.710 1182.040 651.850 ;
        RECT 1181.900 580.565 1182.040 651.710 ;
        RECT 1181.830 580.195 1182.110 580.565 ;
        RECT 1181.370 579.515 1181.650 579.885 ;
        RECT 1181.380 579.370 1181.640 579.515 ;
        RECT 1181.840 579.030 1182.100 579.350 ;
        RECT 1181.900 507.010 1182.040 579.030 ;
        RECT 1181.440 506.870 1182.040 507.010 ;
        RECT 1181.440 435.190 1181.580 506.870 ;
        RECT 1180.920 434.870 1181.180 435.190 ;
        RECT 1181.380 434.870 1181.640 435.190 ;
        RECT 1180.980 386.570 1181.120 434.870 ;
        RECT 1180.920 386.250 1181.180 386.570 ;
        RECT 1181.380 386.250 1181.640 386.570 ;
        RECT 1181.440 337.950 1181.580 386.250 ;
        RECT 1181.380 337.630 1181.640 337.950 ;
        RECT 1181.840 337.630 1182.100 337.950 ;
        RECT 1181.900 241.390 1182.040 337.630 ;
        RECT 1181.380 241.070 1181.640 241.390 ;
        RECT 1181.840 241.070 1182.100 241.390 ;
        RECT 1181.440 145.510 1181.580 241.070 ;
        RECT 1181.380 145.190 1181.640 145.510 ;
        RECT 1180.920 144.850 1181.180 145.170 ;
        RECT 1180.980 96.890 1181.120 144.850 ;
        RECT 1180.920 96.570 1181.180 96.890 ;
        RECT 1181.380 96.570 1181.640 96.890 ;
        RECT 1181.440 18.010 1181.580 96.570 ;
        RECT 1181.380 17.690 1181.640 18.010 ;
        RECT 846.960 17.350 847.220 17.670 ;
        RECT 847.020 2.400 847.160 17.350 ;
        RECT 846.810 -4.800 847.370 2.400 ;
      LAYER via2 ;
        RECT 1181.830 580.240 1182.110 580.520 ;
        RECT 1181.370 579.560 1181.650 579.840 ;
      LAYER met3 ;
        RECT 1181.805 580.530 1182.135 580.545 ;
        RECT 1181.590 580.215 1182.135 580.530 ;
        RECT 1181.590 579.865 1181.890 580.215 ;
        RECT 1181.345 579.550 1181.890 579.865 ;
        RECT 1181.345 579.535 1181.675 579.550 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 906.805 16.405 906.975 18.275 ;
        RECT 931.185 16.405 931.355 17.935 ;
        RECT 955.565 16.065 955.735 17.935 ;
        RECT 1003.865 16.065 1004.035 17.935 ;
        RECT 1043.885 16.405 1044.055 17.935 ;
        RECT 1100.465 16.405 1100.635 17.935 ;
        RECT 1159.345 17.425 1159.515 18.275 ;
      LAYER mcon ;
        RECT 906.805 18.105 906.975 18.275 ;
        RECT 1159.345 18.105 1159.515 18.275 ;
        RECT 931.185 17.765 931.355 17.935 ;
        RECT 955.565 17.765 955.735 17.935 ;
        RECT 1003.865 17.765 1004.035 17.935 ;
        RECT 1043.885 17.765 1044.055 17.935 ;
        RECT 1100.465 17.765 1100.635 17.935 ;
      LAYER met1 ;
        RECT 1193.770 18.600 1194.090 18.660 ;
        RECT 1179.600 18.460 1194.090 18.600 ;
        RECT 864.870 18.260 865.190 18.320 ;
        RECT 906.745 18.260 907.035 18.305 ;
        RECT 864.870 18.120 907.035 18.260 ;
        RECT 864.870 18.060 865.190 18.120 ;
        RECT 906.745 18.075 907.035 18.120 ;
        RECT 1159.285 18.260 1159.575 18.305 ;
        RECT 1179.600 18.260 1179.740 18.460 ;
        RECT 1193.770 18.400 1194.090 18.460 ;
        RECT 1159.285 18.120 1179.740 18.260 ;
        RECT 1159.285 18.075 1159.575 18.120 ;
        RECT 931.125 17.920 931.415 17.965 ;
        RECT 955.505 17.920 955.795 17.965 ;
        RECT 931.125 17.780 955.795 17.920 ;
        RECT 931.125 17.735 931.415 17.780 ;
        RECT 955.505 17.735 955.795 17.780 ;
        RECT 1003.805 17.920 1004.095 17.965 ;
        RECT 1043.825 17.920 1044.115 17.965 ;
        RECT 1003.805 17.780 1044.115 17.920 ;
        RECT 1003.805 17.735 1004.095 17.780 ;
        RECT 1043.825 17.735 1044.115 17.780 ;
        RECT 1100.405 17.920 1100.695 17.965 ;
        RECT 1100.405 17.780 1132.360 17.920 ;
        RECT 1100.405 17.735 1100.695 17.780 ;
        RECT 1132.220 17.580 1132.360 17.780 ;
        RECT 1159.285 17.580 1159.575 17.625 ;
        RECT 1132.220 17.440 1159.575 17.580 ;
        RECT 1159.285 17.395 1159.575 17.440 ;
        RECT 906.745 16.560 907.035 16.605 ;
        RECT 931.125 16.560 931.415 16.605 ;
        RECT 906.745 16.420 931.415 16.560 ;
        RECT 906.745 16.375 907.035 16.420 ;
        RECT 931.125 16.375 931.415 16.420 ;
        RECT 1043.825 16.560 1044.115 16.605 ;
        RECT 1100.405 16.560 1100.695 16.605 ;
        RECT 1043.825 16.420 1100.695 16.560 ;
        RECT 1043.825 16.375 1044.115 16.420 ;
        RECT 1100.405 16.375 1100.695 16.420 ;
        RECT 955.505 16.220 955.795 16.265 ;
        RECT 1003.805 16.220 1004.095 16.265 ;
        RECT 955.505 16.080 1004.095 16.220 ;
        RECT 955.505 16.035 955.795 16.080 ;
        RECT 1003.805 16.035 1004.095 16.080 ;
      LAYER via ;
        RECT 864.900 18.060 865.160 18.320 ;
        RECT 1193.800 18.400 1194.060 18.660 ;
      LAYER met2 ;
        RECT 1194.270 1220.330 1194.830 1228.680 ;
        RECT 1193.860 1220.190 1194.830 1220.330 ;
        RECT 1193.860 18.690 1194.000 1220.190 ;
        RECT 1194.270 1219.680 1194.830 1220.190 ;
        RECT 1193.800 18.370 1194.060 18.690 ;
        RECT 864.900 18.030 865.160 18.350 ;
        RECT 864.960 2.400 865.100 18.030 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 956.025 18.105 956.195 20.655 ;
        RECT 983.625 18.105 983.795 20.655 ;
        RECT 1046.645 18.105 1046.815 19.975 ;
        RECT 1082.525 18.105 1082.695 19.975 ;
        RECT 1126.225 16.745 1126.395 18.275 ;
        RECT 1159.805 16.745 1159.975 17.595 ;
        RECT 1178.665 17.255 1178.835 17.595 ;
        RECT 1179.585 17.425 1182.515 17.595 ;
        RECT 1197.525 17.425 1197.695 18.955 ;
        RECT 1179.585 17.255 1179.755 17.425 ;
        RECT 1178.665 17.085 1179.755 17.255 ;
      LAYER mcon ;
        RECT 956.025 20.485 956.195 20.655 ;
        RECT 983.625 20.485 983.795 20.655 ;
        RECT 1046.645 19.805 1046.815 19.975 ;
        RECT 1082.525 19.805 1082.695 19.975 ;
        RECT 1197.525 18.785 1197.695 18.955 ;
        RECT 1126.225 18.105 1126.395 18.275 ;
        RECT 1159.805 17.425 1159.975 17.595 ;
        RECT 1178.665 17.425 1178.835 17.595 ;
        RECT 1182.345 17.425 1182.515 17.595 ;
      LAYER met1 ;
        RECT 955.965 20.640 956.255 20.685 ;
        RECT 983.565 20.640 983.855 20.685 ;
        RECT 955.965 20.500 983.855 20.640 ;
        RECT 955.965 20.455 956.255 20.500 ;
        RECT 983.565 20.455 983.855 20.500 ;
        RECT 1046.585 19.960 1046.875 20.005 ;
        RECT 1082.465 19.960 1082.755 20.005 ;
        RECT 1046.585 19.820 1082.755 19.960 ;
        RECT 1046.585 19.775 1046.875 19.820 ;
        RECT 1082.465 19.775 1082.755 19.820 ;
        RECT 882.810 18.940 883.130 19.000 ;
        RECT 1197.465 18.940 1197.755 18.985 ;
        RECT 1201.130 18.940 1201.450 19.000 ;
        RECT 882.810 18.800 907.420 18.940 ;
        RECT 882.810 18.740 883.130 18.800 ;
        RECT 907.280 18.260 907.420 18.800 ;
        RECT 1197.465 18.800 1201.450 18.940 ;
        RECT 1197.465 18.755 1197.755 18.800 ;
        RECT 1201.130 18.740 1201.450 18.800 ;
        RECT 955.965 18.260 956.255 18.305 ;
        RECT 907.280 18.120 956.255 18.260 ;
        RECT 955.965 18.075 956.255 18.120 ;
        RECT 983.565 18.260 983.855 18.305 ;
        RECT 1046.585 18.260 1046.875 18.305 ;
        RECT 983.565 18.120 1046.875 18.260 ;
        RECT 983.565 18.075 983.855 18.120 ;
        RECT 1046.585 18.075 1046.875 18.120 ;
        RECT 1082.465 18.260 1082.755 18.305 ;
        RECT 1126.165 18.260 1126.455 18.305 ;
        RECT 1082.465 18.120 1126.455 18.260 ;
        RECT 1082.465 18.075 1082.755 18.120 ;
        RECT 1126.165 18.075 1126.455 18.120 ;
        RECT 1159.745 17.580 1160.035 17.625 ;
        RECT 1178.605 17.580 1178.895 17.625 ;
        RECT 1159.745 17.440 1178.895 17.580 ;
        RECT 1159.745 17.395 1160.035 17.440 ;
        RECT 1178.605 17.395 1178.895 17.440 ;
        RECT 1182.285 17.580 1182.575 17.625 ;
        RECT 1197.465 17.580 1197.755 17.625 ;
        RECT 1182.285 17.440 1197.755 17.580 ;
        RECT 1182.285 17.395 1182.575 17.440 ;
        RECT 1197.465 17.395 1197.755 17.440 ;
        RECT 1126.165 16.900 1126.455 16.945 ;
        RECT 1159.745 16.900 1160.035 16.945 ;
        RECT 1126.165 16.760 1160.035 16.900 ;
        RECT 1126.165 16.715 1126.455 16.760 ;
        RECT 1159.745 16.715 1160.035 16.760 ;
      LAYER via ;
        RECT 882.840 18.740 883.100 19.000 ;
        RECT 1201.160 18.740 1201.420 19.000 ;
      LAYER met2 ;
        RECT 1203.010 1220.330 1203.570 1228.680 ;
        RECT 1201.220 1220.190 1203.570 1220.330 ;
        RECT 1201.220 19.030 1201.360 1220.190 ;
        RECT 1203.010 1219.680 1203.570 1220.190 ;
        RECT 882.840 18.710 883.100 19.030 ;
        RECT 1201.160 18.710 1201.420 19.030 ;
        RECT 882.900 2.400 883.040 18.710 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1179.125 17.425 1179.295 18.615 ;
      LAYER mcon ;
        RECT 1179.125 18.445 1179.295 18.615 ;
      LAYER met1 ;
        RECT 1207.570 1196.700 1207.890 1196.760 ;
        RECT 1210.790 1196.700 1211.110 1196.760 ;
        RECT 1207.570 1196.560 1211.110 1196.700 ;
        RECT 1207.570 1196.500 1207.890 1196.560 ;
        RECT 1210.790 1196.500 1211.110 1196.560 ;
        RECT 900.750 19.280 901.070 19.340 ;
        RECT 900.750 19.140 907.880 19.280 ;
        RECT 900.750 19.080 901.070 19.140 ;
        RECT 907.740 18.600 907.880 19.140 ;
        RECT 1179.065 18.600 1179.355 18.645 ;
        RECT 907.740 18.460 1179.355 18.600 ;
        RECT 1179.065 18.415 1179.355 18.460 ;
        RECT 1207.570 17.920 1207.890 17.980 ;
        RECT 1181.900 17.780 1207.890 17.920 ;
        RECT 1179.065 17.580 1179.355 17.625 ;
        RECT 1181.900 17.580 1182.040 17.780 ;
        RECT 1207.570 17.720 1207.890 17.780 ;
        RECT 1179.065 17.440 1182.040 17.580 ;
        RECT 1179.065 17.395 1179.355 17.440 ;
      LAYER via ;
        RECT 1207.600 1196.500 1207.860 1196.760 ;
        RECT 1210.820 1196.500 1211.080 1196.760 ;
        RECT 900.780 19.080 901.040 19.340 ;
        RECT 1207.600 17.720 1207.860 17.980 ;
      LAYER met2 ;
        RECT 1212.210 1220.330 1212.770 1228.680 ;
        RECT 1210.880 1220.190 1212.770 1220.330 ;
        RECT 1210.880 1196.790 1211.020 1220.190 ;
        RECT 1212.210 1219.680 1212.770 1220.190 ;
        RECT 1207.600 1196.470 1207.860 1196.790 ;
        RECT 1210.820 1196.470 1211.080 1196.790 ;
        RECT 900.780 19.050 901.040 19.370 ;
        RECT 900.840 2.400 900.980 19.050 ;
        RECT 1207.660 18.010 1207.800 1196.470 ;
        RECT 1207.600 17.690 1207.860 18.010 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 955.105 16.745 955.275 18.955 ;
      LAYER mcon ;
        RECT 955.105 18.785 955.275 18.955 ;
      LAYER met1 ;
        RECT 955.045 18.940 955.335 18.985 ;
        RECT 955.045 18.800 1197.220 18.940 ;
        RECT 955.045 18.755 955.335 18.800 ;
        RECT 1197.080 18.600 1197.220 18.800 ;
        RECT 1222.290 18.600 1222.610 18.660 ;
        RECT 1197.080 18.460 1222.610 18.600 ;
        RECT 1222.290 18.400 1222.610 18.460 ;
        RECT 918.690 16.900 919.010 16.960 ;
        RECT 955.045 16.900 955.335 16.945 ;
        RECT 918.690 16.760 955.335 16.900 ;
        RECT 918.690 16.700 919.010 16.760 ;
        RECT 955.045 16.715 955.335 16.760 ;
      LAYER via ;
        RECT 1222.320 18.400 1222.580 18.660 ;
        RECT 918.720 16.700 918.980 16.960 ;
      LAYER met2 ;
        RECT 1221.410 1220.330 1221.970 1228.680 ;
        RECT 1221.410 1220.190 1222.520 1220.330 ;
        RECT 1221.410 1219.680 1221.970 1220.190 ;
        RECT 1222.380 18.690 1222.520 1220.190 ;
        RECT 1222.320 18.370 1222.580 18.690 ;
        RECT 918.720 16.670 918.980 16.990 ;
        RECT 918.780 2.400 918.920 16.670 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 936.170 27.440 936.490 27.500 ;
        RECT 1228.270 27.440 1228.590 27.500 ;
        RECT 936.170 27.300 1228.590 27.440 ;
        RECT 936.170 27.240 936.490 27.300 ;
        RECT 1228.270 27.240 1228.590 27.300 ;
      LAYER via ;
        RECT 936.200 27.240 936.460 27.500 ;
        RECT 1228.300 27.240 1228.560 27.500 ;
      LAYER met2 ;
        RECT 1230.610 1221.010 1231.170 1228.680 ;
        RECT 1228.820 1220.870 1231.170 1221.010 ;
        RECT 1228.820 1196.530 1228.960 1220.870 ;
        RECT 1230.610 1219.680 1231.170 1220.870 ;
        RECT 1228.360 1196.390 1228.960 1196.530 ;
        RECT 1228.360 27.530 1228.500 1196.390 ;
        RECT 936.200 27.210 936.460 27.530 ;
        RECT 1228.300 27.210 1228.560 27.530 ;
        RECT 936.260 2.400 936.400 27.210 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1235.245 386.325 1235.415 434.775 ;
        RECT 1237.085 186.065 1237.255 227.715 ;
        RECT 1237.085 138.125 1237.255 156.655 ;
      LAYER mcon ;
        RECT 1235.245 434.605 1235.415 434.775 ;
        RECT 1237.085 227.545 1237.255 227.715 ;
        RECT 1237.085 156.485 1237.255 156.655 ;
      LAYER met1 ;
        RECT 1236.090 1196.700 1236.410 1196.760 ;
        RECT 1238.850 1196.700 1239.170 1196.760 ;
        RECT 1236.090 1196.560 1239.170 1196.700 ;
        RECT 1236.090 1196.500 1236.410 1196.560 ;
        RECT 1238.850 1196.500 1239.170 1196.560 ;
        RECT 1236.090 1124.760 1236.410 1125.020 ;
        RECT 1236.180 1124.280 1236.320 1124.760 ;
        RECT 1236.550 1124.280 1236.870 1124.340 ;
        RECT 1236.180 1124.140 1236.870 1124.280 ;
        RECT 1236.550 1124.080 1236.870 1124.140 ;
        RECT 1236.550 1062.740 1236.870 1062.800 ;
        RECT 1237.010 1062.740 1237.330 1062.800 ;
        RECT 1236.550 1062.600 1237.330 1062.740 ;
        RECT 1236.550 1062.540 1236.870 1062.600 ;
        RECT 1237.010 1062.540 1237.330 1062.600 ;
        RECT 1235.170 966.180 1235.490 966.240 ;
        RECT 1236.550 966.180 1236.870 966.240 ;
        RECT 1235.170 966.040 1236.870 966.180 ;
        RECT 1235.170 965.980 1235.490 966.040 ;
        RECT 1236.550 965.980 1236.870 966.040 ;
        RECT 1235.170 869.620 1235.490 869.680 ;
        RECT 1236.550 869.620 1236.870 869.680 ;
        RECT 1235.170 869.480 1236.870 869.620 ;
        RECT 1235.170 869.420 1235.490 869.480 ;
        RECT 1236.550 869.420 1236.870 869.480 ;
        RECT 1235.170 821.000 1235.490 821.060 ;
        RECT 1236.090 821.000 1236.410 821.060 ;
        RECT 1235.170 820.860 1236.410 821.000 ;
        RECT 1235.170 820.800 1235.490 820.860 ;
        RECT 1236.090 820.800 1236.410 820.860 ;
        RECT 1236.090 689.900 1236.410 690.160 ;
        RECT 1236.180 689.760 1236.320 689.900 ;
        RECT 1236.550 689.760 1236.870 689.820 ;
        RECT 1236.180 689.620 1236.870 689.760 ;
        RECT 1236.550 689.560 1236.870 689.620 ;
        RECT 1236.090 593.340 1236.410 593.600 ;
        RECT 1236.180 593.200 1236.320 593.340 ;
        RECT 1236.550 593.200 1236.870 593.260 ;
        RECT 1236.180 593.060 1236.870 593.200 ;
        RECT 1236.550 593.000 1236.870 593.060 ;
        RECT 1236.090 496.780 1236.410 497.040 ;
        RECT 1236.180 496.640 1236.320 496.780 ;
        RECT 1236.550 496.640 1236.870 496.700 ;
        RECT 1236.180 496.500 1236.870 496.640 ;
        RECT 1236.550 496.440 1236.870 496.500 ;
        RECT 1235.185 434.760 1235.475 434.805 ;
        RECT 1235.630 434.760 1235.950 434.820 ;
        RECT 1235.185 434.620 1235.950 434.760 ;
        RECT 1235.185 434.575 1235.475 434.620 ;
        RECT 1235.630 434.560 1235.950 434.620 ;
        RECT 1235.170 386.480 1235.490 386.540 ;
        RECT 1234.975 386.340 1235.490 386.480 ;
        RECT 1235.170 386.280 1235.490 386.340 ;
        RECT 1235.630 283.120 1235.950 283.180 ;
        RECT 1236.550 283.120 1236.870 283.180 ;
        RECT 1235.630 282.980 1236.870 283.120 ;
        RECT 1235.630 282.920 1235.950 282.980 ;
        RECT 1236.550 282.920 1236.870 282.980 ;
        RECT 1235.630 234.500 1235.950 234.560 ;
        RECT 1237.010 234.500 1237.330 234.560 ;
        RECT 1235.630 234.360 1237.330 234.500 ;
        RECT 1235.630 234.300 1235.950 234.360 ;
        RECT 1237.010 234.300 1237.330 234.360 ;
        RECT 1237.010 227.700 1237.330 227.760 ;
        RECT 1236.815 227.560 1237.330 227.700 ;
        RECT 1237.010 227.500 1237.330 227.560 ;
        RECT 1237.010 186.220 1237.330 186.280 ;
        RECT 1236.815 186.080 1237.330 186.220 ;
        RECT 1237.010 186.020 1237.330 186.080 ;
        RECT 1237.010 156.640 1237.330 156.700 ;
        RECT 1236.815 156.500 1237.330 156.640 ;
        RECT 1237.010 156.440 1237.330 156.500 ;
        RECT 1237.010 138.280 1237.330 138.340 ;
        RECT 1236.815 138.140 1237.330 138.280 ;
        RECT 1237.010 138.080 1237.330 138.140 ;
        RECT 954.110 22.680 954.430 22.740 ;
        RECT 1236.550 22.680 1236.870 22.740 ;
        RECT 954.110 22.540 1236.870 22.680 ;
        RECT 954.110 22.480 954.430 22.540 ;
        RECT 1236.550 22.480 1236.870 22.540 ;
      LAYER via ;
        RECT 1236.120 1196.500 1236.380 1196.760 ;
        RECT 1238.880 1196.500 1239.140 1196.760 ;
        RECT 1236.120 1124.760 1236.380 1125.020 ;
        RECT 1236.580 1124.080 1236.840 1124.340 ;
        RECT 1236.580 1062.540 1236.840 1062.800 ;
        RECT 1237.040 1062.540 1237.300 1062.800 ;
        RECT 1235.200 965.980 1235.460 966.240 ;
        RECT 1236.580 965.980 1236.840 966.240 ;
        RECT 1235.200 869.420 1235.460 869.680 ;
        RECT 1236.580 869.420 1236.840 869.680 ;
        RECT 1235.200 820.800 1235.460 821.060 ;
        RECT 1236.120 820.800 1236.380 821.060 ;
        RECT 1236.120 689.900 1236.380 690.160 ;
        RECT 1236.580 689.560 1236.840 689.820 ;
        RECT 1236.120 593.340 1236.380 593.600 ;
        RECT 1236.580 593.000 1236.840 593.260 ;
        RECT 1236.120 496.780 1236.380 497.040 ;
        RECT 1236.580 496.440 1236.840 496.700 ;
        RECT 1235.660 434.560 1235.920 434.820 ;
        RECT 1235.200 386.280 1235.460 386.540 ;
        RECT 1235.660 282.920 1235.920 283.180 ;
        RECT 1236.580 282.920 1236.840 283.180 ;
        RECT 1235.660 234.300 1235.920 234.560 ;
        RECT 1237.040 234.300 1237.300 234.560 ;
        RECT 1237.040 227.500 1237.300 227.760 ;
        RECT 1237.040 186.020 1237.300 186.280 ;
        RECT 1237.040 156.440 1237.300 156.700 ;
        RECT 1237.040 138.080 1237.300 138.340 ;
        RECT 954.140 22.480 954.400 22.740 ;
        RECT 1236.580 22.480 1236.840 22.740 ;
      LAYER met2 ;
        RECT 1239.810 1220.330 1240.370 1228.680 ;
        RECT 1238.940 1220.190 1240.370 1220.330 ;
        RECT 1238.940 1196.790 1239.080 1220.190 ;
        RECT 1239.810 1219.680 1240.370 1220.190 ;
        RECT 1236.120 1196.470 1236.380 1196.790 ;
        RECT 1238.880 1196.470 1239.140 1196.790 ;
        RECT 1236.180 1125.050 1236.320 1196.470 ;
        RECT 1236.120 1124.730 1236.380 1125.050 ;
        RECT 1236.580 1124.050 1236.840 1124.370 ;
        RECT 1236.640 1110.850 1236.780 1124.050 ;
        RECT 1236.640 1110.710 1237.240 1110.850 ;
        RECT 1237.100 1062.830 1237.240 1110.710 ;
        RECT 1236.580 1062.510 1236.840 1062.830 ;
        RECT 1237.040 1062.510 1237.300 1062.830 ;
        RECT 1236.640 1027.890 1236.780 1062.510 ;
        RECT 1236.180 1027.750 1236.780 1027.890 ;
        RECT 1236.180 1014.405 1236.320 1027.750 ;
        RECT 1235.190 1014.035 1235.470 1014.405 ;
        RECT 1236.110 1014.035 1236.390 1014.405 ;
        RECT 1235.260 966.270 1235.400 1014.035 ;
        RECT 1235.200 965.950 1235.460 966.270 ;
        RECT 1236.580 965.950 1236.840 966.270 ;
        RECT 1236.640 931.330 1236.780 965.950 ;
        RECT 1236.180 931.190 1236.780 931.330 ;
        RECT 1236.180 917.845 1236.320 931.190 ;
        RECT 1235.190 917.475 1235.470 917.845 ;
        RECT 1236.110 917.475 1236.390 917.845 ;
        RECT 1235.260 869.710 1235.400 917.475 ;
        RECT 1235.200 869.390 1235.460 869.710 ;
        RECT 1236.580 869.390 1236.840 869.710 ;
        RECT 1236.640 834.770 1236.780 869.390 ;
        RECT 1236.180 834.630 1236.780 834.770 ;
        RECT 1236.180 821.090 1236.320 834.630 ;
        RECT 1235.200 820.770 1235.460 821.090 ;
        RECT 1236.120 820.770 1236.380 821.090 ;
        RECT 1235.260 773.005 1235.400 820.770 ;
        RECT 1235.190 772.635 1235.470 773.005 ;
        RECT 1236.570 772.635 1236.850 773.005 ;
        RECT 1236.640 738.210 1236.780 772.635 ;
        RECT 1236.180 738.070 1236.780 738.210 ;
        RECT 1236.180 690.190 1236.320 738.070 ;
        RECT 1236.120 689.870 1236.380 690.190 ;
        RECT 1236.580 689.530 1236.840 689.850 ;
        RECT 1236.640 641.650 1236.780 689.530 ;
        RECT 1236.180 641.510 1236.780 641.650 ;
        RECT 1236.180 593.630 1236.320 641.510 ;
        RECT 1236.120 593.310 1236.380 593.630 ;
        RECT 1236.580 592.970 1236.840 593.290 ;
        RECT 1236.640 545.090 1236.780 592.970 ;
        RECT 1236.180 544.950 1236.780 545.090 ;
        RECT 1236.180 497.070 1236.320 544.950 ;
        RECT 1236.120 496.750 1236.380 497.070 ;
        RECT 1236.580 496.410 1236.840 496.730 ;
        RECT 1236.640 448.530 1236.780 496.410 ;
        RECT 1235.720 448.390 1236.780 448.530 ;
        RECT 1235.720 434.850 1235.860 448.390 ;
        RECT 1235.660 434.530 1235.920 434.850 ;
        RECT 1235.200 386.250 1235.460 386.570 ;
        RECT 1235.260 351.290 1235.400 386.250 ;
        RECT 1235.260 351.150 1235.860 351.290 ;
        RECT 1235.720 283.210 1235.860 351.150 ;
        RECT 1235.660 282.890 1235.920 283.210 ;
        RECT 1236.580 282.890 1236.840 283.210 ;
        RECT 1236.640 235.010 1236.780 282.890 ;
        RECT 1235.720 234.870 1236.780 235.010 ;
        RECT 1235.720 234.590 1235.860 234.870 ;
        RECT 1235.660 234.270 1235.920 234.590 ;
        RECT 1237.040 234.270 1237.300 234.590 ;
        RECT 1237.100 227.790 1237.240 234.270 ;
        RECT 1237.040 227.470 1237.300 227.790 ;
        RECT 1237.040 185.990 1237.300 186.310 ;
        RECT 1237.100 156.730 1237.240 185.990 ;
        RECT 1237.040 156.410 1237.300 156.730 ;
        RECT 1237.040 138.050 1237.300 138.370 ;
        RECT 1237.100 110.570 1237.240 138.050 ;
        RECT 1236.640 110.430 1237.240 110.570 ;
        RECT 1236.640 22.770 1236.780 110.430 ;
        RECT 954.140 22.450 954.400 22.770 ;
        RECT 1236.580 22.450 1236.840 22.770 ;
        RECT 954.200 2.400 954.340 22.450 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER via2 ;
        RECT 1235.190 1014.080 1235.470 1014.360 ;
        RECT 1236.110 1014.080 1236.390 1014.360 ;
        RECT 1235.190 917.520 1235.470 917.800 ;
        RECT 1236.110 917.520 1236.390 917.800 ;
        RECT 1235.190 772.680 1235.470 772.960 ;
        RECT 1236.570 772.680 1236.850 772.960 ;
      LAYER met3 ;
        RECT 1235.165 1014.370 1235.495 1014.385 ;
        RECT 1236.085 1014.370 1236.415 1014.385 ;
        RECT 1235.165 1014.070 1236.415 1014.370 ;
        RECT 1235.165 1014.055 1235.495 1014.070 ;
        RECT 1236.085 1014.055 1236.415 1014.070 ;
        RECT 1235.165 917.810 1235.495 917.825 ;
        RECT 1236.085 917.810 1236.415 917.825 ;
        RECT 1235.165 917.510 1236.415 917.810 ;
        RECT 1235.165 917.495 1235.495 917.510 ;
        RECT 1236.085 917.495 1236.415 917.510 ;
        RECT 1235.165 772.970 1235.495 772.985 ;
        RECT 1236.545 772.970 1236.875 772.985 ;
        RECT 1235.165 772.670 1236.875 772.970 ;
        RECT 1235.165 772.655 1235.495 772.670 ;
        RECT 1236.545 772.655 1236.875 772.670 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 23.360 972.370 23.420 ;
        RECT 1249.890 23.360 1250.210 23.420 ;
        RECT 972.050 23.220 1250.210 23.360 ;
        RECT 972.050 23.160 972.370 23.220 ;
        RECT 1249.890 23.160 1250.210 23.220 ;
      LAYER via ;
        RECT 972.080 23.160 972.340 23.420 ;
        RECT 1249.920 23.160 1250.180 23.420 ;
      LAYER met2 ;
        RECT 1249.010 1220.330 1249.570 1228.680 ;
        RECT 1249.010 1220.190 1250.120 1220.330 ;
        RECT 1249.010 1219.680 1249.570 1220.190 ;
        RECT 1249.980 23.450 1250.120 1220.190 ;
        RECT 972.080 23.130 972.340 23.450 ;
        RECT 1249.920 23.130 1250.180 23.450 ;
        RECT 972.140 2.400 972.280 23.130 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 36.620 651.290 36.680 ;
        RECT 1083.370 36.620 1083.690 36.680 ;
        RECT 650.970 36.480 1083.690 36.620 ;
        RECT 650.970 36.420 651.290 36.480 ;
        RECT 1083.370 36.420 1083.690 36.480 ;
      LAYER via ;
        RECT 651.000 36.420 651.260 36.680 ;
        RECT 1083.400 36.420 1083.660 36.680 ;
      LAYER met2 ;
        RECT 1083.870 1220.330 1084.430 1228.680 ;
        RECT 1083.460 1220.190 1084.430 1220.330 ;
        RECT 1083.460 36.710 1083.600 1220.190 ;
        RECT 1083.870 1219.680 1084.430 1220.190 ;
        RECT 651.000 36.390 651.260 36.710 ;
        RECT 1083.400 36.390 1083.660 36.710 ;
        RECT 651.060 2.400 651.200 36.390 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 990.450 22.000 990.770 22.060 ;
        RECT 1256.330 22.000 1256.650 22.060 ;
        RECT 990.450 21.860 1256.650 22.000 ;
        RECT 990.450 21.800 990.770 21.860 ;
        RECT 1256.330 21.800 1256.650 21.860 ;
      LAYER via ;
        RECT 990.480 21.800 990.740 22.060 ;
        RECT 1256.360 21.800 1256.620 22.060 ;
      LAYER met2 ;
        RECT 1258.210 1220.330 1258.770 1228.680 ;
        RECT 1256.420 1220.190 1258.770 1220.330 ;
        RECT 1256.420 22.090 1256.560 1220.190 ;
        RECT 1258.210 1219.680 1258.770 1220.190 ;
        RECT 990.480 21.770 990.740 22.090 ;
        RECT 1256.360 21.770 1256.620 22.090 ;
        RECT 990.540 11.290 990.680 21.770 ;
        RECT 990.080 11.150 990.680 11.290 ;
        RECT 990.080 2.400 990.220 11.150 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1263.765 786.505 1263.935 821.015 ;
        RECT 1263.765 689.605 1263.935 724.455 ;
        RECT 1263.765 593.045 1263.935 627.895 ;
        RECT 1263.765 496.485 1263.935 531.335 ;
        RECT 1263.765 386.325 1263.935 434.775 ;
        RECT 1263.765 331.245 1263.935 338.555 ;
        RECT 1263.765 89.845 1263.935 137.955 ;
      LAYER mcon ;
        RECT 1263.765 820.845 1263.935 821.015 ;
        RECT 1263.765 724.285 1263.935 724.455 ;
        RECT 1263.765 627.725 1263.935 627.895 ;
        RECT 1263.765 531.165 1263.935 531.335 ;
        RECT 1263.765 434.605 1263.935 434.775 ;
        RECT 1263.765 338.385 1263.935 338.555 ;
        RECT 1263.765 137.785 1263.935 137.955 ;
      LAYER met1 ;
        RECT 1263.230 1124.960 1263.550 1125.020 ;
        RECT 1264.150 1124.960 1264.470 1125.020 ;
        RECT 1263.230 1124.820 1264.470 1124.960 ;
        RECT 1263.230 1124.760 1263.550 1124.820 ;
        RECT 1264.150 1124.760 1264.470 1124.820 ;
        RECT 1263.230 1028.400 1263.550 1028.460 ;
        RECT 1264.150 1028.400 1264.470 1028.460 ;
        RECT 1263.230 1028.260 1264.470 1028.400 ;
        RECT 1263.230 1028.200 1263.550 1028.260 ;
        RECT 1264.150 1028.200 1264.470 1028.260 ;
        RECT 1263.230 931.840 1263.550 931.900 ;
        RECT 1264.150 931.840 1264.470 931.900 ;
        RECT 1263.230 931.700 1264.470 931.840 ;
        RECT 1263.230 931.640 1263.550 931.700 ;
        RECT 1264.150 931.640 1264.470 931.700 ;
        RECT 1262.770 869.620 1263.090 869.680 ;
        RECT 1264.150 869.620 1264.470 869.680 ;
        RECT 1262.770 869.480 1264.470 869.620 ;
        RECT 1262.770 869.420 1263.090 869.480 ;
        RECT 1264.150 869.420 1264.470 869.480 ;
        RECT 1263.230 835.280 1263.550 835.340 ;
        RECT 1264.150 835.280 1264.470 835.340 ;
        RECT 1263.230 835.140 1264.470 835.280 ;
        RECT 1263.230 835.080 1263.550 835.140 ;
        RECT 1264.150 835.080 1264.470 835.140 ;
        RECT 1263.690 821.000 1264.010 821.060 ;
        RECT 1263.495 820.860 1264.010 821.000 ;
        RECT 1263.690 820.800 1264.010 820.860 ;
        RECT 1263.690 786.660 1264.010 786.720 ;
        RECT 1263.495 786.520 1264.010 786.660 ;
        RECT 1263.690 786.460 1264.010 786.520 ;
        RECT 1263.230 738.380 1263.550 738.440 ;
        RECT 1264.150 738.380 1264.470 738.440 ;
        RECT 1263.230 738.240 1264.470 738.380 ;
        RECT 1263.230 738.180 1263.550 738.240 ;
        RECT 1264.150 738.180 1264.470 738.240 ;
        RECT 1263.690 724.440 1264.010 724.500 ;
        RECT 1263.495 724.300 1264.010 724.440 ;
        RECT 1263.690 724.240 1264.010 724.300 ;
        RECT 1263.690 689.760 1264.010 689.820 ;
        RECT 1263.495 689.620 1264.010 689.760 ;
        RECT 1263.690 689.560 1264.010 689.620 ;
        RECT 1263.230 641.820 1263.550 641.880 ;
        RECT 1264.150 641.820 1264.470 641.880 ;
        RECT 1263.230 641.680 1264.470 641.820 ;
        RECT 1263.230 641.620 1263.550 641.680 ;
        RECT 1264.150 641.620 1264.470 641.680 ;
        RECT 1263.690 627.880 1264.010 627.940 ;
        RECT 1263.495 627.740 1264.010 627.880 ;
        RECT 1263.690 627.680 1264.010 627.740 ;
        RECT 1263.690 593.200 1264.010 593.260 ;
        RECT 1263.495 593.060 1264.010 593.200 ;
        RECT 1263.690 593.000 1264.010 593.060 ;
        RECT 1263.230 545.260 1263.550 545.320 ;
        RECT 1264.150 545.260 1264.470 545.320 ;
        RECT 1263.230 545.120 1264.470 545.260 ;
        RECT 1263.230 545.060 1263.550 545.120 ;
        RECT 1264.150 545.060 1264.470 545.120 ;
        RECT 1263.690 531.320 1264.010 531.380 ;
        RECT 1263.495 531.180 1264.010 531.320 ;
        RECT 1263.690 531.120 1264.010 531.180 ;
        RECT 1263.690 496.640 1264.010 496.700 ;
        RECT 1263.495 496.500 1264.010 496.640 ;
        RECT 1263.690 496.440 1264.010 496.500 ;
        RECT 1263.230 448.700 1263.550 448.760 ;
        RECT 1264.150 448.700 1264.470 448.760 ;
        RECT 1263.230 448.560 1264.470 448.700 ;
        RECT 1263.230 448.500 1263.550 448.560 ;
        RECT 1264.150 448.500 1264.470 448.560 ;
        RECT 1263.690 434.760 1264.010 434.820 ;
        RECT 1263.495 434.620 1264.010 434.760 ;
        RECT 1263.690 434.560 1264.010 434.620 ;
        RECT 1263.705 386.480 1263.995 386.525 ;
        RECT 1264.150 386.480 1264.470 386.540 ;
        RECT 1263.705 386.340 1264.470 386.480 ;
        RECT 1263.705 386.295 1263.995 386.340 ;
        RECT 1264.150 386.280 1264.470 386.340 ;
        RECT 1263.705 338.540 1263.995 338.585 ;
        RECT 1264.150 338.540 1264.470 338.600 ;
        RECT 1263.705 338.400 1264.470 338.540 ;
        RECT 1263.705 338.355 1263.995 338.400 ;
        RECT 1264.150 338.340 1264.470 338.400 ;
        RECT 1263.690 331.400 1264.010 331.460 ;
        RECT 1263.495 331.260 1264.010 331.400 ;
        RECT 1263.690 331.200 1264.010 331.260 ;
        RECT 1261.850 285.160 1262.170 285.220 ;
        RECT 1264.150 285.160 1264.470 285.220 ;
        RECT 1261.850 285.020 1264.470 285.160 ;
        RECT 1261.850 284.960 1262.170 285.020 ;
        RECT 1264.150 284.960 1264.470 285.020 ;
        RECT 1261.850 255.240 1262.170 255.300 ;
        RECT 1263.690 255.240 1264.010 255.300 ;
        RECT 1261.850 255.100 1264.010 255.240 ;
        RECT 1261.850 255.040 1262.170 255.100 ;
        RECT 1263.690 255.040 1264.010 255.100 ;
        RECT 1263.230 193.360 1263.550 193.420 ;
        RECT 1264.150 193.360 1264.470 193.420 ;
        RECT 1263.230 193.220 1264.470 193.360 ;
        RECT 1263.230 193.160 1263.550 193.220 ;
        RECT 1264.150 193.160 1264.470 193.220 ;
        RECT 1263.690 137.940 1264.010 138.000 ;
        RECT 1263.495 137.800 1264.010 137.940 ;
        RECT 1263.690 137.740 1264.010 137.800 ;
        RECT 1263.705 90.000 1263.995 90.045 ;
        RECT 1264.150 90.000 1264.470 90.060 ;
        RECT 1263.705 89.860 1264.470 90.000 ;
        RECT 1263.705 89.815 1263.995 89.860 ;
        RECT 1264.150 89.800 1264.470 89.860 ;
        RECT 1007.470 21.660 1007.790 21.720 ;
        RECT 1264.150 21.660 1264.470 21.720 ;
        RECT 1007.470 21.520 1264.470 21.660 ;
        RECT 1007.470 21.460 1007.790 21.520 ;
        RECT 1264.150 21.460 1264.470 21.520 ;
      LAYER via ;
        RECT 1263.260 1124.760 1263.520 1125.020 ;
        RECT 1264.180 1124.760 1264.440 1125.020 ;
        RECT 1263.260 1028.200 1263.520 1028.460 ;
        RECT 1264.180 1028.200 1264.440 1028.460 ;
        RECT 1263.260 931.640 1263.520 931.900 ;
        RECT 1264.180 931.640 1264.440 931.900 ;
        RECT 1262.800 869.420 1263.060 869.680 ;
        RECT 1264.180 869.420 1264.440 869.680 ;
        RECT 1263.260 835.080 1263.520 835.340 ;
        RECT 1264.180 835.080 1264.440 835.340 ;
        RECT 1263.720 820.800 1263.980 821.060 ;
        RECT 1263.720 786.460 1263.980 786.720 ;
        RECT 1263.260 738.180 1263.520 738.440 ;
        RECT 1264.180 738.180 1264.440 738.440 ;
        RECT 1263.720 724.240 1263.980 724.500 ;
        RECT 1263.720 689.560 1263.980 689.820 ;
        RECT 1263.260 641.620 1263.520 641.880 ;
        RECT 1264.180 641.620 1264.440 641.880 ;
        RECT 1263.720 627.680 1263.980 627.940 ;
        RECT 1263.720 593.000 1263.980 593.260 ;
        RECT 1263.260 545.060 1263.520 545.320 ;
        RECT 1264.180 545.060 1264.440 545.320 ;
        RECT 1263.720 531.120 1263.980 531.380 ;
        RECT 1263.720 496.440 1263.980 496.700 ;
        RECT 1263.260 448.500 1263.520 448.760 ;
        RECT 1264.180 448.500 1264.440 448.760 ;
        RECT 1263.720 434.560 1263.980 434.820 ;
        RECT 1264.180 386.280 1264.440 386.540 ;
        RECT 1264.180 338.340 1264.440 338.600 ;
        RECT 1263.720 331.200 1263.980 331.460 ;
        RECT 1261.880 284.960 1262.140 285.220 ;
        RECT 1264.180 284.960 1264.440 285.220 ;
        RECT 1261.880 255.040 1262.140 255.300 ;
        RECT 1263.720 255.040 1263.980 255.300 ;
        RECT 1263.260 193.160 1263.520 193.420 ;
        RECT 1264.180 193.160 1264.440 193.420 ;
        RECT 1263.720 137.740 1263.980 138.000 ;
        RECT 1264.180 89.800 1264.440 90.060 ;
        RECT 1007.500 21.460 1007.760 21.720 ;
        RECT 1264.180 21.460 1264.440 21.720 ;
      LAYER met2 ;
        RECT 1267.410 1220.330 1267.970 1228.680 ;
        RECT 1265.620 1220.190 1267.970 1220.330 ;
        RECT 1265.620 1196.530 1265.760 1220.190 ;
        RECT 1267.410 1219.680 1267.970 1220.190 ;
        RECT 1264.240 1196.390 1265.760 1196.530 ;
        RECT 1264.240 1125.050 1264.380 1196.390 ;
        RECT 1263.260 1124.730 1263.520 1125.050 ;
        RECT 1264.180 1124.730 1264.440 1125.050 ;
        RECT 1263.320 1124.450 1263.460 1124.730 ;
        RECT 1263.320 1124.310 1263.920 1124.450 ;
        RECT 1263.780 1076.850 1263.920 1124.310 ;
        RECT 1263.780 1076.710 1264.380 1076.850 ;
        RECT 1264.240 1028.490 1264.380 1076.710 ;
        RECT 1263.260 1028.170 1263.520 1028.490 ;
        RECT 1264.180 1028.170 1264.440 1028.490 ;
        RECT 1263.320 1027.890 1263.460 1028.170 ;
        RECT 1263.320 1027.750 1263.920 1027.890 ;
        RECT 1263.780 980.290 1263.920 1027.750 ;
        RECT 1263.780 980.150 1264.380 980.290 ;
        RECT 1264.240 931.930 1264.380 980.150 ;
        RECT 1263.260 931.610 1263.520 931.930 ;
        RECT 1264.180 931.610 1264.440 931.930 ;
        RECT 1263.320 931.330 1263.460 931.610 ;
        RECT 1263.320 931.190 1263.920 931.330 ;
        RECT 1263.780 917.845 1263.920 931.190 ;
        RECT 1262.790 917.475 1263.070 917.845 ;
        RECT 1263.710 917.475 1263.990 917.845 ;
        RECT 1262.860 869.710 1263.000 917.475 ;
        RECT 1262.800 869.390 1263.060 869.710 ;
        RECT 1264.180 869.390 1264.440 869.710 ;
        RECT 1264.240 835.370 1264.380 869.390 ;
        RECT 1263.260 835.050 1263.520 835.370 ;
        RECT 1264.180 835.050 1264.440 835.370 ;
        RECT 1263.320 834.770 1263.460 835.050 ;
        RECT 1263.320 834.630 1263.920 834.770 ;
        RECT 1263.780 821.090 1263.920 834.630 ;
        RECT 1263.720 820.770 1263.980 821.090 ;
        RECT 1263.720 786.430 1263.980 786.750 ;
        RECT 1263.780 772.890 1263.920 786.430 ;
        RECT 1263.780 772.750 1264.380 772.890 ;
        RECT 1264.240 738.470 1264.380 772.750 ;
        RECT 1263.260 738.210 1263.520 738.470 ;
        RECT 1263.260 738.150 1263.920 738.210 ;
        RECT 1264.180 738.150 1264.440 738.470 ;
        RECT 1263.320 738.070 1263.920 738.150 ;
        RECT 1263.780 724.530 1263.920 738.070 ;
        RECT 1263.720 724.210 1263.980 724.530 ;
        RECT 1263.720 689.530 1263.980 689.850 ;
        RECT 1263.780 676.330 1263.920 689.530 ;
        RECT 1263.780 676.190 1264.380 676.330 ;
        RECT 1264.240 641.910 1264.380 676.190 ;
        RECT 1263.260 641.650 1263.520 641.910 ;
        RECT 1263.260 641.590 1263.920 641.650 ;
        RECT 1264.180 641.590 1264.440 641.910 ;
        RECT 1263.320 641.510 1263.920 641.590 ;
        RECT 1263.780 627.970 1263.920 641.510 ;
        RECT 1263.720 627.650 1263.980 627.970 ;
        RECT 1263.720 592.970 1263.980 593.290 ;
        RECT 1263.780 579.770 1263.920 592.970 ;
        RECT 1263.780 579.630 1264.380 579.770 ;
        RECT 1264.240 545.350 1264.380 579.630 ;
        RECT 1263.260 545.090 1263.520 545.350 ;
        RECT 1263.260 545.030 1263.920 545.090 ;
        RECT 1264.180 545.030 1264.440 545.350 ;
        RECT 1263.320 544.950 1263.920 545.030 ;
        RECT 1263.780 531.410 1263.920 544.950 ;
        RECT 1263.720 531.090 1263.980 531.410 ;
        RECT 1263.720 496.410 1263.980 496.730 ;
        RECT 1263.780 483.210 1263.920 496.410 ;
        RECT 1263.780 483.070 1264.380 483.210 ;
        RECT 1264.240 448.790 1264.380 483.070 ;
        RECT 1263.260 448.530 1263.520 448.790 ;
        RECT 1263.260 448.470 1263.920 448.530 ;
        RECT 1264.180 448.470 1264.440 448.790 ;
        RECT 1263.320 448.390 1263.920 448.470 ;
        RECT 1263.780 434.850 1263.920 448.390 ;
        RECT 1263.720 434.530 1263.980 434.850 ;
        RECT 1264.180 386.250 1264.440 386.570 ;
        RECT 1264.240 338.630 1264.380 386.250 ;
        RECT 1264.180 338.310 1264.440 338.630 ;
        RECT 1263.720 331.170 1263.980 331.490 ;
        RECT 1263.780 304.370 1263.920 331.170 ;
        RECT 1263.780 304.230 1264.380 304.370 ;
        RECT 1264.240 285.250 1264.380 304.230 ;
        RECT 1261.880 284.930 1262.140 285.250 ;
        RECT 1264.180 284.930 1264.440 285.250 ;
        RECT 1261.940 255.330 1262.080 284.930 ;
        RECT 1261.880 255.010 1262.140 255.330 ;
        RECT 1263.720 255.010 1263.980 255.330 ;
        RECT 1263.780 217.330 1263.920 255.010 ;
        RECT 1263.320 217.190 1263.920 217.330 ;
        RECT 1263.320 193.450 1263.460 217.190 ;
        RECT 1263.260 193.130 1263.520 193.450 ;
        RECT 1264.180 193.130 1264.440 193.450 ;
        RECT 1264.240 159.530 1264.380 193.130 ;
        RECT 1264.240 159.390 1264.840 159.530 ;
        RECT 1264.700 158.170 1264.840 159.390 ;
        RECT 1263.780 158.030 1264.840 158.170 ;
        RECT 1263.780 138.030 1263.920 158.030 ;
        RECT 1263.720 137.710 1263.980 138.030 ;
        RECT 1264.180 89.770 1264.440 90.090 ;
        RECT 1264.240 21.750 1264.380 89.770 ;
        RECT 1007.500 21.430 1007.760 21.750 ;
        RECT 1264.180 21.430 1264.440 21.750 ;
        RECT 1007.560 2.400 1007.700 21.430 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 1262.790 917.520 1263.070 917.800 ;
        RECT 1263.710 917.520 1263.990 917.800 ;
      LAYER met3 ;
        RECT 1262.765 917.810 1263.095 917.825 ;
        RECT 1263.685 917.810 1264.015 917.825 ;
        RECT 1262.765 917.510 1264.015 917.810 ;
        RECT 1262.765 917.495 1263.095 917.510 ;
        RECT 1263.685 917.495 1264.015 917.510 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1025.410 21.320 1025.730 21.380 ;
        RECT 1277.030 21.320 1277.350 21.380 ;
        RECT 1025.410 21.180 1277.350 21.320 ;
        RECT 1025.410 21.120 1025.730 21.180 ;
        RECT 1277.030 21.120 1277.350 21.180 ;
      LAYER via ;
        RECT 1025.440 21.120 1025.700 21.380 ;
        RECT 1277.060 21.120 1277.320 21.380 ;
      LAYER met2 ;
        RECT 1276.610 1220.330 1277.170 1228.680 ;
        RECT 1276.610 1219.680 1277.260 1220.330 ;
        RECT 1277.120 21.410 1277.260 1219.680 ;
        RECT 1025.440 21.090 1025.700 21.410 ;
        RECT 1277.060 21.090 1277.320 21.410 ;
        RECT 1025.500 2.400 1025.640 21.090 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 19.280 1043.670 19.340 ;
        RECT 1283.930 19.280 1284.250 19.340 ;
        RECT 1043.350 19.140 1284.250 19.280 ;
        RECT 1043.350 19.080 1043.670 19.140 ;
        RECT 1283.930 19.080 1284.250 19.140 ;
      LAYER via ;
        RECT 1043.380 19.080 1043.640 19.340 ;
        RECT 1283.960 19.080 1284.220 19.340 ;
      LAYER met2 ;
        RECT 1285.810 1220.330 1286.370 1228.680 ;
        RECT 1284.020 1220.190 1286.370 1220.330 ;
        RECT 1284.020 19.370 1284.160 1220.190 ;
        RECT 1285.810 1219.680 1286.370 1220.190 ;
        RECT 1043.380 19.050 1043.640 19.370 ;
        RECT 1283.960 19.050 1284.220 19.370 ;
        RECT 1043.440 2.400 1043.580 19.050 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1290.445 386.325 1290.615 434.775 ;
        RECT 1290.905 241.485 1291.075 289.595 ;
      LAYER mcon ;
        RECT 1290.445 434.605 1290.615 434.775 ;
        RECT 1290.905 289.425 1291.075 289.595 ;
      LAYER met1 ;
        RECT 1290.830 1076.340 1291.150 1076.400 ;
        RECT 1291.750 1076.340 1292.070 1076.400 ;
        RECT 1290.830 1076.200 1292.070 1076.340 ;
        RECT 1290.830 1076.140 1291.150 1076.200 ;
        RECT 1291.750 1076.140 1292.070 1076.200 ;
        RECT 1290.370 966.180 1290.690 966.240 ;
        RECT 1291.750 966.180 1292.070 966.240 ;
        RECT 1290.370 966.040 1292.070 966.180 ;
        RECT 1290.370 965.980 1290.690 966.040 ;
        RECT 1291.750 965.980 1292.070 966.040 ;
        RECT 1290.370 869.620 1290.690 869.680 ;
        RECT 1291.750 869.620 1292.070 869.680 ;
        RECT 1290.370 869.480 1292.070 869.620 ;
        RECT 1290.370 869.420 1290.690 869.480 ;
        RECT 1291.750 869.420 1292.070 869.480 ;
        RECT 1290.370 821.000 1290.690 821.060 ;
        RECT 1291.290 821.000 1291.610 821.060 ;
        RECT 1290.370 820.860 1291.610 821.000 ;
        RECT 1290.370 820.800 1290.690 820.860 ;
        RECT 1291.290 820.800 1291.610 820.860 ;
        RECT 1290.385 434.760 1290.675 434.805 ;
        RECT 1290.830 434.760 1291.150 434.820 ;
        RECT 1290.385 434.620 1291.150 434.760 ;
        RECT 1290.385 434.575 1290.675 434.620 ;
        RECT 1290.830 434.560 1291.150 434.620 ;
        RECT 1290.370 386.480 1290.690 386.540 ;
        RECT 1290.175 386.340 1290.690 386.480 ;
        RECT 1290.370 386.280 1290.690 386.340 ;
        RECT 1290.830 303.520 1291.150 303.580 ;
        RECT 1291.750 303.520 1292.070 303.580 ;
        RECT 1290.830 303.380 1292.070 303.520 ;
        RECT 1290.830 303.320 1291.150 303.380 ;
        RECT 1291.750 303.320 1292.070 303.380 ;
        RECT 1290.845 289.580 1291.135 289.625 ;
        RECT 1291.750 289.580 1292.070 289.640 ;
        RECT 1290.845 289.440 1292.070 289.580 ;
        RECT 1290.845 289.395 1291.135 289.440 ;
        RECT 1291.750 289.380 1292.070 289.440 ;
        RECT 1290.830 241.640 1291.150 241.700 ;
        RECT 1290.635 241.500 1291.150 241.640 ;
        RECT 1290.830 241.440 1291.150 241.500 ;
        RECT 1291.290 193.840 1291.610 194.100 ;
        RECT 1291.380 193.420 1291.520 193.840 ;
        RECT 1291.290 193.160 1291.610 193.420 ;
        RECT 1290.830 34.920 1291.150 34.980 ;
        RECT 1290.460 34.780 1291.150 34.920 ;
        RECT 1290.460 34.640 1290.600 34.780 ;
        RECT 1290.830 34.720 1291.150 34.780 ;
        RECT 1290.370 34.380 1290.690 34.640 ;
        RECT 1061.290 20.980 1061.610 21.040 ;
        RECT 1290.370 20.980 1290.690 21.040 ;
        RECT 1061.290 20.840 1290.690 20.980 ;
        RECT 1061.290 20.780 1061.610 20.840 ;
        RECT 1290.370 20.780 1290.690 20.840 ;
      LAYER via ;
        RECT 1290.860 1076.140 1291.120 1076.400 ;
        RECT 1291.780 1076.140 1292.040 1076.400 ;
        RECT 1290.400 965.980 1290.660 966.240 ;
        RECT 1291.780 965.980 1292.040 966.240 ;
        RECT 1290.400 869.420 1290.660 869.680 ;
        RECT 1291.780 869.420 1292.040 869.680 ;
        RECT 1290.400 820.800 1290.660 821.060 ;
        RECT 1291.320 820.800 1291.580 821.060 ;
        RECT 1290.860 434.560 1291.120 434.820 ;
        RECT 1290.400 386.280 1290.660 386.540 ;
        RECT 1290.860 303.320 1291.120 303.580 ;
        RECT 1291.780 303.320 1292.040 303.580 ;
        RECT 1291.780 289.380 1292.040 289.640 ;
        RECT 1290.860 241.440 1291.120 241.700 ;
        RECT 1291.320 193.840 1291.580 194.100 ;
        RECT 1291.320 193.160 1291.580 193.420 ;
        RECT 1290.860 34.720 1291.120 34.980 ;
        RECT 1290.400 34.380 1290.660 34.640 ;
        RECT 1061.320 20.780 1061.580 21.040 ;
        RECT 1290.400 20.780 1290.660 21.040 ;
      LAYER met2 ;
        RECT 1295.010 1220.330 1295.570 1228.680 ;
        RECT 1293.220 1220.190 1295.570 1220.330 ;
        RECT 1293.220 1207.410 1293.360 1220.190 ;
        RECT 1295.010 1219.680 1295.570 1220.190 ;
        RECT 1291.380 1207.270 1293.360 1207.410 ;
        RECT 1291.380 1097.250 1291.520 1207.270 ;
        RECT 1290.920 1097.110 1291.520 1097.250 ;
        RECT 1290.920 1076.430 1291.060 1097.110 ;
        RECT 1290.860 1076.110 1291.120 1076.430 ;
        RECT 1291.780 1076.110 1292.040 1076.430 ;
        RECT 1291.840 1027.890 1291.980 1076.110 ;
        RECT 1291.380 1027.750 1291.980 1027.890 ;
        RECT 1291.380 1014.405 1291.520 1027.750 ;
        RECT 1290.390 1014.035 1290.670 1014.405 ;
        RECT 1291.310 1014.035 1291.590 1014.405 ;
        RECT 1290.460 966.270 1290.600 1014.035 ;
        RECT 1290.400 965.950 1290.660 966.270 ;
        RECT 1291.780 965.950 1292.040 966.270 ;
        RECT 1291.840 931.330 1291.980 965.950 ;
        RECT 1291.380 931.190 1291.980 931.330 ;
        RECT 1291.380 917.845 1291.520 931.190 ;
        RECT 1290.390 917.475 1290.670 917.845 ;
        RECT 1291.310 917.475 1291.590 917.845 ;
        RECT 1290.460 869.710 1290.600 917.475 ;
        RECT 1290.400 869.390 1290.660 869.710 ;
        RECT 1291.780 869.390 1292.040 869.710 ;
        RECT 1291.840 834.770 1291.980 869.390 ;
        RECT 1291.380 834.630 1291.980 834.770 ;
        RECT 1291.380 821.090 1291.520 834.630 ;
        RECT 1290.400 820.770 1290.660 821.090 ;
        RECT 1291.320 820.770 1291.580 821.090 ;
        RECT 1290.460 773.005 1290.600 820.770 ;
        RECT 1290.390 772.635 1290.670 773.005 ;
        RECT 1291.770 772.635 1292.050 773.005 ;
        RECT 1291.840 738.210 1291.980 772.635 ;
        RECT 1291.380 738.070 1291.980 738.210 ;
        RECT 1291.380 700.130 1291.520 738.070 ;
        RECT 1290.460 699.990 1291.520 700.130 ;
        RECT 1290.460 676.445 1290.600 699.990 ;
        RECT 1290.390 676.075 1290.670 676.445 ;
        RECT 1291.770 676.075 1292.050 676.445 ;
        RECT 1291.840 641.650 1291.980 676.075 ;
        RECT 1291.380 641.510 1291.980 641.650 ;
        RECT 1291.380 603.570 1291.520 641.510 ;
        RECT 1290.460 603.430 1291.520 603.570 ;
        RECT 1290.460 579.885 1290.600 603.430 ;
        RECT 1290.390 579.515 1290.670 579.885 ;
        RECT 1291.770 579.515 1292.050 579.885 ;
        RECT 1291.840 545.090 1291.980 579.515 ;
        RECT 1291.380 544.950 1291.980 545.090 ;
        RECT 1291.380 507.010 1291.520 544.950 ;
        RECT 1290.460 506.870 1291.520 507.010 ;
        RECT 1290.460 483.325 1290.600 506.870 ;
        RECT 1290.390 482.955 1290.670 483.325 ;
        RECT 1291.770 482.955 1292.050 483.325 ;
        RECT 1291.840 448.530 1291.980 482.955 ;
        RECT 1290.920 448.390 1291.980 448.530 ;
        RECT 1290.920 434.850 1291.060 448.390 ;
        RECT 1290.860 434.530 1291.120 434.850 ;
        RECT 1290.400 386.250 1290.660 386.570 ;
        RECT 1290.460 351.290 1290.600 386.250 ;
        RECT 1290.460 351.150 1291.060 351.290 ;
        RECT 1290.920 303.610 1291.060 351.150 ;
        RECT 1290.860 303.290 1291.120 303.610 ;
        RECT 1291.780 303.290 1292.040 303.610 ;
        RECT 1291.840 289.670 1291.980 303.290 ;
        RECT 1291.780 289.350 1292.040 289.670 ;
        RECT 1290.860 241.410 1291.120 241.730 ;
        RECT 1290.920 226.170 1291.060 241.410 ;
        RECT 1290.920 226.030 1291.520 226.170 ;
        RECT 1291.380 194.130 1291.520 226.030 ;
        RECT 1291.320 193.810 1291.580 194.130 ;
        RECT 1291.320 193.130 1291.580 193.450 ;
        RECT 1291.380 192.850 1291.520 193.130 ;
        RECT 1290.920 192.710 1291.520 192.850 ;
        RECT 1290.920 158.170 1291.060 192.710 ;
        RECT 1290.920 158.030 1291.980 158.170 ;
        RECT 1291.840 110.570 1291.980 158.030 ;
        RECT 1290.920 110.430 1291.980 110.570 ;
        RECT 1290.920 35.010 1291.060 110.430 ;
        RECT 1290.860 34.690 1291.120 35.010 ;
        RECT 1290.400 34.350 1290.660 34.670 ;
        RECT 1290.460 21.070 1290.600 34.350 ;
        RECT 1061.320 20.750 1061.580 21.070 ;
        RECT 1290.400 20.750 1290.660 21.070 ;
        RECT 1061.380 2.400 1061.520 20.750 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
      LAYER via2 ;
        RECT 1290.390 1014.080 1290.670 1014.360 ;
        RECT 1291.310 1014.080 1291.590 1014.360 ;
        RECT 1290.390 917.520 1290.670 917.800 ;
        RECT 1291.310 917.520 1291.590 917.800 ;
        RECT 1290.390 772.680 1290.670 772.960 ;
        RECT 1291.770 772.680 1292.050 772.960 ;
        RECT 1290.390 676.120 1290.670 676.400 ;
        RECT 1291.770 676.120 1292.050 676.400 ;
        RECT 1290.390 579.560 1290.670 579.840 ;
        RECT 1291.770 579.560 1292.050 579.840 ;
        RECT 1290.390 483.000 1290.670 483.280 ;
        RECT 1291.770 483.000 1292.050 483.280 ;
      LAYER met3 ;
        RECT 1290.365 1014.370 1290.695 1014.385 ;
        RECT 1291.285 1014.370 1291.615 1014.385 ;
        RECT 1290.365 1014.070 1291.615 1014.370 ;
        RECT 1290.365 1014.055 1290.695 1014.070 ;
        RECT 1291.285 1014.055 1291.615 1014.070 ;
        RECT 1290.365 917.810 1290.695 917.825 ;
        RECT 1291.285 917.810 1291.615 917.825 ;
        RECT 1290.365 917.510 1291.615 917.810 ;
        RECT 1290.365 917.495 1290.695 917.510 ;
        RECT 1291.285 917.495 1291.615 917.510 ;
        RECT 1290.365 772.970 1290.695 772.985 ;
        RECT 1291.745 772.970 1292.075 772.985 ;
        RECT 1290.365 772.670 1292.075 772.970 ;
        RECT 1290.365 772.655 1290.695 772.670 ;
        RECT 1291.745 772.655 1292.075 772.670 ;
        RECT 1290.365 676.410 1290.695 676.425 ;
        RECT 1291.745 676.410 1292.075 676.425 ;
        RECT 1290.365 676.110 1292.075 676.410 ;
        RECT 1290.365 676.095 1290.695 676.110 ;
        RECT 1291.745 676.095 1292.075 676.110 ;
        RECT 1290.365 579.850 1290.695 579.865 ;
        RECT 1291.745 579.850 1292.075 579.865 ;
        RECT 1290.365 579.550 1292.075 579.850 ;
        RECT 1290.365 579.535 1290.695 579.550 ;
        RECT 1291.745 579.535 1292.075 579.550 ;
        RECT 1290.365 483.290 1290.695 483.305 ;
        RECT 1291.745 483.290 1292.075 483.305 ;
        RECT 1290.365 482.990 1292.075 483.290 ;
        RECT 1290.365 482.975 1290.695 482.990 ;
        RECT 1291.745 482.975 1292.075 482.990 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.230 19.620 1079.550 19.680 ;
        RECT 1305.090 19.620 1305.410 19.680 ;
        RECT 1079.230 19.480 1305.410 19.620 ;
        RECT 1079.230 19.420 1079.550 19.480 ;
        RECT 1305.090 19.420 1305.410 19.480 ;
      LAYER via ;
        RECT 1079.260 19.420 1079.520 19.680 ;
        RECT 1305.120 19.420 1305.380 19.680 ;
      LAYER met2 ;
        RECT 1304.210 1220.330 1304.770 1228.680 ;
        RECT 1304.210 1220.190 1305.320 1220.330 ;
        RECT 1304.210 1219.680 1304.770 1220.190 ;
        RECT 1305.180 19.710 1305.320 1220.190 ;
        RECT 1079.260 19.390 1079.520 19.710 ;
        RECT 1305.120 19.390 1305.380 19.710 ;
        RECT 1079.320 2.400 1079.460 19.390 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 19.960 1097.030 20.020 ;
        RECT 1311.990 19.960 1312.310 20.020 ;
        RECT 1096.710 19.820 1312.310 19.960 ;
        RECT 1096.710 19.760 1097.030 19.820 ;
        RECT 1311.990 19.760 1312.310 19.820 ;
      LAYER via ;
        RECT 1096.740 19.760 1097.000 20.020 ;
        RECT 1312.020 19.760 1312.280 20.020 ;
      LAYER met2 ;
        RECT 1313.410 1220.330 1313.970 1228.680 ;
        RECT 1312.080 1220.190 1313.970 1220.330 ;
        RECT 1312.080 20.050 1312.220 1220.190 ;
        RECT 1313.410 1219.680 1313.970 1220.190 ;
        RECT 1096.740 19.730 1097.000 20.050 ;
        RECT 1312.020 19.730 1312.280 20.050 ;
        RECT 1096.800 2.400 1096.940 19.730 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1318.965 1062.585 1319.135 1076.355 ;
        RECT 1318.965 741.625 1319.135 772.735 ;
        RECT 1318.965 662.405 1319.135 710.515 ;
        RECT 1318.965 571.285 1319.135 613.955 ;
        RECT 1318.965 484.245 1319.135 524.195 ;
        RECT 1318.505 241.485 1318.675 331.075 ;
      LAYER mcon ;
        RECT 1318.965 1076.185 1319.135 1076.355 ;
        RECT 1318.965 772.565 1319.135 772.735 ;
        RECT 1318.965 710.345 1319.135 710.515 ;
        RECT 1318.965 613.785 1319.135 613.955 ;
        RECT 1318.965 524.025 1319.135 524.195 ;
        RECT 1318.505 330.905 1318.675 331.075 ;
      LAYER met1 ;
        RECT 1318.890 1076.340 1319.210 1076.400 ;
        RECT 1318.695 1076.200 1319.210 1076.340 ;
        RECT 1318.890 1076.140 1319.210 1076.200 ;
        RECT 1318.890 1062.740 1319.210 1062.800 ;
        RECT 1318.695 1062.600 1319.210 1062.740 ;
        RECT 1318.890 1062.540 1319.210 1062.600 ;
        RECT 1317.970 966.180 1318.290 966.240 ;
        RECT 1318.890 966.180 1319.210 966.240 ;
        RECT 1317.970 966.040 1319.210 966.180 ;
        RECT 1317.970 965.980 1318.290 966.040 ;
        RECT 1318.890 965.980 1319.210 966.040 ;
        RECT 1317.970 869.620 1318.290 869.680 ;
        RECT 1318.890 869.620 1319.210 869.680 ;
        RECT 1317.970 869.480 1319.210 869.620 ;
        RECT 1317.970 869.420 1318.290 869.480 ;
        RECT 1318.890 869.420 1319.210 869.480 ;
        RECT 1318.890 772.720 1319.210 772.780 ;
        RECT 1318.695 772.580 1319.210 772.720 ;
        RECT 1318.890 772.520 1319.210 772.580 ;
        RECT 1318.890 741.780 1319.210 741.840 ;
        RECT 1318.695 741.640 1319.210 741.780 ;
        RECT 1318.890 741.580 1319.210 741.640 ;
        RECT 1318.890 710.500 1319.210 710.560 ;
        RECT 1318.695 710.360 1319.210 710.500 ;
        RECT 1318.890 710.300 1319.210 710.360 ;
        RECT 1318.890 662.560 1319.210 662.620 ;
        RECT 1318.695 662.420 1319.210 662.560 ;
        RECT 1318.890 662.360 1319.210 662.420 ;
        RECT 1318.890 613.940 1319.210 614.000 ;
        RECT 1318.695 613.800 1319.210 613.940 ;
        RECT 1318.890 613.740 1319.210 613.800 ;
        RECT 1318.890 571.440 1319.210 571.500 ;
        RECT 1318.695 571.300 1319.210 571.440 ;
        RECT 1318.890 571.240 1319.210 571.300 ;
        RECT 1318.890 524.180 1319.210 524.240 ;
        RECT 1318.695 524.040 1319.210 524.180 ;
        RECT 1318.890 523.980 1319.210 524.040 ;
        RECT 1318.890 484.400 1319.210 484.460 ;
        RECT 1318.695 484.260 1319.210 484.400 ;
        RECT 1318.890 484.200 1319.210 484.260 ;
        RECT 1318.445 331.060 1318.735 331.105 ;
        RECT 1318.890 331.060 1319.210 331.120 ;
        RECT 1318.445 330.920 1319.210 331.060 ;
        RECT 1318.445 330.875 1318.735 330.920 ;
        RECT 1318.890 330.860 1319.210 330.920 ;
        RECT 1318.430 241.640 1318.750 241.700 ;
        RECT 1318.235 241.500 1318.750 241.640 ;
        RECT 1318.430 241.440 1318.750 241.500 ;
        RECT 1114.650 20.640 1114.970 20.700 ;
        RECT 1318.430 20.640 1318.750 20.700 ;
        RECT 1114.650 20.500 1318.750 20.640 ;
        RECT 1114.650 20.440 1114.970 20.500 ;
        RECT 1318.430 20.440 1318.750 20.500 ;
      LAYER via ;
        RECT 1318.920 1076.140 1319.180 1076.400 ;
        RECT 1318.920 1062.540 1319.180 1062.800 ;
        RECT 1318.000 965.980 1318.260 966.240 ;
        RECT 1318.920 965.980 1319.180 966.240 ;
        RECT 1318.000 869.420 1318.260 869.680 ;
        RECT 1318.920 869.420 1319.180 869.680 ;
        RECT 1318.920 772.520 1319.180 772.780 ;
        RECT 1318.920 741.580 1319.180 741.840 ;
        RECT 1318.920 710.300 1319.180 710.560 ;
        RECT 1318.920 662.360 1319.180 662.620 ;
        RECT 1318.920 613.740 1319.180 614.000 ;
        RECT 1318.920 571.240 1319.180 571.500 ;
        RECT 1318.920 523.980 1319.180 524.240 ;
        RECT 1318.920 484.200 1319.180 484.460 ;
        RECT 1318.920 330.860 1319.180 331.120 ;
        RECT 1318.460 241.440 1318.720 241.700 ;
        RECT 1114.680 20.440 1114.940 20.700 ;
        RECT 1318.460 20.440 1318.720 20.700 ;
      LAYER met2 ;
        RECT 1322.150 1220.330 1322.710 1228.680 ;
        RECT 1320.820 1220.190 1322.710 1220.330 ;
        RECT 1320.820 1196.530 1320.960 1220.190 ;
        RECT 1322.150 1219.680 1322.710 1220.190 ;
        RECT 1318.980 1196.390 1320.960 1196.530 ;
        RECT 1318.980 1076.430 1319.120 1196.390 ;
        RECT 1318.920 1076.110 1319.180 1076.430 ;
        RECT 1318.920 1062.510 1319.180 1062.830 ;
        RECT 1318.980 1014.405 1319.120 1062.510 ;
        RECT 1317.990 1014.035 1318.270 1014.405 ;
        RECT 1318.910 1014.035 1319.190 1014.405 ;
        RECT 1318.060 966.270 1318.200 1014.035 ;
        RECT 1318.000 965.950 1318.260 966.270 ;
        RECT 1318.920 965.950 1319.180 966.270 ;
        RECT 1318.980 917.845 1319.120 965.950 ;
        RECT 1317.990 917.475 1318.270 917.845 ;
        RECT 1318.910 917.475 1319.190 917.845 ;
        RECT 1318.060 869.710 1318.200 917.475 ;
        RECT 1318.000 869.390 1318.260 869.710 ;
        RECT 1318.920 869.390 1319.180 869.710 ;
        RECT 1318.980 787.170 1319.120 869.390 ;
        RECT 1318.520 787.030 1319.120 787.170 ;
        RECT 1318.520 786.490 1318.660 787.030 ;
        RECT 1318.520 786.350 1319.120 786.490 ;
        RECT 1318.980 772.810 1319.120 786.350 ;
        RECT 1318.920 772.490 1319.180 772.810 ;
        RECT 1318.920 741.550 1319.180 741.870 ;
        RECT 1318.980 718.605 1319.120 741.550 ;
        RECT 1318.910 718.235 1319.190 718.605 ;
        RECT 1318.910 717.555 1319.190 717.925 ;
        RECT 1318.980 710.590 1319.120 717.555 ;
        RECT 1318.920 710.270 1319.180 710.590 ;
        RECT 1318.920 662.330 1319.180 662.650 ;
        RECT 1318.980 621.930 1319.120 662.330 ;
        RECT 1318.520 621.790 1319.120 621.930 ;
        RECT 1318.520 621.250 1318.660 621.790 ;
        RECT 1318.520 621.110 1319.120 621.250 ;
        RECT 1318.980 614.030 1319.120 621.110 ;
        RECT 1318.920 613.710 1319.180 614.030 ;
        RECT 1318.920 571.210 1319.180 571.530 ;
        RECT 1318.980 524.270 1319.120 571.210 ;
        RECT 1318.920 523.950 1319.180 524.270 ;
        RECT 1318.920 484.170 1319.180 484.490 ;
        RECT 1318.980 339.165 1319.120 484.170 ;
        RECT 1318.910 338.795 1319.190 339.165 ;
        RECT 1318.910 338.115 1319.190 338.485 ;
        RECT 1318.980 331.150 1319.120 338.115 ;
        RECT 1318.920 330.830 1319.180 331.150 ;
        RECT 1318.460 241.410 1318.720 241.730 ;
        RECT 1318.520 241.245 1318.660 241.410 ;
        RECT 1318.450 240.875 1318.730 241.245 ;
        RECT 1318.910 240.195 1319.190 240.565 ;
        RECT 1318.980 110.570 1319.120 240.195 ;
        RECT 1318.520 110.430 1319.120 110.570 ;
        RECT 1318.520 20.730 1318.660 110.430 ;
        RECT 1114.680 20.410 1114.940 20.730 ;
        RECT 1318.460 20.410 1318.720 20.730 ;
        RECT 1114.740 2.400 1114.880 20.410 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
      LAYER via2 ;
        RECT 1317.990 1014.080 1318.270 1014.360 ;
        RECT 1318.910 1014.080 1319.190 1014.360 ;
        RECT 1317.990 917.520 1318.270 917.800 ;
        RECT 1318.910 917.520 1319.190 917.800 ;
        RECT 1318.910 718.280 1319.190 718.560 ;
        RECT 1318.910 717.600 1319.190 717.880 ;
        RECT 1318.910 338.840 1319.190 339.120 ;
        RECT 1318.910 338.160 1319.190 338.440 ;
        RECT 1318.450 240.920 1318.730 241.200 ;
        RECT 1318.910 240.240 1319.190 240.520 ;
      LAYER met3 ;
        RECT 1317.965 1014.370 1318.295 1014.385 ;
        RECT 1318.885 1014.370 1319.215 1014.385 ;
        RECT 1317.965 1014.070 1319.215 1014.370 ;
        RECT 1317.965 1014.055 1318.295 1014.070 ;
        RECT 1318.885 1014.055 1319.215 1014.070 ;
        RECT 1317.965 917.810 1318.295 917.825 ;
        RECT 1318.885 917.810 1319.215 917.825 ;
        RECT 1317.965 917.510 1319.215 917.810 ;
        RECT 1317.965 917.495 1318.295 917.510 ;
        RECT 1318.885 917.495 1319.215 917.510 ;
        RECT 1318.885 718.570 1319.215 718.585 ;
        RECT 1318.670 718.255 1319.215 718.570 ;
        RECT 1318.670 717.905 1318.970 718.255 ;
        RECT 1318.670 717.590 1319.215 717.905 ;
        RECT 1318.885 717.575 1319.215 717.590 ;
        RECT 1318.885 339.130 1319.215 339.145 ;
        RECT 1318.885 338.830 1319.890 339.130 ;
        RECT 1318.885 338.815 1319.215 338.830 ;
        RECT 1318.885 338.450 1319.215 338.465 ;
        RECT 1319.590 338.450 1319.890 338.830 ;
        RECT 1318.885 338.150 1319.890 338.450 ;
        RECT 1318.885 338.135 1319.215 338.150 ;
        RECT 1318.425 241.210 1318.755 241.225 ;
        RECT 1317.750 240.910 1318.755 241.210 ;
        RECT 1317.750 240.530 1318.050 240.910 ;
        RECT 1318.425 240.895 1318.755 240.910 ;
        RECT 1318.885 240.530 1319.215 240.545 ;
        RECT 1317.750 240.230 1319.215 240.530 ;
        RECT 1318.885 240.215 1319.215 240.230 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1325.405 1062.585 1325.575 1077.035 ;
        RECT 1324.945 565.845 1325.115 613.955 ;
        RECT 1325.405 303.365 1325.575 331.075 ;
        RECT 1324.945 89.845 1325.115 137.955 ;
      LAYER mcon ;
        RECT 1325.405 1076.865 1325.575 1077.035 ;
        RECT 1324.945 613.785 1325.115 613.955 ;
        RECT 1325.405 330.905 1325.575 331.075 ;
        RECT 1324.945 137.785 1325.115 137.955 ;
      LAYER met1 ;
        RECT 1325.790 1174.260 1326.110 1174.320 ;
        RECT 1329.930 1174.260 1330.250 1174.320 ;
        RECT 1325.790 1174.120 1330.250 1174.260 ;
        RECT 1325.790 1174.060 1326.110 1174.120 ;
        RECT 1329.930 1174.060 1330.250 1174.120 ;
        RECT 1325.790 1111.020 1326.110 1111.080 ;
        RECT 1326.710 1111.020 1327.030 1111.080 ;
        RECT 1325.790 1110.880 1327.030 1111.020 ;
        RECT 1325.790 1110.820 1326.110 1110.880 ;
        RECT 1326.710 1110.820 1327.030 1110.880 ;
        RECT 1325.345 1077.020 1325.635 1077.065 ;
        RECT 1325.790 1077.020 1326.110 1077.080 ;
        RECT 1325.345 1076.880 1326.110 1077.020 ;
        RECT 1325.345 1076.835 1325.635 1076.880 ;
        RECT 1325.790 1076.820 1326.110 1076.880 ;
        RECT 1325.330 1062.740 1325.650 1062.800 ;
        RECT 1325.135 1062.600 1325.650 1062.740 ;
        RECT 1325.330 1062.540 1325.650 1062.600 ;
        RECT 1325.330 834.740 1325.650 835.000 ;
        RECT 1325.420 834.320 1325.560 834.740 ;
        RECT 1325.330 834.060 1325.650 834.320 ;
        RECT 1325.330 814.200 1325.650 814.260 ;
        RECT 1326.250 814.200 1326.570 814.260 ;
        RECT 1325.330 814.060 1326.570 814.200 ;
        RECT 1325.330 814.000 1325.650 814.060 ;
        RECT 1326.250 814.000 1326.570 814.060 ;
        RECT 1324.870 613.940 1325.190 614.000 ;
        RECT 1324.675 613.800 1325.190 613.940 ;
        RECT 1324.870 613.740 1325.190 613.800 ;
        RECT 1324.885 566.000 1325.175 566.045 ;
        RECT 1325.330 566.000 1325.650 566.060 ;
        RECT 1324.885 565.860 1325.650 566.000 ;
        RECT 1324.885 565.815 1325.175 565.860 ;
        RECT 1325.330 565.800 1325.650 565.860 ;
        RECT 1324.870 448.500 1325.190 448.760 ;
        RECT 1324.960 448.360 1325.100 448.500 ;
        RECT 1325.330 448.360 1325.650 448.420 ;
        RECT 1324.960 448.220 1325.650 448.360 ;
        RECT 1325.330 448.160 1325.650 448.220 ;
        RECT 1325.330 386.280 1325.650 386.540 ;
        RECT 1325.420 385.860 1325.560 386.280 ;
        RECT 1325.330 385.600 1325.650 385.860 ;
        RECT 1325.330 338.680 1325.650 338.940 ;
        RECT 1325.420 338.260 1325.560 338.680 ;
        RECT 1325.330 338.000 1325.650 338.260 ;
        RECT 1325.330 331.060 1325.650 331.120 ;
        RECT 1325.135 330.920 1325.650 331.060 ;
        RECT 1325.330 330.860 1325.650 330.920 ;
        RECT 1325.330 303.520 1325.650 303.580 ;
        RECT 1325.135 303.380 1325.650 303.520 ;
        RECT 1325.330 303.320 1325.650 303.380 ;
        RECT 1324.870 193.360 1325.190 193.420 ;
        RECT 1325.330 193.360 1325.650 193.420 ;
        RECT 1324.870 193.220 1325.650 193.360 ;
        RECT 1324.870 193.160 1325.190 193.220 ;
        RECT 1325.330 193.160 1325.650 193.220 ;
        RECT 1324.870 145.420 1325.190 145.480 ;
        RECT 1325.330 145.420 1325.650 145.480 ;
        RECT 1324.870 145.280 1325.650 145.420 ;
        RECT 1324.870 145.220 1325.190 145.280 ;
        RECT 1325.330 145.220 1325.650 145.280 ;
        RECT 1324.870 137.940 1325.190 138.000 ;
        RECT 1324.675 137.800 1325.190 137.940 ;
        RECT 1324.870 137.740 1325.190 137.800 ;
        RECT 1324.885 90.000 1325.175 90.045 ;
        RECT 1325.330 90.000 1325.650 90.060 ;
        RECT 1324.885 89.860 1325.650 90.000 ;
        RECT 1324.885 89.815 1325.175 89.860 ;
        RECT 1325.330 89.800 1325.650 89.860 ;
        RECT 1132.590 14.860 1132.910 14.920 ;
        RECT 1324.870 14.860 1325.190 14.920 ;
        RECT 1132.590 14.720 1325.190 14.860 ;
        RECT 1132.590 14.660 1132.910 14.720 ;
        RECT 1324.870 14.660 1325.190 14.720 ;
      LAYER via ;
        RECT 1325.820 1174.060 1326.080 1174.320 ;
        RECT 1329.960 1174.060 1330.220 1174.320 ;
        RECT 1325.820 1110.820 1326.080 1111.080 ;
        RECT 1326.740 1110.820 1327.000 1111.080 ;
        RECT 1325.820 1076.820 1326.080 1077.080 ;
        RECT 1325.360 1062.540 1325.620 1062.800 ;
        RECT 1325.360 834.740 1325.620 835.000 ;
        RECT 1325.360 834.060 1325.620 834.320 ;
        RECT 1325.360 814.000 1325.620 814.260 ;
        RECT 1326.280 814.000 1326.540 814.260 ;
        RECT 1324.900 613.740 1325.160 614.000 ;
        RECT 1325.360 565.800 1325.620 566.060 ;
        RECT 1324.900 448.500 1325.160 448.760 ;
        RECT 1325.360 448.160 1325.620 448.420 ;
        RECT 1325.360 386.280 1325.620 386.540 ;
        RECT 1325.360 385.600 1325.620 385.860 ;
        RECT 1325.360 338.680 1325.620 338.940 ;
        RECT 1325.360 338.000 1325.620 338.260 ;
        RECT 1325.360 330.860 1325.620 331.120 ;
        RECT 1325.360 303.320 1325.620 303.580 ;
        RECT 1324.900 193.160 1325.160 193.420 ;
        RECT 1325.360 193.160 1325.620 193.420 ;
        RECT 1324.900 145.220 1325.160 145.480 ;
        RECT 1325.360 145.220 1325.620 145.480 ;
        RECT 1324.900 137.740 1325.160 138.000 ;
        RECT 1325.360 89.800 1325.620 90.060 ;
        RECT 1132.620 14.660 1132.880 14.920 ;
        RECT 1324.900 14.660 1325.160 14.920 ;
      LAYER met2 ;
        RECT 1331.350 1220.330 1331.910 1228.680 ;
        RECT 1330.020 1220.190 1331.910 1220.330 ;
        RECT 1330.020 1174.350 1330.160 1220.190 ;
        RECT 1331.350 1219.680 1331.910 1220.190 ;
        RECT 1325.820 1174.030 1326.080 1174.350 ;
        RECT 1329.960 1174.030 1330.220 1174.350 ;
        RECT 1325.880 1159.245 1326.020 1174.030 ;
        RECT 1325.810 1158.875 1326.090 1159.245 ;
        RECT 1326.730 1158.875 1327.010 1159.245 ;
        RECT 1326.800 1111.110 1326.940 1158.875 ;
        RECT 1325.820 1110.790 1326.080 1111.110 ;
        RECT 1326.740 1110.790 1327.000 1111.110 ;
        RECT 1325.880 1077.110 1326.020 1110.790 ;
        RECT 1325.820 1076.790 1326.080 1077.110 ;
        RECT 1325.360 1062.510 1325.620 1062.830 ;
        RECT 1325.420 1028.570 1325.560 1062.510 ;
        RECT 1324.960 1028.430 1325.560 1028.570 ;
        RECT 1324.960 1027.890 1325.100 1028.430 ;
        RECT 1324.960 1027.750 1325.560 1027.890 ;
        RECT 1325.420 932.010 1325.560 1027.750 ;
        RECT 1324.960 931.870 1325.560 932.010 ;
        RECT 1324.960 931.330 1325.100 931.870 ;
        RECT 1324.960 931.190 1325.560 931.330 ;
        RECT 1325.420 835.030 1325.560 931.190 ;
        RECT 1325.360 834.710 1325.620 835.030 ;
        RECT 1325.360 834.030 1325.620 834.350 ;
        RECT 1325.420 814.290 1325.560 834.030 ;
        RECT 1325.360 813.970 1325.620 814.290 ;
        RECT 1326.280 813.970 1326.540 814.290 ;
        RECT 1326.340 724.725 1326.480 813.970 ;
        RECT 1325.350 724.355 1325.630 724.725 ;
        RECT 1326.270 724.355 1326.550 724.725 ;
        RECT 1325.420 723.930 1325.560 724.355 ;
        RECT 1325.420 723.790 1326.480 723.930 ;
        RECT 1326.340 676.445 1326.480 723.790 ;
        RECT 1325.350 676.075 1325.630 676.445 ;
        RECT 1326.270 676.075 1326.550 676.445 ;
        RECT 1325.420 644.370 1325.560 676.075 ;
        RECT 1324.960 644.230 1325.560 644.370 ;
        RECT 1324.960 614.030 1325.100 644.230 ;
        RECT 1324.900 613.710 1325.160 614.030 ;
        RECT 1325.360 565.770 1325.620 566.090 ;
        RECT 1325.420 554.610 1325.560 565.770 ;
        RECT 1324.960 554.470 1325.560 554.610 ;
        RECT 1324.960 448.790 1325.100 554.470 ;
        RECT 1324.900 448.470 1325.160 448.790 ;
        RECT 1325.360 448.130 1325.620 448.450 ;
        RECT 1325.420 386.570 1325.560 448.130 ;
        RECT 1325.360 386.250 1325.620 386.570 ;
        RECT 1325.360 385.570 1325.620 385.890 ;
        RECT 1325.420 338.970 1325.560 385.570 ;
        RECT 1325.360 338.650 1325.620 338.970 ;
        RECT 1325.360 337.970 1325.620 338.290 ;
        RECT 1325.420 331.150 1325.560 337.970 ;
        RECT 1325.360 330.830 1325.620 331.150 ;
        RECT 1325.360 303.290 1325.620 303.610 ;
        RECT 1325.420 255.410 1325.560 303.290 ;
        RECT 1324.960 255.270 1325.560 255.410 ;
        RECT 1324.960 193.450 1325.100 255.270 ;
        RECT 1324.900 193.130 1325.160 193.450 ;
        RECT 1325.360 193.130 1325.620 193.450 ;
        RECT 1325.420 145.510 1325.560 193.130 ;
        RECT 1324.900 145.190 1325.160 145.510 ;
        RECT 1325.360 145.190 1325.620 145.510 ;
        RECT 1324.960 138.030 1325.100 145.190 ;
        RECT 1324.900 137.710 1325.160 138.030 ;
        RECT 1325.360 89.770 1325.620 90.090 ;
        RECT 1325.420 62.290 1325.560 89.770 ;
        RECT 1324.960 62.150 1325.560 62.290 ;
        RECT 1324.960 14.950 1325.100 62.150 ;
        RECT 1132.620 14.630 1132.880 14.950 ;
        RECT 1324.900 14.630 1325.160 14.950 ;
        RECT 1132.680 2.400 1132.820 14.630 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
      LAYER via2 ;
        RECT 1325.810 1158.920 1326.090 1159.200 ;
        RECT 1326.730 1158.920 1327.010 1159.200 ;
        RECT 1325.350 724.400 1325.630 724.680 ;
        RECT 1326.270 724.400 1326.550 724.680 ;
        RECT 1325.350 676.120 1325.630 676.400 ;
        RECT 1326.270 676.120 1326.550 676.400 ;
      LAYER met3 ;
        RECT 1325.785 1159.210 1326.115 1159.225 ;
        RECT 1326.705 1159.210 1327.035 1159.225 ;
        RECT 1325.785 1158.910 1327.035 1159.210 ;
        RECT 1325.785 1158.895 1326.115 1158.910 ;
        RECT 1326.705 1158.895 1327.035 1158.910 ;
        RECT 1325.325 724.690 1325.655 724.705 ;
        RECT 1326.245 724.690 1326.575 724.705 ;
        RECT 1325.325 724.390 1326.575 724.690 ;
        RECT 1325.325 724.375 1325.655 724.390 ;
        RECT 1326.245 724.375 1326.575 724.390 ;
        RECT 1325.325 676.410 1325.655 676.425 ;
        RECT 1326.245 676.410 1326.575 676.425 ;
        RECT 1325.325 676.110 1326.575 676.410 ;
        RECT 1325.325 676.095 1325.655 676.110 ;
        RECT 1326.245 676.095 1326.575 676.110 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 15.200 1150.850 15.260 ;
        RECT 1339.130 15.200 1339.450 15.260 ;
        RECT 1150.530 15.060 1339.450 15.200 ;
        RECT 1150.530 15.000 1150.850 15.060 ;
        RECT 1339.130 15.000 1339.450 15.060 ;
      LAYER via ;
        RECT 1150.560 15.000 1150.820 15.260 ;
        RECT 1339.160 15.000 1339.420 15.260 ;
      LAYER met2 ;
        RECT 1340.550 1220.330 1341.110 1228.680 ;
        RECT 1339.220 1220.190 1341.110 1220.330 ;
        RECT 1339.220 15.290 1339.360 1220.190 ;
        RECT 1340.550 1219.680 1341.110 1220.190 ;
        RECT 1150.560 14.970 1150.820 15.290 ;
        RECT 1339.160 14.970 1339.420 15.290 ;
        RECT 1150.620 2.400 1150.760 14.970 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 36.280 669.230 36.340 ;
        RECT 1090.730 36.280 1091.050 36.340 ;
        RECT 668.910 36.140 1091.050 36.280 ;
        RECT 668.910 36.080 669.230 36.140 ;
        RECT 1090.730 36.080 1091.050 36.140 ;
      LAYER via ;
        RECT 668.940 36.080 669.200 36.340 ;
        RECT 1090.760 36.080 1091.020 36.340 ;
      LAYER met2 ;
        RECT 1093.070 1220.330 1093.630 1228.680 ;
        RECT 1091.740 1220.190 1093.630 1220.330 ;
        RECT 1091.740 1196.700 1091.880 1220.190 ;
        RECT 1093.070 1219.680 1093.630 1220.190 ;
        RECT 1090.820 1196.560 1091.880 1196.700 ;
        RECT 1090.820 36.370 1090.960 1196.560 ;
        RECT 668.940 36.050 669.200 36.370 ;
        RECT 1090.760 36.050 1091.020 36.370 ;
        RECT 669.000 2.400 669.140 36.050 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.030 1193.640 1346.350 1193.700 ;
        RECT 1347.870 1193.640 1348.190 1193.700 ;
        RECT 1346.030 1193.500 1348.190 1193.640 ;
        RECT 1346.030 1193.440 1346.350 1193.500 ;
        RECT 1347.870 1193.440 1348.190 1193.500 ;
        RECT 1168.470 24.040 1168.790 24.100 ;
        RECT 1346.030 24.040 1346.350 24.100 ;
        RECT 1168.470 23.900 1346.350 24.040 ;
        RECT 1168.470 23.840 1168.790 23.900 ;
        RECT 1346.030 23.840 1346.350 23.900 ;
      LAYER via ;
        RECT 1346.060 1193.440 1346.320 1193.700 ;
        RECT 1347.900 1193.440 1348.160 1193.700 ;
        RECT 1168.500 23.840 1168.760 24.100 ;
        RECT 1346.060 23.840 1346.320 24.100 ;
      LAYER met2 ;
        RECT 1349.750 1220.330 1350.310 1228.680 ;
        RECT 1347.960 1220.190 1350.310 1220.330 ;
        RECT 1347.960 1193.730 1348.100 1220.190 ;
        RECT 1349.750 1219.680 1350.310 1220.190 ;
        RECT 1346.060 1193.410 1346.320 1193.730 ;
        RECT 1347.900 1193.410 1348.160 1193.730 ;
        RECT 1346.120 24.130 1346.260 1193.410 ;
        RECT 1168.500 23.810 1168.760 24.130 ;
        RECT 1346.060 23.810 1346.320 24.130 ;
        RECT 1168.560 2.400 1168.700 23.810 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1353.005 1062.585 1353.175 1077.035 ;
        RECT 1352.545 469.285 1352.715 517.395 ;
        RECT 1352.545 379.525 1352.715 427.635 ;
        RECT 1353.005 241.485 1353.175 255.935 ;
        RECT 1353.005 138.125 1353.175 159.375 ;
        RECT 1352.545 48.365 1352.715 96.815 ;
      LAYER mcon ;
        RECT 1353.005 1076.865 1353.175 1077.035 ;
        RECT 1352.545 517.225 1352.715 517.395 ;
        RECT 1352.545 427.465 1352.715 427.635 ;
        RECT 1353.005 255.765 1353.175 255.935 ;
        RECT 1353.005 159.205 1353.175 159.375 ;
        RECT 1352.545 96.645 1352.715 96.815 ;
      LAYER met1 ;
        RECT 1352.470 1196.700 1352.790 1196.760 ;
        RECT 1357.530 1196.700 1357.850 1196.760 ;
        RECT 1352.470 1196.560 1357.850 1196.700 ;
        RECT 1352.470 1196.500 1352.790 1196.560 ;
        RECT 1357.530 1196.500 1357.850 1196.560 ;
        RECT 1352.470 1172.900 1352.790 1172.960 ;
        RECT 1353.390 1172.900 1353.710 1172.960 ;
        RECT 1352.470 1172.760 1353.710 1172.900 ;
        RECT 1352.470 1172.700 1352.790 1172.760 ;
        RECT 1353.390 1172.700 1353.710 1172.760 ;
        RECT 1352.945 1077.020 1353.235 1077.065 ;
        RECT 1353.390 1077.020 1353.710 1077.080 ;
        RECT 1352.945 1076.880 1353.710 1077.020 ;
        RECT 1352.945 1076.835 1353.235 1076.880 ;
        RECT 1353.390 1076.820 1353.710 1076.880 ;
        RECT 1352.930 1062.740 1353.250 1062.800 ;
        RECT 1352.735 1062.600 1353.250 1062.740 ;
        RECT 1352.930 1062.540 1353.250 1062.600 ;
        RECT 1352.930 834.740 1353.250 835.000 ;
        RECT 1353.020 834.320 1353.160 834.740 ;
        RECT 1352.930 834.060 1353.250 834.320 ;
        RECT 1352.930 814.200 1353.250 814.260 ;
        RECT 1353.850 814.200 1354.170 814.260 ;
        RECT 1352.930 814.060 1354.170 814.200 ;
        RECT 1352.930 814.000 1353.250 814.060 ;
        RECT 1353.850 814.000 1354.170 814.060 ;
        RECT 1352.470 517.380 1352.790 517.440 ;
        RECT 1352.275 517.240 1352.790 517.380 ;
        RECT 1352.470 517.180 1352.790 517.240 ;
        RECT 1352.485 469.440 1352.775 469.485 ;
        RECT 1352.930 469.440 1353.250 469.500 ;
        RECT 1352.485 469.300 1353.250 469.440 ;
        RECT 1352.485 469.255 1352.775 469.300 ;
        RECT 1352.930 469.240 1353.250 469.300 ;
        RECT 1352.470 427.620 1352.790 427.680 ;
        RECT 1352.275 427.480 1352.790 427.620 ;
        RECT 1352.470 427.420 1352.790 427.480 ;
        RECT 1352.485 379.680 1352.775 379.725 ;
        RECT 1352.930 379.680 1353.250 379.740 ;
        RECT 1352.485 379.540 1353.250 379.680 ;
        RECT 1352.485 379.495 1352.775 379.540 ;
        RECT 1352.930 379.480 1353.250 379.540 ;
        RECT 1352.930 255.920 1353.250 255.980 ;
        RECT 1352.735 255.780 1353.250 255.920 ;
        RECT 1352.930 255.720 1353.250 255.780 ;
        RECT 1352.930 241.640 1353.250 241.700 ;
        RECT 1352.735 241.500 1353.250 241.640 ;
        RECT 1352.930 241.440 1353.250 241.500 ;
        RECT 1352.930 159.360 1353.250 159.420 ;
        RECT 1352.735 159.220 1353.250 159.360 ;
        RECT 1352.930 159.160 1353.250 159.220 ;
        RECT 1352.930 138.280 1353.250 138.340 ;
        RECT 1352.735 138.140 1353.250 138.280 ;
        RECT 1352.930 138.080 1353.250 138.140 ;
        RECT 1352.485 96.800 1352.775 96.845 ;
        RECT 1352.930 96.800 1353.250 96.860 ;
        RECT 1352.485 96.660 1353.250 96.800 ;
        RECT 1352.485 96.615 1352.775 96.660 ;
        RECT 1352.930 96.600 1353.250 96.660 ;
        RECT 1352.485 48.520 1352.775 48.565 ;
        RECT 1352.930 48.520 1353.250 48.580 ;
        RECT 1352.485 48.380 1353.250 48.520 ;
        RECT 1352.485 48.335 1352.775 48.380 ;
        RECT 1352.930 48.320 1353.250 48.380 ;
        RECT 1185.950 24.380 1186.270 24.440 ;
        RECT 1352.930 24.380 1353.250 24.440 ;
        RECT 1185.950 24.240 1353.250 24.380 ;
        RECT 1185.950 24.180 1186.270 24.240 ;
        RECT 1352.930 24.180 1353.250 24.240 ;
      LAYER via ;
        RECT 1352.500 1196.500 1352.760 1196.760 ;
        RECT 1357.560 1196.500 1357.820 1196.760 ;
        RECT 1352.500 1172.700 1352.760 1172.960 ;
        RECT 1353.420 1172.700 1353.680 1172.960 ;
        RECT 1353.420 1076.820 1353.680 1077.080 ;
        RECT 1352.960 1062.540 1353.220 1062.800 ;
        RECT 1352.960 834.740 1353.220 835.000 ;
        RECT 1352.960 834.060 1353.220 834.320 ;
        RECT 1352.960 814.000 1353.220 814.260 ;
        RECT 1353.880 814.000 1354.140 814.260 ;
        RECT 1352.500 517.180 1352.760 517.440 ;
        RECT 1352.960 469.240 1353.220 469.500 ;
        RECT 1352.500 427.420 1352.760 427.680 ;
        RECT 1352.960 379.480 1353.220 379.740 ;
        RECT 1352.960 255.720 1353.220 255.980 ;
        RECT 1352.960 241.440 1353.220 241.700 ;
        RECT 1352.960 159.160 1353.220 159.420 ;
        RECT 1352.960 138.080 1353.220 138.340 ;
        RECT 1352.960 96.600 1353.220 96.860 ;
        RECT 1352.960 48.320 1353.220 48.580 ;
        RECT 1185.980 24.180 1186.240 24.440 ;
        RECT 1352.960 24.180 1353.220 24.440 ;
      LAYER met2 ;
        RECT 1358.950 1220.330 1359.510 1228.680 ;
        RECT 1357.620 1220.190 1359.510 1220.330 ;
        RECT 1357.620 1196.790 1357.760 1220.190 ;
        RECT 1358.950 1219.680 1359.510 1220.190 ;
        RECT 1352.500 1196.470 1352.760 1196.790 ;
        RECT 1357.560 1196.470 1357.820 1196.790 ;
        RECT 1352.560 1172.990 1352.700 1196.470 ;
        RECT 1352.500 1172.670 1352.760 1172.990 ;
        RECT 1353.420 1172.670 1353.680 1172.990 ;
        RECT 1353.480 1159.245 1353.620 1172.670 ;
        RECT 1352.490 1158.875 1352.770 1159.245 ;
        RECT 1353.410 1158.875 1353.690 1159.245 ;
        RECT 1352.560 1121.730 1352.700 1158.875 ;
        RECT 1352.560 1121.590 1353.620 1121.730 ;
        RECT 1353.480 1077.110 1353.620 1121.590 ;
        RECT 1353.420 1076.790 1353.680 1077.110 ;
        RECT 1352.960 1062.510 1353.220 1062.830 ;
        RECT 1353.020 1028.570 1353.160 1062.510 ;
        RECT 1352.560 1028.430 1353.160 1028.570 ;
        RECT 1352.560 1027.890 1352.700 1028.430 ;
        RECT 1352.560 1027.750 1353.160 1027.890 ;
        RECT 1353.020 932.010 1353.160 1027.750 ;
        RECT 1352.560 931.870 1353.160 932.010 ;
        RECT 1352.560 931.330 1352.700 931.870 ;
        RECT 1352.560 931.190 1353.160 931.330 ;
        RECT 1353.020 835.030 1353.160 931.190 ;
        RECT 1352.960 834.710 1353.220 835.030 ;
        RECT 1352.960 834.030 1353.220 834.350 ;
        RECT 1353.020 814.290 1353.160 834.030 ;
        RECT 1352.960 813.970 1353.220 814.290 ;
        RECT 1353.880 813.970 1354.140 814.290 ;
        RECT 1353.940 724.725 1354.080 813.970 ;
        RECT 1352.490 724.355 1352.770 724.725 ;
        RECT 1353.870 724.355 1354.150 724.725 ;
        RECT 1352.560 676.330 1352.700 724.355 ;
        RECT 1352.560 676.190 1353.160 676.330 ;
        RECT 1353.020 641.650 1353.160 676.190 ;
        RECT 1352.560 641.510 1353.160 641.650 ;
        RECT 1352.560 579.770 1352.700 641.510 ;
        RECT 1352.560 579.630 1353.160 579.770 ;
        RECT 1353.020 548.490 1353.160 579.630 ;
        RECT 1352.560 548.350 1353.160 548.490 ;
        RECT 1352.560 517.470 1352.700 548.350 ;
        RECT 1352.500 517.150 1352.760 517.470 ;
        RECT 1352.960 469.210 1353.220 469.530 ;
        RECT 1353.020 451.930 1353.160 469.210 ;
        RECT 1352.560 451.790 1353.160 451.930 ;
        RECT 1352.560 427.710 1352.700 451.790 ;
        RECT 1352.500 427.390 1352.760 427.710 ;
        RECT 1352.960 379.450 1353.220 379.770 ;
        RECT 1353.020 351.970 1353.160 379.450 ;
        RECT 1352.560 351.830 1353.160 351.970 ;
        RECT 1352.560 351.290 1352.700 351.830 ;
        RECT 1352.560 351.150 1353.160 351.290 ;
        RECT 1353.020 256.010 1353.160 351.150 ;
        RECT 1352.960 255.690 1353.220 256.010 ;
        RECT 1352.960 241.410 1353.220 241.730 ;
        RECT 1353.020 159.450 1353.160 241.410 ;
        RECT 1352.960 159.130 1353.220 159.450 ;
        RECT 1352.960 138.050 1353.220 138.370 ;
        RECT 1353.020 96.890 1353.160 138.050 ;
        RECT 1352.960 96.570 1353.220 96.890 ;
        RECT 1352.960 48.290 1353.220 48.610 ;
        RECT 1353.020 24.470 1353.160 48.290 ;
        RECT 1185.980 24.150 1186.240 24.470 ;
        RECT 1352.960 24.150 1353.220 24.470 ;
        RECT 1186.040 2.400 1186.180 24.150 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 1352.490 1158.920 1352.770 1159.200 ;
        RECT 1353.410 1158.920 1353.690 1159.200 ;
        RECT 1352.490 724.400 1352.770 724.680 ;
        RECT 1353.870 724.400 1354.150 724.680 ;
      LAYER met3 ;
        RECT 1352.465 1159.210 1352.795 1159.225 ;
        RECT 1353.385 1159.210 1353.715 1159.225 ;
        RECT 1352.465 1158.910 1353.715 1159.210 ;
        RECT 1352.465 1158.895 1352.795 1158.910 ;
        RECT 1353.385 1158.895 1353.715 1158.910 ;
        RECT 1352.465 724.690 1352.795 724.705 ;
        RECT 1353.845 724.690 1354.175 724.705 ;
        RECT 1352.465 724.390 1354.175 724.690 ;
        RECT 1352.465 724.375 1352.795 724.390 ;
        RECT 1353.845 724.375 1354.175 724.390 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 1209.280 1207.430 1209.340 ;
        RECT 1368.110 1209.280 1368.430 1209.340 ;
        RECT 1207.110 1209.140 1368.430 1209.280 ;
        RECT 1207.110 1209.080 1207.430 1209.140 ;
        RECT 1368.110 1209.080 1368.430 1209.140 ;
        RECT 1203.890 18.940 1204.210 19.000 ;
        RECT 1207.110 18.940 1207.430 19.000 ;
        RECT 1203.890 18.800 1207.430 18.940 ;
        RECT 1203.890 18.740 1204.210 18.800 ;
        RECT 1207.110 18.740 1207.430 18.800 ;
      LAYER via ;
        RECT 1207.140 1209.080 1207.400 1209.340 ;
        RECT 1368.140 1209.080 1368.400 1209.340 ;
        RECT 1203.920 18.740 1204.180 19.000 ;
        RECT 1207.140 18.740 1207.400 19.000 ;
      LAYER met2 ;
        RECT 1368.150 1219.680 1368.710 1228.680 ;
        RECT 1368.200 1209.370 1368.340 1219.680 ;
        RECT 1207.140 1209.050 1207.400 1209.370 ;
        RECT 1368.140 1209.050 1368.400 1209.370 ;
        RECT 1207.200 19.030 1207.340 1209.050 ;
        RECT 1203.920 18.710 1204.180 19.030 ;
        RECT 1207.140 18.710 1207.400 19.030 ;
        RECT 1203.980 2.400 1204.120 18.710 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1268.825 16.405 1274.055 16.575 ;
        RECT 1284.465 16.405 1284.635 19.295 ;
      LAYER mcon ;
        RECT 1284.465 19.125 1284.635 19.295 ;
        RECT 1273.885 16.405 1274.055 16.575 ;
      LAYER met1 ;
        RECT 1342.350 1210.300 1342.670 1210.360 ;
        RECT 1377.310 1210.300 1377.630 1210.360 ;
        RECT 1342.350 1210.160 1377.630 1210.300 ;
        RECT 1342.350 1210.100 1342.670 1210.160 ;
        RECT 1377.310 1210.100 1377.630 1210.160 ;
        RECT 1341.430 20.300 1341.750 20.360 ;
        RECT 1312.540 20.160 1341.750 20.300 ;
        RECT 1312.540 19.620 1312.680 20.160 ;
        RECT 1341.430 20.100 1341.750 20.160 ;
        RECT 1305.640 19.480 1312.680 19.620 ;
        RECT 1284.405 19.280 1284.695 19.325 ;
        RECT 1305.640 19.280 1305.780 19.480 ;
        RECT 1284.405 19.140 1305.780 19.280 ;
        RECT 1284.405 19.095 1284.695 19.140 ;
        RECT 1268.765 16.560 1269.055 16.605 ;
        RECT 1245.840 16.420 1269.055 16.560 ;
        RECT 1221.830 16.220 1222.150 16.280 ;
        RECT 1245.840 16.220 1245.980 16.420 ;
        RECT 1268.765 16.375 1269.055 16.420 ;
        RECT 1273.825 16.560 1274.115 16.605 ;
        RECT 1284.405 16.560 1284.695 16.605 ;
        RECT 1273.825 16.420 1284.695 16.560 ;
        RECT 1273.825 16.375 1274.115 16.420 ;
        RECT 1284.405 16.375 1284.695 16.420 ;
        RECT 1221.830 16.080 1245.980 16.220 ;
        RECT 1221.830 16.020 1222.150 16.080 ;
      LAYER via ;
        RECT 1342.380 1210.100 1342.640 1210.360 ;
        RECT 1377.340 1210.100 1377.600 1210.360 ;
        RECT 1341.460 20.100 1341.720 20.360 ;
        RECT 1221.860 16.020 1222.120 16.280 ;
      LAYER met2 ;
        RECT 1377.350 1219.680 1377.910 1228.680 ;
        RECT 1377.400 1210.390 1377.540 1219.680 ;
        RECT 1342.380 1210.070 1342.640 1210.390 ;
        RECT 1377.340 1210.070 1377.600 1210.390 ;
        RECT 1342.440 1208.770 1342.580 1210.070 ;
        RECT 1341.980 1208.630 1342.580 1208.770 ;
        RECT 1341.980 20.810 1342.120 1208.630 ;
        RECT 1341.520 20.670 1342.120 20.810 ;
        RECT 1341.520 20.390 1341.660 20.670 ;
        RECT 1341.460 20.070 1341.720 20.390 ;
        RECT 1221.860 15.990 1222.120 16.310 ;
        RECT 1221.920 2.400 1222.060 15.990 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1240.765 959.225 1240.935 1007.335 ;
        RECT 1241.685 766.105 1241.855 814.215 ;
        RECT 1241.685 669.545 1241.855 717.655 ;
        RECT 1241.685 572.645 1241.855 620.755 ;
        RECT 1241.685 476.085 1241.855 524.195 ;
        RECT 1241.685 379.525 1241.855 427.635 ;
        RECT 1241.685 282.965 1241.855 331.075 ;
        RECT 1241.685 186.405 1241.855 234.515 ;
        RECT 1239.845 48.365 1240.015 96.475 ;
      LAYER mcon ;
        RECT 1240.765 1007.165 1240.935 1007.335 ;
        RECT 1241.685 814.045 1241.855 814.215 ;
        RECT 1241.685 717.485 1241.855 717.655 ;
        RECT 1241.685 620.585 1241.855 620.755 ;
        RECT 1241.685 524.025 1241.855 524.195 ;
        RECT 1241.685 427.465 1241.855 427.635 ;
        RECT 1241.685 330.905 1241.855 331.075 ;
        RECT 1241.685 234.345 1241.855 234.515 ;
        RECT 1239.845 96.305 1240.015 96.475 ;
      LAYER met1 ;
        RECT 1241.610 1212.340 1241.930 1212.400 ;
        RECT 1386.510 1212.340 1386.830 1212.400 ;
        RECT 1241.610 1212.200 1386.830 1212.340 ;
        RECT 1241.610 1212.140 1241.930 1212.200 ;
        RECT 1386.510 1212.140 1386.830 1212.200 ;
        RECT 1240.690 1152.500 1241.010 1152.560 ;
        RECT 1241.150 1152.500 1241.470 1152.560 ;
        RECT 1240.690 1152.360 1241.470 1152.500 ;
        RECT 1240.690 1152.300 1241.010 1152.360 ;
        RECT 1241.150 1152.300 1241.470 1152.360 ;
        RECT 1239.770 1104.220 1240.090 1104.280 ;
        RECT 1241.610 1104.220 1241.930 1104.280 ;
        RECT 1239.770 1104.080 1241.930 1104.220 ;
        RECT 1239.770 1104.020 1240.090 1104.080 ;
        RECT 1241.610 1104.020 1241.930 1104.080 ;
        RECT 1240.690 1055.940 1241.010 1056.000 ;
        RECT 1241.150 1055.940 1241.470 1056.000 ;
        RECT 1240.690 1055.800 1241.470 1055.940 ;
        RECT 1240.690 1055.740 1241.010 1055.800 ;
        RECT 1241.150 1055.740 1241.470 1055.800 ;
        RECT 1240.690 1014.460 1241.010 1014.520 ;
        RECT 1241.610 1014.460 1241.930 1014.520 ;
        RECT 1240.690 1014.320 1241.930 1014.460 ;
        RECT 1240.690 1014.260 1241.010 1014.320 ;
        RECT 1241.610 1014.260 1241.930 1014.320 ;
        RECT 1240.705 1007.320 1240.995 1007.365 ;
        RECT 1241.610 1007.320 1241.930 1007.380 ;
        RECT 1240.705 1007.180 1241.930 1007.320 ;
        RECT 1240.705 1007.135 1240.995 1007.180 ;
        RECT 1241.610 1007.120 1241.930 1007.180 ;
        RECT 1240.690 959.380 1241.010 959.440 ;
        RECT 1240.495 959.240 1241.010 959.380 ;
        RECT 1240.690 959.180 1241.010 959.240 ;
        RECT 1240.690 917.900 1241.010 917.960 ;
        RECT 1241.610 917.900 1241.930 917.960 ;
        RECT 1240.690 917.760 1241.930 917.900 ;
        RECT 1240.690 917.700 1241.010 917.760 ;
        RECT 1241.610 917.700 1241.930 917.760 ;
        RECT 1240.690 910.760 1241.010 910.820 ;
        RECT 1241.610 910.760 1241.930 910.820 ;
        RECT 1240.690 910.620 1241.930 910.760 ;
        RECT 1240.690 910.560 1241.010 910.620 ;
        RECT 1241.610 910.560 1241.930 910.620 ;
        RECT 1241.610 814.200 1241.930 814.260 ;
        RECT 1241.415 814.060 1241.930 814.200 ;
        RECT 1241.610 814.000 1241.930 814.060 ;
        RECT 1241.610 766.260 1241.930 766.320 ;
        RECT 1241.415 766.120 1241.930 766.260 ;
        RECT 1241.610 766.060 1241.930 766.120 ;
        RECT 1241.610 717.640 1241.930 717.700 ;
        RECT 1241.415 717.500 1241.930 717.640 ;
        RECT 1241.610 717.440 1241.930 717.500 ;
        RECT 1241.610 669.700 1241.930 669.760 ;
        RECT 1241.415 669.560 1241.930 669.700 ;
        RECT 1241.610 669.500 1241.930 669.560 ;
        RECT 1241.610 620.740 1241.930 620.800 ;
        RECT 1241.415 620.600 1241.930 620.740 ;
        RECT 1241.610 620.540 1241.930 620.600 ;
        RECT 1241.610 572.800 1241.930 572.860 ;
        RECT 1241.415 572.660 1241.930 572.800 ;
        RECT 1241.610 572.600 1241.930 572.660 ;
        RECT 1241.610 524.180 1241.930 524.240 ;
        RECT 1241.415 524.040 1241.930 524.180 ;
        RECT 1241.610 523.980 1241.930 524.040 ;
        RECT 1241.610 476.240 1241.930 476.300 ;
        RECT 1241.415 476.100 1241.930 476.240 ;
        RECT 1241.610 476.040 1241.930 476.100 ;
        RECT 1241.610 427.620 1241.930 427.680 ;
        RECT 1241.415 427.480 1241.930 427.620 ;
        RECT 1241.610 427.420 1241.930 427.480 ;
        RECT 1241.610 379.680 1241.930 379.740 ;
        RECT 1241.415 379.540 1241.930 379.680 ;
        RECT 1241.610 379.480 1241.930 379.540 ;
        RECT 1241.610 338.680 1241.930 338.940 ;
        RECT 1241.700 338.260 1241.840 338.680 ;
        RECT 1241.610 338.000 1241.930 338.260 ;
        RECT 1241.610 331.060 1241.930 331.120 ;
        RECT 1241.415 330.920 1241.930 331.060 ;
        RECT 1241.610 330.860 1241.930 330.920 ;
        RECT 1241.610 283.120 1241.930 283.180 ;
        RECT 1241.415 282.980 1241.930 283.120 ;
        RECT 1241.610 282.920 1241.930 282.980 ;
        RECT 1241.610 234.500 1241.930 234.560 ;
        RECT 1241.415 234.360 1241.930 234.500 ;
        RECT 1241.610 234.300 1241.930 234.360 ;
        RECT 1241.610 186.560 1241.930 186.620 ;
        RECT 1241.415 186.420 1241.930 186.560 ;
        RECT 1241.610 186.360 1241.930 186.420 ;
        RECT 1239.785 96.460 1240.075 96.505 ;
        RECT 1241.610 96.460 1241.930 96.520 ;
        RECT 1239.785 96.320 1241.930 96.460 ;
        RECT 1239.785 96.275 1240.075 96.320 ;
        RECT 1241.610 96.260 1241.930 96.320 ;
        RECT 1239.770 48.520 1240.090 48.580 ;
        RECT 1239.575 48.380 1240.090 48.520 ;
        RECT 1239.770 48.320 1240.090 48.380 ;
      LAYER via ;
        RECT 1241.640 1212.140 1241.900 1212.400 ;
        RECT 1386.540 1212.140 1386.800 1212.400 ;
        RECT 1240.720 1152.300 1240.980 1152.560 ;
        RECT 1241.180 1152.300 1241.440 1152.560 ;
        RECT 1239.800 1104.020 1240.060 1104.280 ;
        RECT 1241.640 1104.020 1241.900 1104.280 ;
        RECT 1240.720 1055.740 1240.980 1056.000 ;
        RECT 1241.180 1055.740 1241.440 1056.000 ;
        RECT 1240.720 1014.260 1240.980 1014.520 ;
        RECT 1241.640 1014.260 1241.900 1014.520 ;
        RECT 1241.640 1007.120 1241.900 1007.380 ;
        RECT 1240.720 959.180 1240.980 959.440 ;
        RECT 1240.720 917.700 1240.980 917.960 ;
        RECT 1241.640 917.700 1241.900 917.960 ;
        RECT 1240.720 910.560 1240.980 910.820 ;
        RECT 1241.640 910.560 1241.900 910.820 ;
        RECT 1241.640 814.000 1241.900 814.260 ;
        RECT 1241.640 766.060 1241.900 766.320 ;
        RECT 1241.640 717.440 1241.900 717.700 ;
        RECT 1241.640 669.500 1241.900 669.760 ;
        RECT 1241.640 620.540 1241.900 620.800 ;
        RECT 1241.640 572.600 1241.900 572.860 ;
        RECT 1241.640 523.980 1241.900 524.240 ;
        RECT 1241.640 476.040 1241.900 476.300 ;
        RECT 1241.640 427.420 1241.900 427.680 ;
        RECT 1241.640 379.480 1241.900 379.740 ;
        RECT 1241.640 338.680 1241.900 338.940 ;
        RECT 1241.640 338.000 1241.900 338.260 ;
        RECT 1241.640 330.860 1241.900 331.120 ;
        RECT 1241.640 282.920 1241.900 283.180 ;
        RECT 1241.640 234.300 1241.900 234.560 ;
        RECT 1241.640 186.360 1241.900 186.620 ;
        RECT 1241.640 96.260 1241.900 96.520 ;
        RECT 1239.800 48.320 1240.060 48.580 ;
      LAYER met2 ;
        RECT 1386.550 1219.680 1387.110 1228.680 ;
        RECT 1386.600 1212.430 1386.740 1219.680 ;
        RECT 1241.640 1212.110 1241.900 1212.430 ;
        RECT 1386.540 1212.110 1386.800 1212.430 ;
        RECT 1241.700 1200.610 1241.840 1212.110 ;
        RECT 1241.240 1200.470 1241.840 1200.610 ;
        RECT 1241.240 1152.590 1241.380 1200.470 ;
        RECT 1240.720 1152.445 1240.980 1152.590 ;
        RECT 1239.790 1152.075 1240.070 1152.445 ;
        RECT 1240.710 1152.075 1240.990 1152.445 ;
        RECT 1241.180 1152.270 1241.440 1152.590 ;
        RECT 1239.860 1104.310 1240.000 1152.075 ;
        RECT 1241.700 1104.310 1241.840 1104.465 ;
        RECT 1239.800 1103.990 1240.060 1104.310 ;
        RECT 1241.640 1104.050 1241.900 1104.310 ;
        RECT 1241.240 1103.990 1241.900 1104.050 ;
        RECT 1241.240 1103.910 1241.840 1103.990 ;
        RECT 1241.240 1056.030 1241.380 1103.910 ;
        RECT 1240.720 1055.710 1240.980 1056.030 ;
        RECT 1241.180 1055.710 1241.440 1056.030 ;
        RECT 1240.780 1014.550 1240.920 1055.710 ;
        RECT 1240.720 1014.230 1240.980 1014.550 ;
        RECT 1241.640 1014.230 1241.900 1014.550 ;
        RECT 1241.700 1007.410 1241.840 1014.230 ;
        RECT 1241.640 1007.090 1241.900 1007.410 ;
        RECT 1240.720 959.150 1240.980 959.470 ;
        RECT 1240.780 917.990 1240.920 959.150 ;
        RECT 1240.720 917.670 1240.980 917.990 ;
        RECT 1241.640 917.670 1241.900 917.990 ;
        RECT 1241.700 910.850 1241.840 917.670 ;
        RECT 1240.720 910.530 1240.980 910.850 ;
        RECT 1241.640 910.530 1241.900 910.850 ;
        RECT 1240.780 862.765 1240.920 910.530 ;
        RECT 1240.710 862.395 1240.990 862.765 ;
        RECT 1241.630 862.395 1241.910 862.765 ;
        RECT 1241.700 814.290 1241.840 862.395 ;
        RECT 1241.640 813.970 1241.900 814.290 ;
        RECT 1241.640 766.030 1241.900 766.350 ;
        RECT 1241.700 717.730 1241.840 766.030 ;
        RECT 1241.640 717.410 1241.900 717.730 ;
        RECT 1241.640 669.470 1241.900 669.790 ;
        RECT 1241.700 620.830 1241.840 669.470 ;
        RECT 1241.640 620.510 1241.900 620.830 ;
        RECT 1241.640 572.570 1241.900 572.890 ;
        RECT 1241.700 524.270 1241.840 572.570 ;
        RECT 1241.640 523.950 1241.900 524.270 ;
        RECT 1241.640 476.010 1241.900 476.330 ;
        RECT 1241.700 427.710 1241.840 476.010 ;
        RECT 1241.640 427.390 1241.900 427.710 ;
        RECT 1241.640 379.450 1241.900 379.770 ;
        RECT 1241.700 338.970 1241.840 379.450 ;
        RECT 1241.640 338.650 1241.900 338.970 ;
        RECT 1241.640 337.970 1241.900 338.290 ;
        RECT 1241.700 331.150 1241.840 337.970 ;
        RECT 1241.640 330.830 1241.900 331.150 ;
        RECT 1241.640 282.890 1241.900 283.210 ;
        RECT 1241.700 234.590 1241.840 282.890 ;
        RECT 1241.640 234.270 1241.900 234.590 ;
        RECT 1241.640 186.330 1241.900 186.650 ;
        RECT 1241.700 96.550 1241.840 186.330 ;
        RECT 1241.640 96.230 1241.900 96.550 ;
        RECT 1239.800 48.290 1240.060 48.610 ;
        RECT 1239.860 2.400 1240.000 48.290 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 1239.790 1152.120 1240.070 1152.400 ;
        RECT 1240.710 1152.120 1240.990 1152.400 ;
        RECT 1240.710 862.440 1240.990 862.720 ;
        RECT 1241.630 862.440 1241.910 862.720 ;
      LAYER met3 ;
        RECT 1239.765 1152.410 1240.095 1152.425 ;
        RECT 1240.685 1152.410 1241.015 1152.425 ;
        RECT 1239.765 1152.110 1241.015 1152.410 ;
        RECT 1239.765 1152.095 1240.095 1152.110 ;
        RECT 1240.685 1152.095 1241.015 1152.110 ;
        RECT 1240.685 862.730 1241.015 862.745 ;
        RECT 1241.605 862.730 1241.935 862.745 ;
        RECT 1240.685 862.430 1241.935 862.730 ;
        RECT 1240.685 862.415 1241.015 862.430 ;
        RECT 1241.605 862.415 1241.935 862.430 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 1210.980 1262.630 1211.040 ;
        RECT 1395.710 1210.980 1396.030 1211.040 ;
        RECT 1262.310 1210.840 1396.030 1210.980 ;
        RECT 1262.310 1210.780 1262.630 1210.840 ;
        RECT 1395.710 1210.780 1396.030 1210.840 ;
        RECT 1262.310 290.060 1262.630 290.320 ;
        RECT 1262.400 289.640 1262.540 290.060 ;
        RECT 1262.310 289.380 1262.630 289.640 ;
        RECT 1257.250 18.940 1257.570 19.000 ;
        RECT 1262.310 18.940 1262.630 19.000 ;
        RECT 1257.250 18.800 1262.630 18.940 ;
        RECT 1257.250 18.740 1257.570 18.800 ;
        RECT 1262.310 18.740 1262.630 18.800 ;
      LAYER via ;
        RECT 1262.340 1210.780 1262.600 1211.040 ;
        RECT 1395.740 1210.780 1396.000 1211.040 ;
        RECT 1262.340 290.060 1262.600 290.320 ;
        RECT 1262.340 289.380 1262.600 289.640 ;
        RECT 1257.280 18.740 1257.540 19.000 ;
        RECT 1262.340 18.740 1262.600 19.000 ;
      LAYER met2 ;
        RECT 1395.750 1219.680 1396.310 1228.680 ;
        RECT 1395.800 1211.070 1395.940 1219.680 ;
        RECT 1262.340 1210.750 1262.600 1211.070 ;
        RECT 1395.740 1210.750 1396.000 1211.070 ;
        RECT 1262.400 290.350 1262.540 1210.750 ;
        RECT 1262.340 290.030 1262.600 290.350 ;
        RECT 1262.340 289.350 1262.600 289.670 ;
        RECT 1262.400 19.030 1262.540 289.350 ;
        RECT 1257.280 18.710 1257.540 19.030 ;
        RECT 1262.340 18.710 1262.600 19.030 ;
        RECT 1257.340 2.400 1257.480 18.710 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 1212.000 1276.430 1212.060 ;
        RECT 1404.910 1212.000 1405.230 1212.060 ;
        RECT 1276.110 1211.860 1405.230 1212.000 ;
        RECT 1276.110 1211.800 1276.430 1211.860 ;
        RECT 1404.910 1211.800 1405.230 1211.860 ;
      LAYER via ;
        RECT 1276.140 1211.800 1276.400 1212.060 ;
        RECT 1404.940 1211.800 1405.200 1212.060 ;
      LAYER met2 ;
        RECT 1404.950 1219.680 1405.510 1228.680 ;
        RECT 1405.000 1212.090 1405.140 1219.680 ;
        RECT 1276.140 1211.770 1276.400 1212.090 ;
        RECT 1404.940 1211.770 1405.200 1212.090 ;
        RECT 1276.200 3.130 1276.340 1211.770 ;
        RECT 1275.280 2.990 1276.340 3.130 ;
        RECT 1275.280 2.400 1275.420 2.990 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 1213.360 1297.130 1213.420 ;
        RECT 1414.110 1213.360 1414.430 1213.420 ;
        RECT 1296.810 1213.220 1414.430 1213.360 ;
        RECT 1296.810 1213.160 1297.130 1213.220 ;
        RECT 1414.110 1213.160 1414.430 1213.220 ;
        RECT 1293.130 16.900 1293.450 16.960 ;
        RECT 1296.810 16.900 1297.130 16.960 ;
        RECT 1293.130 16.760 1297.130 16.900 ;
        RECT 1293.130 16.700 1293.450 16.760 ;
        RECT 1296.810 16.700 1297.130 16.760 ;
      LAYER via ;
        RECT 1296.840 1213.160 1297.100 1213.420 ;
        RECT 1414.140 1213.160 1414.400 1213.420 ;
        RECT 1293.160 16.700 1293.420 16.960 ;
        RECT 1296.840 16.700 1297.100 16.960 ;
      LAYER met2 ;
        RECT 1414.150 1219.680 1414.710 1228.680 ;
        RECT 1414.200 1213.450 1414.340 1219.680 ;
        RECT 1296.840 1213.130 1297.100 1213.450 ;
        RECT 1414.140 1213.130 1414.400 1213.450 ;
        RECT 1296.900 16.990 1297.040 1213.130 ;
        RECT 1293.160 16.670 1293.420 16.990 ;
        RECT 1296.840 16.670 1297.100 16.990 ;
        RECT 1293.220 2.400 1293.360 16.670 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1341.505 1207.425 1341.675 1213.035 ;
      LAYER mcon ;
        RECT 1341.505 1212.865 1341.675 1213.035 ;
      LAYER met1 ;
        RECT 1341.445 1213.020 1341.735 1213.065 ;
        RECT 1423.310 1213.020 1423.630 1213.080 ;
        RECT 1341.445 1212.880 1423.630 1213.020 ;
        RECT 1341.445 1212.835 1341.735 1212.880 ;
        RECT 1423.310 1212.820 1423.630 1212.880 ;
        RECT 1317.510 1207.580 1317.830 1207.640 ;
        RECT 1341.445 1207.580 1341.735 1207.625 ;
        RECT 1317.510 1207.440 1341.735 1207.580 ;
        RECT 1317.510 1207.380 1317.830 1207.440 ;
        RECT 1341.445 1207.395 1341.735 1207.440 ;
        RECT 1311.070 16.900 1311.390 16.960 ;
        RECT 1317.510 16.900 1317.830 16.960 ;
        RECT 1311.070 16.760 1317.830 16.900 ;
        RECT 1311.070 16.700 1311.390 16.760 ;
        RECT 1317.510 16.700 1317.830 16.760 ;
      LAYER via ;
        RECT 1423.340 1212.820 1423.600 1213.080 ;
        RECT 1317.540 1207.380 1317.800 1207.640 ;
        RECT 1311.100 16.700 1311.360 16.960 ;
        RECT 1317.540 16.700 1317.800 16.960 ;
      LAYER met2 ;
        RECT 1423.350 1219.680 1423.910 1228.680 ;
        RECT 1423.400 1213.110 1423.540 1219.680 ;
        RECT 1423.340 1212.790 1423.600 1213.110 ;
        RECT 1317.540 1207.350 1317.800 1207.670 ;
        RECT 1317.600 16.990 1317.740 1207.350 ;
        RECT 1311.100 16.670 1311.360 16.990 ;
        RECT 1317.540 16.670 1317.800 16.990 ;
        RECT 1311.160 2.400 1311.300 16.670 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1338.285 1212.865 1338.455 1214.055 ;
        RECT 1365.885 1213.885 1366.055 1214.735 ;
      LAYER mcon ;
        RECT 1365.885 1214.565 1366.055 1214.735 ;
        RECT 1338.285 1213.885 1338.455 1214.055 ;
      LAYER met1 ;
        RECT 1365.825 1214.720 1366.115 1214.765 ;
        RECT 1365.825 1214.580 1366.960 1214.720 ;
        RECT 1365.825 1214.535 1366.115 1214.580 ;
        RECT 1366.820 1214.380 1366.960 1214.580 ;
        RECT 1432.510 1214.380 1432.830 1214.440 ;
        RECT 1366.820 1214.240 1432.830 1214.380 ;
        RECT 1432.510 1214.180 1432.830 1214.240 ;
        RECT 1338.225 1214.040 1338.515 1214.085 ;
        RECT 1365.825 1214.040 1366.115 1214.085 ;
        RECT 1338.225 1213.900 1366.115 1214.040 ;
        RECT 1338.225 1213.855 1338.515 1213.900 ;
        RECT 1365.825 1213.855 1366.115 1213.900 ;
        RECT 1331.310 1213.020 1331.630 1213.080 ;
        RECT 1338.225 1213.020 1338.515 1213.065 ;
        RECT 1331.310 1212.880 1338.515 1213.020 ;
        RECT 1331.310 1212.820 1331.630 1212.880 ;
        RECT 1338.225 1212.835 1338.515 1212.880 ;
        RECT 1329.010 20.640 1329.330 20.700 ;
        RECT 1331.310 20.640 1331.630 20.700 ;
        RECT 1329.010 20.500 1331.630 20.640 ;
        RECT 1329.010 20.440 1329.330 20.500 ;
        RECT 1331.310 20.440 1331.630 20.500 ;
      LAYER via ;
        RECT 1432.540 1214.180 1432.800 1214.440 ;
        RECT 1331.340 1212.820 1331.600 1213.080 ;
        RECT 1329.040 20.440 1329.300 20.700 ;
        RECT 1331.340 20.440 1331.600 20.700 ;
      LAYER met2 ;
        RECT 1432.550 1219.680 1433.110 1228.680 ;
        RECT 1432.600 1214.470 1432.740 1219.680 ;
        RECT 1432.540 1214.150 1432.800 1214.470 ;
        RECT 1331.340 1212.790 1331.600 1213.110 ;
        RECT 1331.400 20.730 1331.540 1212.790 ;
        RECT 1329.040 20.410 1329.300 20.730 ;
        RECT 1331.340 20.410 1331.600 20.730 ;
        RECT 1329.100 2.400 1329.240 20.410 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1097.705 900.065 1097.875 917.575 ;
        RECT 1097.705 812.005 1097.875 855.355 ;
        RECT 1097.705 752.165 1097.875 800.275 ;
        RECT 1098.165 427.805 1098.335 475.915 ;
        RECT 1097.705 234.685 1097.875 331.075 ;
        RECT 1097.245 186.065 1097.415 227.715 ;
      LAYER mcon ;
        RECT 1097.705 917.405 1097.875 917.575 ;
        RECT 1097.705 855.185 1097.875 855.355 ;
        RECT 1097.705 800.105 1097.875 800.275 ;
        RECT 1098.165 475.745 1098.335 475.915 ;
        RECT 1097.705 330.905 1097.875 331.075 ;
        RECT 1097.245 227.545 1097.415 227.715 ;
      LAYER met1 ;
        RECT 1097.630 1055.400 1097.950 1055.660 ;
        RECT 1097.720 1055.260 1097.860 1055.400 ;
        RECT 1098.090 1055.260 1098.410 1055.320 ;
        RECT 1097.720 1055.120 1098.410 1055.260 ;
        RECT 1098.090 1055.060 1098.410 1055.120 ;
        RECT 1097.630 917.560 1097.950 917.620 ;
        RECT 1097.435 917.420 1097.950 917.560 ;
        RECT 1097.630 917.360 1097.950 917.420 ;
        RECT 1097.645 900.220 1097.935 900.265 ;
        RECT 1098.090 900.220 1098.410 900.280 ;
        RECT 1097.645 900.080 1098.410 900.220 ;
        RECT 1097.645 900.035 1097.935 900.080 ;
        RECT 1098.090 900.020 1098.410 900.080 ;
        RECT 1097.645 855.340 1097.935 855.385 ;
        RECT 1098.090 855.340 1098.410 855.400 ;
        RECT 1097.645 855.200 1098.410 855.340 ;
        RECT 1097.645 855.155 1097.935 855.200 ;
        RECT 1098.090 855.140 1098.410 855.200 ;
        RECT 1097.630 812.160 1097.950 812.220 ;
        RECT 1097.435 812.020 1097.950 812.160 ;
        RECT 1097.630 811.960 1097.950 812.020 ;
        RECT 1097.630 800.260 1097.950 800.320 ;
        RECT 1097.435 800.120 1097.950 800.260 ;
        RECT 1097.630 800.060 1097.950 800.120 ;
        RECT 1097.645 752.320 1097.935 752.365 ;
        RECT 1098.090 752.320 1098.410 752.380 ;
        RECT 1097.645 752.180 1098.410 752.320 ;
        RECT 1097.645 752.135 1097.935 752.180 ;
        RECT 1098.090 752.120 1098.410 752.180 ;
        RECT 1097.630 627.880 1097.950 627.940 ;
        RECT 1098.550 627.880 1098.870 627.940 ;
        RECT 1097.630 627.740 1098.870 627.880 ;
        RECT 1097.630 627.680 1097.950 627.740 ;
        RECT 1098.550 627.680 1098.870 627.740 ;
        RECT 1098.090 545.400 1098.410 545.660 ;
        RECT 1098.180 544.980 1098.320 545.400 ;
        RECT 1098.090 544.720 1098.410 544.980 ;
        RECT 1098.090 475.900 1098.410 475.960 ;
        RECT 1097.895 475.760 1098.410 475.900 ;
        RECT 1098.090 475.700 1098.410 475.760 ;
        RECT 1098.090 427.960 1098.410 428.020 ;
        RECT 1097.895 427.820 1098.410 427.960 ;
        RECT 1098.090 427.760 1098.410 427.820 ;
        RECT 1098.090 352.820 1098.410 352.880 ;
        RECT 1097.720 352.680 1098.410 352.820 ;
        RECT 1097.720 351.860 1097.860 352.680 ;
        RECT 1098.090 352.620 1098.410 352.680 ;
        RECT 1097.630 351.600 1097.950 351.860 ;
        RECT 1097.630 331.060 1097.950 331.120 ;
        RECT 1097.435 330.920 1097.950 331.060 ;
        RECT 1097.630 330.860 1097.950 330.920 ;
        RECT 1097.630 234.840 1097.950 234.900 ;
        RECT 1097.435 234.700 1097.950 234.840 ;
        RECT 1097.630 234.640 1097.950 234.700 ;
        RECT 1097.185 227.700 1097.475 227.745 ;
        RECT 1097.630 227.700 1097.950 227.760 ;
        RECT 1097.185 227.560 1097.950 227.700 ;
        RECT 1097.185 227.515 1097.475 227.560 ;
        RECT 1097.630 227.500 1097.950 227.560 ;
        RECT 1097.185 186.220 1097.475 186.265 ;
        RECT 1097.630 186.220 1097.950 186.280 ;
        RECT 1097.185 186.080 1097.950 186.220 ;
        RECT 1097.185 186.035 1097.475 186.080 ;
        RECT 1097.630 186.020 1097.950 186.080 ;
        RECT 1097.630 96.940 1097.950 97.200 ;
        RECT 1097.720 96.520 1097.860 96.940 ;
        RECT 1097.630 96.260 1097.950 96.520 ;
        RECT 686.390 35.940 686.710 36.000 ;
        RECT 1097.630 35.940 1097.950 36.000 ;
        RECT 686.390 35.800 1097.950 35.940 ;
        RECT 686.390 35.740 686.710 35.800 ;
        RECT 1097.630 35.740 1097.950 35.800 ;
      LAYER via ;
        RECT 1097.660 1055.400 1097.920 1055.660 ;
        RECT 1098.120 1055.060 1098.380 1055.320 ;
        RECT 1097.660 917.360 1097.920 917.620 ;
        RECT 1098.120 900.020 1098.380 900.280 ;
        RECT 1098.120 855.140 1098.380 855.400 ;
        RECT 1097.660 811.960 1097.920 812.220 ;
        RECT 1097.660 800.060 1097.920 800.320 ;
        RECT 1098.120 752.120 1098.380 752.380 ;
        RECT 1097.660 627.680 1097.920 627.940 ;
        RECT 1098.580 627.680 1098.840 627.940 ;
        RECT 1098.120 545.400 1098.380 545.660 ;
        RECT 1098.120 544.720 1098.380 544.980 ;
        RECT 1098.120 475.700 1098.380 475.960 ;
        RECT 1098.120 427.760 1098.380 428.020 ;
        RECT 1098.120 352.620 1098.380 352.880 ;
        RECT 1097.660 351.600 1097.920 351.860 ;
        RECT 1097.660 330.860 1097.920 331.120 ;
        RECT 1097.660 234.640 1097.920 234.900 ;
        RECT 1097.660 227.500 1097.920 227.760 ;
        RECT 1097.660 186.020 1097.920 186.280 ;
        RECT 1097.660 96.940 1097.920 97.200 ;
        RECT 1097.660 96.260 1097.920 96.520 ;
        RECT 686.420 35.740 686.680 36.000 ;
        RECT 1097.660 35.740 1097.920 36.000 ;
      LAYER met2 ;
        RECT 1102.270 1220.330 1102.830 1228.680 ;
        RECT 1100.940 1220.190 1102.830 1220.330 ;
        RECT 1100.940 1196.700 1101.080 1220.190 ;
        RECT 1102.270 1219.680 1102.830 1220.190 ;
        RECT 1097.720 1196.560 1101.080 1196.700 ;
        RECT 1097.720 1152.445 1097.860 1196.560 ;
        RECT 1097.650 1152.075 1097.930 1152.445 ;
        RECT 1098.570 1152.075 1098.850 1152.445 ;
        RECT 1098.640 1055.885 1098.780 1152.075 ;
        RECT 1097.650 1055.515 1097.930 1055.885 ;
        RECT 1098.570 1055.515 1098.850 1055.885 ;
        RECT 1097.660 1055.370 1097.920 1055.515 ;
        RECT 1098.120 1055.030 1098.380 1055.350 ;
        RECT 1098.180 942.210 1098.320 1055.030 ;
        RECT 1097.720 942.070 1098.320 942.210 ;
        RECT 1097.720 917.650 1097.860 942.070 ;
        RECT 1097.660 917.330 1097.920 917.650 ;
        RECT 1098.120 899.990 1098.380 900.310 ;
        RECT 1098.180 855.430 1098.320 899.990 ;
        RECT 1098.120 855.110 1098.380 855.430 ;
        RECT 1097.660 811.930 1097.920 812.250 ;
        RECT 1097.720 800.350 1097.860 811.930 ;
        RECT 1097.660 800.030 1097.920 800.350 ;
        RECT 1098.120 752.090 1098.380 752.410 ;
        RECT 1098.180 742.290 1098.320 752.090 ;
        RECT 1098.180 742.150 1098.780 742.290 ;
        RECT 1098.640 688.570 1098.780 742.150 ;
        RECT 1098.180 688.430 1098.780 688.570 ;
        RECT 1098.180 628.050 1098.320 688.430 ;
        RECT 1097.720 627.970 1098.320 628.050 ;
        RECT 1097.660 627.910 1098.320 627.970 ;
        RECT 1097.660 627.650 1097.920 627.910 ;
        RECT 1098.580 627.650 1098.840 627.970 ;
        RECT 1098.640 596.770 1098.780 627.650 ;
        RECT 1098.180 596.630 1098.780 596.770 ;
        RECT 1098.180 545.690 1098.320 596.630 ;
        RECT 1098.120 545.370 1098.380 545.690 ;
        RECT 1098.120 544.690 1098.380 545.010 ;
        RECT 1098.180 475.990 1098.320 544.690 ;
        RECT 1098.120 475.670 1098.380 475.990 ;
        RECT 1098.120 427.730 1098.380 428.050 ;
        RECT 1098.180 352.910 1098.320 427.730 ;
        RECT 1098.120 352.590 1098.380 352.910 ;
        RECT 1097.660 351.570 1097.920 351.890 ;
        RECT 1097.720 331.150 1097.860 351.570 ;
        RECT 1097.660 330.830 1097.920 331.150 ;
        RECT 1097.660 234.610 1097.920 234.930 ;
        RECT 1097.720 227.790 1097.860 234.610 ;
        RECT 1097.660 227.470 1097.920 227.790 ;
        RECT 1097.660 185.990 1097.920 186.310 ;
        RECT 1097.720 97.230 1097.860 185.990 ;
        RECT 1097.660 96.910 1097.920 97.230 ;
        RECT 1097.660 96.230 1097.920 96.550 ;
        RECT 1097.720 36.030 1097.860 96.230 ;
        RECT 686.420 35.710 686.680 36.030 ;
        RECT 1097.660 35.710 1097.920 36.030 ;
        RECT 686.480 2.400 686.620 35.710 ;
        RECT 686.270 -4.800 686.830 2.400 ;
      LAYER via2 ;
        RECT 1097.650 1152.120 1097.930 1152.400 ;
        RECT 1098.570 1152.120 1098.850 1152.400 ;
        RECT 1097.650 1055.560 1097.930 1055.840 ;
        RECT 1098.570 1055.560 1098.850 1055.840 ;
      LAYER met3 ;
        RECT 1097.625 1152.410 1097.955 1152.425 ;
        RECT 1098.545 1152.410 1098.875 1152.425 ;
        RECT 1097.625 1152.110 1098.875 1152.410 ;
        RECT 1097.625 1152.095 1097.955 1152.110 ;
        RECT 1098.545 1152.095 1098.875 1152.110 ;
        RECT 1097.625 1055.850 1097.955 1055.865 ;
        RECT 1098.545 1055.850 1098.875 1055.865 ;
        RECT 1097.625 1055.550 1098.875 1055.850 ;
        RECT 1097.625 1055.535 1097.955 1055.550 ;
        RECT 1098.545 1055.535 1098.875 1055.550 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.010 1208.600 1352.330 1208.660 ;
        RECT 1439.870 1208.600 1440.190 1208.660 ;
        RECT 1352.010 1208.460 1440.190 1208.600 ;
        RECT 1352.010 1208.400 1352.330 1208.460 ;
        RECT 1439.870 1208.400 1440.190 1208.460 ;
        RECT 1346.490 20.640 1346.810 20.700 ;
        RECT 1352.010 20.640 1352.330 20.700 ;
        RECT 1346.490 20.500 1352.330 20.640 ;
        RECT 1346.490 20.440 1346.810 20.500 ;
        RECT 1352.010 20.440 1352.330 20.500 ;
      LAYER via ;
        RECT 1352.040 1208.400 1352.300 1208.660 ;
        RECT 1439.900 1208.400 1440.160 1208.660 ;
        RECT 1346.520 20.440 1346.780 20.700 ;
        RECT 1352.040 20.440 1352.300 20.700 ;
      LAYER met2 ;
        RECT 1441.290 1220.330 1441.850 1228.680 ;
        RECT 1439.960 1220.190 1441.850 1220.330 ;
        RECT 1439.960 1208.690 1440.100 1220.190 ;
        RECT 1441.290 1219.680 1441.850 1220.190 ;
        RECT 1352.040 1208.370 1352.300 1208.690 ;
        RECT 1439.900 1208.370 1440.160 1208.690 ;
        RECT 1352.100 20.730 1352.240 1208.370 ;
        RECT 1346.520 20.410 1346.780 20.730 ;
        RECT 1352.040 20.410 1352.300 20.730 ;
        RECT 1346.580 2.400 1346.720 20.410 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 1208.940 1366.130 1209.000 ;
        RECT 1450.450 1208.940 1450.770 1209.000 ;
        RECT 1365.810 1208.800 1450.770 1208.940 ;
        RECT 1365.810 1208.740 1366.130 1208.800 ;
        RECT 1450.450 1208.740 1450.770 1208.800 ;
      LAYER via ;
        RECT 1365.840 1208.740 1366.100 1209.000 ;
        RECT 1450.480 1208.740 1450.740 1209.000 ;
      LAYER met2 ;
        RECT 1450.490 1219.680 1451.050 1228.680 ;
        RECT 1450.540 1209.030 1450.680 1219.680 ;
        RECT 1365.840 1208.710 1366.100 1209.030 ;
        RECT 1450.480 1208.710 1450.740 1209.030 ;
        RECT 1365.900 3.130 1366.040 1208.710 ;
        RECT 1364.520 2.990 1366.040 3.130 ;
        RECT 1364.520 2.400 1364.660 2.990 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.970 1212.340 1387.290 1212.400 ;
        RECT 1459.650 1212.340 1459.970 1212.400 ;
        RECT 1386.970 1212.200 1459.970 1212.340 ;
        RECT 1386.970 1212.140 1387.290 1212.200 ;
        RECT 1459.650 1212.140 1459.970 1212.200 ;
        RECT 1382.370 17.240 1382.690 17.300 ;
        RECT 1386.510 17.240 1386.830 17.300 ;
        RECT 1382.370 17.100 1386.830 17.240 ;
        RECT 1382.370 17.040 1382.690 17.100 ;
        RECT 1386.510 17.040 1386.830 17.100 ;
      LAYER via ;
        RECT 1387.000 1212.140 1387.260 1212.400 ;
        RECT 1459.680 1212.140 1459.940 1212.400 ;
        RECT 1382.400 17.040 1382.660 17.300 ;
        RECT 1386.540 17.040 1386.800 17.300 ;
      LAYER met2 ;
        RECT 1459.690 1219.680 1460.250 1228.680 ;
        RECT 1459.740 1212.430 1459.880 1219.680 ;
        RECT 1387.000 1212.110 1387.260 1212.430 ;
        RECT 1459.680 1212.110 1459.940 1212.430 ;
        RECT 1387.060 1211.490 1387.200 1212.110 ;
        RECT 1386.600 1211.350 1387.200 1211.490 ;
        RECT 1386.600 17.330 1386.740 1211.350 ;
        RECT 1382.400 17.010 1382.660 17.330 ;
        RECT 1386.540 17.010 1386.800 17.330 ;
        RECT 1382.460 2.400 1382.600 17.010 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 1210.980 1400.630 1211.040 ;
        RECT 1468.850 1210.980 1469.170 1211.040 ;
        RECT 1400.310 1210.840 1469.170 1210.980 ;
        RECT 1400.310 1210.780 1400.630 1210.840 ;
        RECT 1468.850 1210.780 1469.170 1210.840 ;
      LAYER via ;
        RECT 1400.340 1210.780 1400.600 1211.040 ;
        RECT 1468.880 1210.780 1469.140 1211.040 ;
      LAYER met2 ;
        RECT 1468.890 1219.680 1469.450 1228.680 ;
        RECT 1468.940 1211.070 1469.080 1219.680 ;
        RECT 1400.340 1210.750 1400.600 1211.070 ;
        RECT 1468.880 1210.750 1469.140 1211.070 ;
        RECT 1400.400 2.400 1400.540 1210.750 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1211.660 1421.330 1211.720 ;
        RECT 1478.050 1211.660 1478.370 1211.720 ;
        RECT 1421.010 1211.520 1478.370 1211.660 ;
        RECT 1421.010 1211.460 1421.330 1211.520 ;
        RECT 1478.050 1211.460 1478.370 1211.520 ;
        RECT 1418.250 14.860 1418.570 14.920 ;
        RECT 1421.010 14.860 1421.330 14.920 ;
        RECT 1418.250 14.720 1421.330 14.860 ;
        RECT 1418.250 14.660 1418.570 14.720 ;
        RECT 1421.010 14.660 1421.330 14.720 ;
      LAYER via ;
        RECT 1421.040 1211.460 1421.300 1211.720 ;
        RECT 1478.080 1211.460 1478.340 1211.720 ;
        RECT 1418.280 14.660 1418.540 14.920 ;
        RECT 1421.040 14.660 1421.300 14.920 ;
      LAYER met2 ;
        RECT 1478.090 1219.680 1478.650 1228.680 ;
        RECT 1478.140 1211.750 1478.280 1219.680 ;
        RECT 1421.040 1211.430 1421.300 1211.750 ;
        RECT 1478.080 1211.430 1478.340 1211.750 ;
        RECT 1421.100 14.950 1421.240 1211.430 ;
        RECT 1418.280 14.630 1418.540 14.950 ;
        RECT 1421.040 14.630 1421.300 14.950 ;
        RECT 1418.340 2.400 1418.480 14.630 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1441.250 1212.680 1441.570 1212.740 ;
        RECT 1487.250 1212.680 1487.570 1212.740 ;
        RECT 1441.250 1212.540 1487.570 1212.680 ;
        RECT 1441.250 1212.480 1441.570 1212.540 ;
        RECT 1487.250 1212.480 1487.570 1212.540 ;
        RECT 1435.730 15.200 1436.050 15.260 ;
        RECT 1441.250 15.200 1441.570 15.260 ;
        RECT 1435.730 15.060 1441.570 15.200 ;
        RECT 1435.730 15.000 1436.050 15.060 ;
        RECT 1441.250 15.000 1441.570 15.060 ;
      LAYER via ;
        RECT 1441.280 1212.480 1441.540 1212.740 ;
        RECT 1487.280 1212.480 1487.540 1212.740 ;
        RECT 1435.760 15.000 1436.020 15.260 ;
        RECT 1441.280 15.000 1441.540 15.260 ;
      LAYER met2 ;
        RECT 1487.290 1219.680 1487.850 1228.680 ;
        RECT 1487.340 1212.770 1487.480 1219.680 ;
        RECT 1441.280 1212.450 1441.540 1212.770 ;
        RECT 1487.280 1212.450 1487.540 1212.770 ;
        RECT 1441.340 15.290 1441.480 1212.450 ;
        RECT 1435.760 14.970 1436.020 15.290 ;
        RECT 1441.280 14.970 1441.540 15.290 ;
        RECT 1435.820 2.400 1435.960 14.970 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1453.745 2.805 1453.915 14.195 ;
      LAYER mcon ;
        RECT 1453.745 14.025 1453.915 14.195 ;
      LAYER met1 ;
        RECT 1455.510 1208.940 1455.830 1209.000 ;
        RECT 1496.450 1208.940 1496.770 1209.000 ;
        RECT 1455.510 1208.800 1496.770 1208.940 ;
        RECT 1455.510 1208.740 1455.830 1208.800 ;
        RECT 1496.450 1208.740 1496.770 1208.800 ;
        RECT 1453.685 14.180 1453.975 14.225 ;
        RECT 1455.510 14.180 1455.830 14.240 ;
        RECT 1453.685 14.040 1455.830 14.180 ;
        RECT 1453.685 13.995 1453.975 14.040 ;
        RECT 1455.510 13.980 1455.830 14.040 ;
        RECT 1453.670 2.960 1453.990 3.020 ;
        RECT 1453.475 2.820 1453.990 2.960 ;
        RECT 1453.670 2.760 1453.990 2.820 ;
      LAYER via ;
        RECT 1455.540 1208.740 1455.800 1209.000 ;
        RECT 1496.480 1208.740 1496.740 1209.000 ;
        RECT 1455.540 13.980 1455.800 14.240 ;
        RECT 1453.700 2.760 1453.960 3.020 ;
      LAYER met2 ;
        RECT 1496.490 1219.680 1497.050 1228.680 ;
        RECT 1496.540 1209.030 1496.680 1219.680 ;
        RECT 1455.540 1208.710 1455.800 1209.030 ;
        RECT 1496.480 1208.710 1496.740 1209.030 ;
        RECT 1455.600 14.270 1455.740 1208.710 ;
        RECT 1455.540 13.950 1455.800 14.270 ;
        RECT 1453.700 2.730 1453.960 3.050 ;
        RECT 1453.760 2.400 1453.900 2.730 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1487.250 1207.920 1487.570 1207.980 ;
        RECT 1505.650 1207.920 1505.970 1207.980 ;
        RECT 1487.250 1207.780 1505.970 1207.920 ;
        RECT 1487.250 1207.720 1487.570 1207.780 ;
        RECT 1505.650 1207.720 1505.970 1207.780 ;
        RECT 1471.610 16.900 1471.930 16.960 ;
        RECT 1487.250 16.900 1487.570 16.960 ;
        RECT 1471.610 16.760 1487.570 16.900 ;
        RECT 1471.610 16.700 1471.930 16.760 ;
        RECT 1487.250 16.700 1487.570 16.760 ;
      LAYER via ;
        RECT 1487.280 1207.720 1487.540 1207.980 ;
        RECT 1505.680 1207.720 1505.940 1207.980 ;
        RECT 1471.640 16.700 1471.900 16.960 ;
        RECT 1487.280 16.700 1487.540 16.960 ;
      LAYER met2 ;
        RECT 1505.690 1219.680 1506.250 1228.680 ;
        RECT 1505.740 1208.010 1505.880 1219.680 ;
        RECT 1487.280 1207.690 1487.540 1208.010 ;
        RECT 1505.680 1207.690 1505.940 1208.010 ;
        RECT 1487.340 16.990 1487.480 1207.690 ;
        RECT 1471.640 16.670 1471.900 16.990 ;
        RECT 1487.280 16.670 1487.540 16.990 ;
        RECT 1471.700 2.400 1471.840 16.670 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.950 1207.580 1508.270 1207.640 ;
        RECT 1514.850 1207.580 1515.170 1207.640 ;
        RECT 1507.950 1207.440 1515.170 1207.580 ;
        RECT 1507.950 1207.380 1508.270 1207.440 ;
        RECT 1514.850 1207.380 1515.170 1207.440 ;
        RECT 1489.550 17.240 1489.870 17.300 ;
        RECT 1507.950 17.240 1508.270 17.300 ;
        RECT 1489.550 17.100 1508.270 17.240 ;
        RECT 1489.550 17.040 1489.870 17.100 ;
        RECT 1507.950 17.040 1508.270 17.100 ;
      LAYER via ;
        RECT 1507.980 1207.380 1508.240 1207.640 ;
        RECT 1514.880 1207.380 1515.140 1207.640 ;
        RECT 1489.580 17.040 1489.840 17.300 ;
        RECT 1507.980 17.040 1508.240 17.300 ;
      LAYER met2 ;
        RECT 1514.890 1219.680 1515.450 1228.680 ;
        RECT 1514.940 1207.670 1515.080 1219.680 ;
        RECT 1507.980 1207.350 1508.240 1207.670 ;
        RECT 1514.880 1207.350 1515.140 1207.670 ;
        RECT 1508.040 17.330 1508.180 1207.350 ;
        RECT 1489.580 17.010 1489.840 17.330 ;
        RECT 1507.980 17.010 1508.240 17.330 ;
        RECT 1489.640 2.400 1489.780 17.010 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1514.390 1208.260 1514.710 1208.320 ;
        RECT 1524.050 1208.260 1524.370 1208.320 ;
        RECT 1514.390 1208.120 1524.370 1208.260 ;
        RECT 1514.390 1208.060 1514.710 1208.120 ;
        RECT 1524.050 1208.060 1524.370 1208.120 ;
        RECT 1507.030 17.580 1507.350 17.640 ;
        RECT 1514.390 17.580 1514.710 17.640 ;
        RECT 1507.030 17.440 1514.710 17.580 ;
        RECT 1507.030 17.380 1507.350 17.440 ;
        RECT 1514.390 17.380 1514.710 17.440 ;
      LAYER via ;
        RECT 1514.420 1208.060 1514.680 1208.320 ;
        RECT 1524.080 1208.060 1524.340 1208.320 ;
        RECT 1507.060 17.380 1507.320 17.640 ;
        RECT 1514.420 17.380 1514.680 17.640 ;
      LAYER met2 ;
        RECT 1524.090 1219.680 1524.650 1228.680 ;
        RECT 1524.140 1208.350 1524.280 1219.680 ;
        RECT 1514.420 1208.030 1514.680 1208.350 ;
        RECT 1524.080 1208.030 1524.340 1208.350 ;
        RECT 1514.480 17.670 1514.620 1208.030 ;
        RECT 1507.060 17.350 1507.320 17.670 ;
        RECT 1514.420 17.350 1514.680 17.670 ;
        RECT 1507.120 2.400 1507.260 17.350 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 35.600 704.650 35.660 ;
        RECT 1111.430 35.600 1111.750 35.660 ;
        RECT 704.330 35.460 1111.750 35.600 ;
        RECT 704.330 35.400 704.650 35.460 ;
        RECT 1111.430 35.400 1111.750 35.460 ;
      LAYER via ;
        RECT 704.360 35.400 704.620 35.660 ;
        RECT 1111.460 35.400 1111.720 35.660 ;
      LAYER met2 ;
        RECT 1111.470 1219.680 1112.030 1228.680 ;
        RECT 1111.520 35.690 1111.660 1219.680 ;
        RECT 704.360 35.370 704.620 35.690 ;
        RECT 1111.460 35.370 1111.720 35.690 ;
        RECT 704.420 2.400 704.560 35.370 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.970 20.640 1525.290 20.700 ;
        RECT 1530.950 20.640 1531.270 20.700 ;
        RECT 1524.970 20.500 1531.270 20.640 ;
        RECT 1524.970 20.440 1525.290 20.500 ;
        RECT 1530.950 20.440 1531.270 20.500 ;
      LAYER via ;
        RECT 1525.000 20.440 1525.260 20.700 ;
        RECT 1530.980 20.440 1531.240 20.700 ;
      LAYER met2 ;
        RECT 1533.290 1220.330 1533.850 1228.680 ;
        RECT 1531.960 1220.190 1533.850 1220.330 ;
        RECT 1531.960 1207.920 1532.100 1220.190 ;
        RECT 1533.290 1219.680 1533.850 1220.190 ;
        RECT 1531.040 1207.780 1532.100 1207.920 ;
        RECT 1531.040 20.730 1531.180 1207.780 ;
        RECT 1525.000 20.410 1525.260 20.730 ;
        RECT 1530.980 20.410 1531.240 20.730 ;
        RECT 1525.060 2.400 1525.200 20.410 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1539.765 786.505 1539.935 821.015 ;
        RECT 1539.765 689.605 1539.935 724.455 ;
        RECT 1539.765 593.045 1539.935 627.895 ;
        RECT 1539.765 496.485 1539.935 531.335 ;
        RECT 1539.765 386.325 1539.935 434.775 ;
        RECT 1539.305 241.485 1539.475 289.595 ;
        RECT 1539.765 144.925 1539.935 193.035 ;
      LAYER mcon ;
        RECT 1539.765 820.845 1539.935 821.015 ;
        RECT 1539.765 724.285 1539.935 724.455 ;
        RECT 1539.765 627.725 1539.935 627.895 ;
        RECT 1539.765 531.165 1539.935 531.335 ;
        RECT 1539.765 434.605 1539.935 434.775 ;
        RECT 1539.305 289.425 1539.475 289.595 ;
        RECT 1539.765 192.865 1539.935 193.035 ;
      LAYER met1 ;
        RECT 1539.230 1124.960 1539.550 1125.020 ;
        RECT 1540.150 1124.960 1540.470 1125.020 ;
        RECT 1539.230 1124.820 1540.470 1124.960 ;
        RECT 1539.230 1124.760 1539.550 1124.820 ;
        RECT 1540.150 1124.760 1540.470 1124.820 ;
        RECT 1539.230 1028.400 1539.550 1028.460 ;
        RECT 1540.150 1028.400 1540.470 1028.460 ;
        RECT 1539.230 1028.260 1540.470 1028.400 ;
        RECT 1539.230 1028.200 1539.550 1028.260 ;
        RECT 1540.150 1028.200 1540.470 1028.260 ;
        RECT 1539.230 931.840 1539.550 931.900 ;
        RECT 1540.150 931.840 1540.470 931.900 ;
        RECT 1539.230 931.700 1540.470 931.840 ;
        RECT 1539.230 931.640 1539.550 931.700 ;
        RECT 1540.150 931.640 1540.470 931.700 ;
        RECT 1540.150 869.620 1540.470 869.680 ;
        RECT 1541.070 869.620 1541.390 869.680 ;
        RECT 1540.150 869.480 1541.390 869.620 ;
        RECT 1540.150 869.420 1540.470 869.480 ;
        RECT 1541.070 869.420 1541.390 869.480 ;
        RECT 1539.230 835.280 1539.550 835.340 ;
        RECT 1540.150 835.280 1540.470 835.340 ;
        RECT 1539.230 835.140 1540.470 835.280 ;
        RECT 1539.230 835.080 1539.550 835.140 ;
        RECT 1540.150 835.080 1540.470 835.140 ;
        RECT 1539.690 821.000 1540.010 821.060 ;
        RECT 1539.495 820.860 1540.010 821.000 ;
        RECT 1539.690 820.800 1540.010 820.860 ;
        RECT 1539.690 786.660 1540.010 786.720 ;
        RECT 1539.495 786.520 1540.010 786.660 ;
        RECT 1539.690 786.460 1540.010 786.520 ;
        RECT 1539.230 738.380 1539.550 738.440 ;
        RECT 1540.150 738.380 1540.470 738.440 ;
        RECT 1539.230 738.240 1540.470 738.380 ;
        RECT 1539.230 738.180 1539.550 738.240 ;
        RECT 1540.150 738.180 1540.470 738.240 ;
        RECT 1539.690 724.440 1540.010 724.500 ;
        RECT 1539.495 724.300 1540.010 724.440 ;
        RECT 1539.690 724.240 1540.010 724.300 ;
        RECT 1539.690 689.760 1540.010 689.820 ;
        RECT 1539.495 689.620 1540.010 689.760 ;
        RECT 1539.690 689.560 1540.010 689.620 ;
        RECT 1539.230 641.820 1539.550 641.880 ;
        RECT 1540.150 641.820 1540.470 641.880 ;
        RECT 1539.230 641.680 1540.470 641.820 ;
        RECT 1539.230 641.620 1539.550 641.680 ;
        RECT 1540.150 641.620 1540.470 641.680 ;
        RECT 1539.690 627.880 1540.010 627.940 ;
        RECT 1539.495 627.740 1540.010 627.880 ;
        RECT 1539.690 627.680 1540.010 627.740 ;
        RECT 1539.690 593.200 1540.010 593.260 ;
        RECT 1539.495 593.060 1540.010 593.200 ;
        RECT 1539.690 593.000 1540.010 593.060 ;
        RECT 1539.230 545.260 1539.550 545.320 ;
        RECT 1540.150 545.260 1540.470 545.320 ;
        RECT 1539.230 545.120 1540.470 545.260 ;
        RECT 1539.230 545.060 1539.550 545.120 ;
        RECT 1540.150 545.060 1540.470 545.120 ;
        RECT 1539.690 531.320 1540.010 531.380 ;
        RECT 1539.495 531.180 1540.010 531.320 ;
        RECT 1539.690 531.120 1540.010 531.180 ;
        RECT 1539.690 496.640 1540.010 496.700 ;
        RECT 1539.495 496.500 1540.010 496.640 ;
        RECT 1539.690 496.440 1540.010 496.500 ;
        RECT 1539.230 448.700 1539.550 448.760 ;
        RECT 1540.150 448.700 1540.470 448.760 ;
        RECT 1539.230 448.560 1540.470 448.700 ;
        RECT 1539.230 448.500 1539.550 448.560 ;
        RECT 1540.150 448.500 1540.470 448.560 ;
        RECT 1539.690 434.760 1540.010 434.820 ;
        RECT 1539.495 434.620 1540.010 434.760 ;
        RECT 1539.690 434.560 1540.010 434.620 ;
        RECT 1539.705 386.480 1539.995 386.525 ;
        RECT 1540.150 386.480 1540.470 386.540 ;
        RECT 1539.705 386.340 1540.470 386.480 ;
        RECT 1539.705 386.295 1539.995 386.340 ;
        RECT 1540.150 386.280 1540.470 386.340 ;
        RECT 1539.690 338.540 1540.010 338.600 ;
        RECT 1540.150 338.540 1540.470 338.600 ;
        RECT 1539.690 338.400 1540.470 338.540 ;
        RECT 1539.690 338.340 1540.010 338.400 ;
        RECT 1540.150 338.340 1540.470 338.400 ;
        RECT 1538.310 337.860 1538.630 337.920 ;
        RECT 1539.690 337.860 1540.010 337.920 ;
        RECT 1538.310 337.720 1540.010 337.860 ;
        RECT 1538.310 337.660 1538.630 337.720 ;
        RECT 1539.690 337.660 1540.010 337.720 ;
        RECT 1539.230 289.580 1539.550 289.640 ;
        RECT 1539.035 289.440 1539.550 289.580 ;
        RECT 1539.230 289.380 1539.550 289.440 ;
        RECT 1539.245 241.640 1539.535 241.685 ;
        RECT 1539.690 241.640 1540.010 241.700 ;
        RECT 1539.245 241.500 1540.010 241.640 ;
        RECT 1539.245 241.455 1539.535 241.500 ;
        RECT 1539.690 241.440 1540.010 241.500 ;
        RECT 1539.705 193.020 1539.995 193.065 ;
        RECT 1540.150 193.020 1540.470 193.080 ;
        RECT 1539.705 192.880 1540.470 193.020 ;
        RECT 1539.705 192.835 1539.995 192.880 ;
        RECT 1540.150 192.820 1540.470 192.880 ;
        RECT 1539.690 145.080 1540.010 145.140 ;
        RECT 1539.495 144.940 1540.010 145.080 ;
        RECT 1539.690 144.880 1540.010 144.940 ;
        RECT 1540.150 20.640 1540.470 20.700 ;
        RECT 1542.910 20.640 1543.230 20.700 ;
        RECT 1540.150 20.500 1543.230 20.640 ;
        RECT 1540.150 20.440 1540.470 20.500 ;
        RECT 1542.910 20.440 1543.230 20.500 ;
      LAYER via ;
        RECT 1539.260 1124.760 1539.520 1125.020 ;
        RECT 1540.180 1124.760 1540.440 1125.020 ;
        RECT 1539.260 1028.200 1539.520 1028.460 ;
        RECT 1540.180 1028.200 1540.440 1028.460 ;
        RECT 1539.260 931.640 1539.520 931.900 ;
        RECT 1540.180 931.640 1540.440 931.900 ;
        RECT 1540.180 869.420 1540.440 869.680 ;
        RECT 1541.100 869.420 1541.360 869.680 ;
        RECT 1539.260 835.080 1539.520 835.340 ;
        RECT 1540.180 835.080 1540.440 835.340 ;
        RECT 1539.720 820.800 1539.980 821.060 ;
        RECT 1539.720 786.460 1539.980 786.720 ;
        RECT 1539.260 738.180 1539.520 738.440 ;
        RECT 1540.180 738.180 1540.440 738.440 ;
        RECT 1539.720 724.240 1539.980 724.500 ;
        RECT 1539.720 689.560 1539.980 689.820 ;
        RECT 1539.260 641.620 1539.520 641.880 ;
        RECT 1540.180 641.620 1540.440 641.880 ;
        RECT 1539.720 627.680 1539.980 627.940 ;
        RECT 1539.720 593.000 1539.980 593.260 ;
        RECT 1539.260 545.060 1539.520 545.320 ;
        RECT 1540.180 545.060 1540.440 545.320 ;
        RECT 1539.720 531.120 1539.980 531.380 ;
        RECT 1539.720 496.440 1539.980 496.700 ;
        RECT 1539.260 448.500 1539.520 448.760 ;
        RECT 1540.180 448.500 1540.440 448.760 ;
        RECT 1539.720 434.560 1539.980 434.820 ;
        RECT 1540.180 386.280 1540.440 386.540 ;
        RECT 1539.720 338.340 1539.980 338.600 ;
        RECT 1540.180 338.340 1540.440 338.600 ;
        RECT 1538.340 337.660 1538.600 337.920 ;
        RECT 1539.720 337.660 1539.980 337.920 ;
        RECT 1539.260 289.380 1539.520 289.640 ;
        RECT 1539.720 241.440 1539.980 241.700 ;
        RECT 1540.180 192.820 1540.440 193.080 ;
        RECT 1539.720 144.880 1539.980 145.140 ;
        RECT 1540.180 20.440 1540.440 20.700 ;
        RECT 1542.940 20.440 1543.200 20.700 ;
      LAYER met2 ;
        RECT 1542.490 1220.330 1543.050 1228.680 ;
        RECT 1540.240 1220.190 1543.050 1220.330 ;
        RECT 1540.240 1125.050 1540.380 1220.190 ;
        RECT 1542.490 1219.680 1543.050 1220.190 ;
        RECT 1539.260 1124.730 1539.520 1125.050 ;
        RECT 1540.180 1124.730 1540.440 1125.050 ;
        RECT 1539.320 1124.450 1539.460 1124.730 ;
        RECT 1539.320 1124.310 1539.920 1124.450 ;
        RECT 1539.780 1076.850 1539.920 1124.310 ;
        RECT 1539.780 1076.710 1540.380 1076.850 ;
        RECT 1540.240 1028.490 1540.380 1076.710 ;
        RECT 1539.260 1028.170 1539.520 1028.490 ;
        RECT 1540.180 1028.170 1540.440 1028.490 ;
        RECT 1539.320 1027.890 1539.460 1028.170 ;
        RECT 1539.320 1027.750 1539.920 1027.890 ;
        RECT 1539.780 980.290 1539.920 1027.750 ;
        RECT 1539.780 980.150 1540.380 980.290 ;
        RECT 1540.240 931.930 1540.380 980.150 ;
        RECT 1539.260 931.610 1539.520 931.930 ;
        RECT 1540.180 931.610 1540.440 931.930 ;
        RECT 1539.320 931.330 1539.460 931.610 ;
        RECT 1539.320 931.190 1539.920 931.330 ;
        RECT 1539.780 917.845 1539.920 931.190 ;
        RECT 1539.710 917.475 1539.990 917.845 ;
        RECT 1541.090 917.475 1541.370 917.845 ;
        RECT 1541.160 869.710 1541.300 917.475 ;
        RECT 1540.180 869.390 1540.440 869.710 ;
        RECT 1541.100 869.390 1541.360 869.710 ;
        RECT 1540.240 835.370 1540.380 869.390 ;
        RECT 1539.260 835.050 1539.520 835.370 ;
        RECT 1540.180 835.050 1540.440 835.370 ;
        RECT 1539.320 834.770 1539.460 835.050 ;
        RECT 1539.320 834.630 1539.920 834.770 ;
        RECT 1539.780 821.090 1539.920 834.630 ;
        RECT 1539.720 820.770 1539.980 821.090 ;
        RECT 1539.720 786.430 1539.980 786.750 ;
        RECT 1539.780 772.890 1539.920 786.430 ;
        RECT 1539.780 772.750 1540.380 772.890 ;
        RECT 1540.240 738.470 1540.380 772.750 ;
        RECT 1539.260 738.210 1539.520 738.470 ;
        RECT 1539.260 738.150 1539.920 738.210 ;
        RECT 1540.180 738.150 1540.440 738.470 ;
        RECT 1539.320 738.070 1539.920 738.150 ;
        RECT 1539.780 724.530 1539.920 738.070 ;
        RECT 1539.720 724.210 1539.980 724.530 ;
        RECT 1539.720 689.530 1539.980 689.850 ;
        RECT 1539.780 676.330 1539.920 689.530 ;
        RECT 1539.780 676.190 1540.380 676.330 ;
        RECT 1540.240 641.910 1540.380 676.190 ;
        RECT 1539.260 641.650 1539.520 641.910 ;
        RECT 1539.260 641.590 1539.920 641.650 ;
        RECT 1540.180 641.590 1540.440 641.910 ;
        RECT 1539.320 641.510 1539.920 641.590 ;
        RECT 1539.780 627.970 1539.920 641.510 ;
        RECT 1539.720 627.650 1539.980 627.970 ;
        RECT 1539.720 592.970 1539.980 593.290 ;
        RECT 1539.780 579.770 1539.920 592.970 ;
        RECT 1539.780 579.630 1540.380 579.770 ;
        RECT 1540.240 545.350 1540.380 579.630 ;
        RECT 1539.260 545.090 1539.520 545.350 ;
        RECT 1539.260 545.030 1539.920 545.090 ;
        RECT 1540.180 545.030 1540.440 545.350 ;
        RECT 1539.320 544.950 1539.920 545.030 ;
        RECT 1539.780 531.410 1539.920 544.950 ;
        RECT 1539.720 531.090 1539.980 531.410 ;
        RECT 1539.720 496.410 1539.980 496.730 ;
        RECT 1539.780 483.210 1539.920 496.410 ;
        RECT 1539.780 483.070 1540.380 483.210 ;
        RECT 1540.240 448.790 1540.380 483.070 ;
        RECT 1539.260 448.530 1539.520 448.790 ;
        RECT 1539.260 448.470 1539.920 448.530 ;
        RECT 1540.180 448.470 1540.440 448.790 ;
        RECT 1539.320 448.390 1539.920 448.470 ;
        RECT 1539.780 434.850 1539.920 448.390 ;
        RECT 1539.720 434.530 1539.980 434.850 ;
        RECT 1540.180 386.250 1540.440 386.570 ;
        RECT 1540.240 338.630 1540.380 386.250 ;
        RECT 1539.720 338.310 1539.980 338.630 ;
        RECT 1540.180 338.310 1540.440 338.630 ;
        RECT 1539.780 337.950 1539.920 338.310 ;
        RECT 1538.340 337.630 1538.600 337.950 ;
        RECT 1539.720 337.630 1539.980 337.950 ;
        RECT 1538.400 290.205 1538.540 337.630 ;
        RECT 1538.330 289.835 1538.610 290.205 ;
        RECT 1539.250 289.835 1539.530 290.205 ;
        RECT 1539.320 289.670 1539.460 289.835 ;
        RECT 1539.260 289.350 1539.520 289.670 ;
        RECT 1539.720 241.410 1539.980 241.730 ;
        RECT 1539.780 241.245 1539.920 241.410 ;
        RECT 1539.710 240.875 1539.990 241.245 ;
        RECT 1540.170 193.275 1540.450 193.645 ;
        RECT 1540.240 193.110 1540.380 193.275 ;
        RECT 1540.180 192.790 1540.440 193.110 ;
        RECT 1539.720 144.850 1539.980 145.170 ;
        RECT 1539.780 144.570 1539.920 144.850 ;
        RECT 1539.780 144.430 1540.380 144.570 ;
        RECT 1540.240 109.890 1540.380 144.430 ;
        RECT 1539.780 109.750 1540.380 109.890 ;
        RECT 1539.780 62.290 1539.920 109.750 ;
        RECT 1539.780 62.150 1540.380 62.290 ;
        RECT 1540.240 20.730 1540.380 62.150 ;
        RECT 1540.180 20.410 1540.440 20.730 ;
        RECT 1542.940 20.410 1543.200 20.730 ;
        RECT 1543.000 2.400 1543.140 20.410 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 1539.710 917.520 1539.990 917.800 ;
        RECT 1541.090 917.520 1541.370 917.800 ;
        RECT 1538.330 289.880 1538.610 290.160 ;
        RECT 1539.250 289.880 1539.530 290.160 ;
        RECT 1539.710 240.920 1539.990 241.200 ;
        RECT 1540.170 193.320 1540.450 193.600 ;
      LAYER met3 ;
        RECT 1539.685 917.810 1540.015 917.825 ;
        RECT 1541.065 917.810 1541.395 917.825 ;
        RECT 1539.685 917.510 1541.395 917.810 ;
        RECT 1539.685 917.495 1540.015 917.510 ;
        RECT 1541.065 917.495 1541.395 917.510 ;
        RECT 1538.305 290.170 1538.635 290.185 ;
        RECT 1539.225 290.170 1539.555 290.185 ;
        RECT 1538.305 289.870 1539.555 290.170 ;
        RECT 1538.305 289.855 1538.635 289.870 ;
        RECT 1539.225 289.855 1539.555 289.870 ;
        RECT 1539.685 241.220 1540.015 241.225 ;
        RECT 1539.430 241.210 1540.015 241.220 ;
        RECT 1539.430 240.910 1540.240 241.210 ;
        RECT 1539.430 240.900 1540.015 240.910 ;
        RECT 1539.685 240.895 1540.015 240.900 ;
        RECT 1539.430 193.610 1539.810 193.620 ;
        RECT 1540.145 193.610 1540.475 193.625 ;
        RECT 1539.430 193.310 1540.475 193.610 ;
        RECT 1539.430 193.300 1539.810 193.310 ;
        RECT 1540.145 193.295 1540.475 193.310 ;
      LAYER via3 ;
        RECT 1539.460 240.900 1539.780 241.220 ;
        RECT 1539.460 193.300 1539.780 193.620 ;
      LAYER met4 ;
        RECT 1539.455 240.895 1539.785 241.225 ;
        RECT 1539.470 193.625 1539.770 240.895 ;
        RECT 1539.455 193.295 1539.785 193.625 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1551.650 1207.920 1551.970 1207.980 ;
        RECT 1559.470 1207.920 1559.790 1207.980 ;
        RECT 1551.650 1207.780 1559.790 1207.920 ;
        RECT 1551.650 1207.720 1551.970 1207.780 ;
        RECT 1559.470 1207.720 1559.790 1207.780 ;
      LAYER via ;
        RECT 1551.680 1207.720 1551.940 1207.980 ;
        RECT 1559.500 1207.720 1559.760 1207.980 ;
      LAYER met2 ;
        RECT 1551.690 1219.680 1552.250 1228.680 ;
        RECT 1551.740 1208.010 1551.880 1219.680 ;
        RECT 1551.680 1207.690 1551.940 1208.010 ;
        RECT 1559.500 1207.690 1559.760 1208.010 ;
        RECT 1559.560 16.730 1559.700 1207.690 ;
        RECT 1559.560 16.590 1561.080 16.730 ;
        RECT 1560.940 2.400 1561.080 16.590 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1560.850 1207.920 1561.170 1207.980 ;
        RECT 1574.190 1207.920 1574.510 1207.980 ;
        RECT 1560.850 1207.780 1574.510 1207.920 ;
        RECT 1560.850 1207.720 1561.170 1207.780 ;
        RECT 1574.190 1207.720 1574.510 1207.780 ;
      LAYER via ;
        RECT 1560.880 1207.720 1561.140 1207.980 ;
        RECT 1574.220 1207.720 1574.480 1207.980 ;
      LAYER met2 ;
        RECT 1560.890 1219.680 1561.450 1228.680 ;
        RECT 1560.940 1208.010 1561.080 1219.680 ;
        RECT 1560.880 1207.690 1561.140 1208.010 ;
        RECT 1574.220 1207.690 1574.480 1208.010 ;
        RECT 1574.280 17.410 1574.420 1207.690 ;
        RECT 1574.280 17.270 1579.020 17.410 ;
        RECT 1578.880 2.400 1579.020 17.270 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1569.590 1213.360 1569.910 1213.420 ;
        RECT 1595.350 1213.360 1595.670 1213.420 ;
        RECT 1569.590 1213.220 1595.670 1213.360 ;
        RECT 1569.590 1213.160 1569.910 1213.220 ;
        RECT 1595.350 1213.160 1595.670 1213.220 ;
      LAYER via ;
        RECT 1569.620 1213.160 1569.880 1213.420 ;
        RECT 1595.380 1213.160 1595.640 1213.420 ;
      LAYER met2 ;
        RECT 1569.630 1219.680 1570.190 1228.680 ;
        RECT 1569.680 1213.450 1569.820 1219.680 ;
        RECT 1569.620 1213.130 1569.880 1213.450 ;
        RECT 1595.380 1213.130 1595.640 1213.450 ;
        RECT 1595.440 3.130 1595.580 1213.130 ;
        RECT 1595.440 2.990 1596.040 3.130 ;
        RECT 1595.900 2.960 1596.040 2.990 ;
        RECT 1595.900 2.820 1596.500 2.960 ;
        RECT 1596.360 2.400 1596.500 2.820 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 17.240 1580.030 17.300 ;
        RECT 1614.210 17.240 1614.530 17.300 ;
        RECT 1579.710 17.100 1614.530 17.240 ;
        RECT 1579.710 17.040 1580.030 17.100 ;
        RECT 1614.210 17.040 1614.530 17.100 ;
      LAYER via ;
        RECT 1579.740 17.040 1580.000 17.300 ;
        RECT 1614.240 17.040 1614.500 17.300 ;
      LAYER met2 ;
        RECT 1578.830 1220.330 1579.390 1228.680 ;
        RECT 1578.830 1220.190 1579.940 1220.330 ;
        RECT 1578.830 1219.680 1579.390 1220.190 ;
        RECT 1579.800 17.330 1579.940 1220.190 ;
        RECT 1579.740 17.010 1580.000 17.330 ;
        RECT 1614.240 17.010 1614.500 17.330 ;
        RECT 1614.300 2.400 1614.440 17.010 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.990 1211.320 1588.310 1211.380 ;
        RECT 1628.930 1211.320 1629.250 1211.380 ;
        RECT 1587.990 1211.180 1629.250 1211.320 ;
        RECT 1587.990 1211.120 1588.310 1211.180 ;
        RECT 1628.930 1211.120 1629.250 1211.180 ;
        RECT 1628.930 2.960 1629.250 3.020 ;
        RECT 1632.150 2.960 1632.470 3.020 ;
        RECT 1628.930 2.820 1632.470 2.960 ;
        RECT 1628.930 2.760 1629.250 2.820 ;
        RECT 1632.150 2.760 1632.470 2.820 ;
      LAYER via ;
        RECT 1588.020 1211.120 1588.280 1211.380 ;
        RECT 1628.960 1211.120 1629.220 1211.380 ;
        RECT 1628.960 2.760 1629.220 3.020 ;
        RECT 1632.180 2.760 1632.440 3.020 ;
      LAYER met2 ;
        RECT 1588.030 1219.680 1588.590 1228.680 ;
        RECT 1588.080 1211.410 1588.220 1219.680 ;
        RECT 1588.020 1211.090 1588.280 1211.410 ;
        RECT 1628.960 1211.090 1629.220 1211.410 ;
        RECT 1629.020 3.050 1629.160 1211.090 ;
        RECT 1628.960 2.730 1629.220 3.050 ;
        RECT 1632.180 2.730 1632.440 3.050 ;
        RECT 1632.240 2.400 1632.380 2.730 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1599.950 19.280 1600.270 19.340 ;
        RECT 1650.090 19.280 1650.410 19.340 ;
        RECT 1599.950 19.140 1650.410 19.280 ;
        RECT 1599.950 19.080 1600.270 19.140 ;
        RECT 1650.090 19.080 1650.410 19.140 ;
      LAYER via ;
        RECT 1599.980 19.080 1600.240 19.340 ;
        RECT 1650.120 19.080 1650.380 19.340 ;
      LAYER met2 ;
        RECT 1597.230 1220.330 1597.790 1228.680 ;
        RECT 1597.230 1220.190 1600.180 1220.330 ;
        RECT 1597.230 1219.680 1597.790 1220.190 ;
        RECT 1600.040 19.370 1600.180 1220.190 ;
        RECT 1599.980 19.050 1600.240 19.370 ;
        RECT 1650.120 19.050 1650.380 19.370 ;
        RECT 1650.180 2.400 1650.320 19.050 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1606.850 18.600 1607.170 18.660 ;
        RECT 1668.030 18.600 1668.350 18.660 ;
        RECT 1606.850 18.460 1668.350 18.600 ;
        RECT 1606.850 18.400 1607.170 18.460 ;
        RECT 1668.030 18.400 1668.350 18.460 ;
      LAYER via ;
        RECT 1606.880 18.400 1607.140 18.660 ;
        RECT 1668.060 18.400 1668.320 18.660 ;
      LAYER met2 ;
        RECT 1606.430 1220.330 1606.990 1228.680 ;
        RECT 1606.430 1219.680 1607.080 1220.330 ;
        RECT 1606.940 18.690 1607.080 1219.680 ;
        RECT 1606.880 18.370 1607.140 18.690 ;
        RECT 1668.060 18.370 1668.320 18.690 ;
        RECT 1668.120 2.400 1668.260 18.370 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1615.590 1207.580 1615.910 1207.640 ;
        RECT 1620.650 1207.580 1620.970 1207.640 ;
        RECT 1615.590 1207.440 1620.970 1207.580 ;
        RECT 1615.590 1207.380 1615.910 1207.440 ;
        RECT 1620.650 1207.380 1620.970 1207.440 ;
        RECT 1620.650 20.640 1620.970 20.700 ;
        RECT 1685.510 20.640 1685.830 20.700 ;
        RECT 1620.650 20.500 1685.830 20.640 ;
        RECT 1620.650 20.440 1620.970 20.500 ;
        RECT 1685.510 20.440 1685.830 20.500 ;
      LAYER via ;
        RECT 1615.620 1207.380 1615.880 1207.640 ;
        RECT 1620.680 1207.380 1620.940 1207.640 ;
        RECT 1620.680 20.440 1620.940 20.700 ;
        RECT 1685.540 20.440 1685.800 20.700 ;
      LAYER met2 ;
        RECT 1615.630 1219.680 1616.190 1228.680 ;
        RECT 1615.680 1207.670 1615.820 1219.680 ;
        RECT 1615.620 1207.350 1615.880 1207.670 ;
        RECT 1620.680 1207.350 1620.940 1207.670 ;
        RECT 1620.740 20.730 1620.880 1207.350 ;
        RECT 1620.680 20.410 1620.940 20.730 ;
        RECT 1685.540 20.410 1685.800 20.730 ;
        RECT 1685.600 2.400 1685.740 20.410 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 35.260 722.590 35.320 ;
        RECT 1117.870 35.260 1118.190 35.320 ;
        RECT 722.270 35.120 1118.190 35.260 ;
        RECT 722.270 35.060 722.590 35.120 ;
        RECT 1117.870 35.060 1118.190 35.120 ;
      LAYER via ;
        RECT 722.300 35.060 722.560 35.320 ;
        RECT 1117.900 35.060 1118.160 35.320 ;
      LAYER met2 ;
        RECT 1120.670 1221.010 1121.230 1228.680 ;
        RECT 1118.420 1220.870 1121.230 1221.010 ;
        RECT 1118.420 1196.700 1118.560 1220.870 ;
        RECT 1120.670 1219.680 1121.230 1220.870 ;
        RECT 1117.960 1196.560 1118.560 1196.700 ;
        RECT 1117.960 35.350 1118.100 1196.560 ;
        RECT 722.300 35.030 722.560 35.350 ;
        RECT 1117.900 35.030 1118.160 35.350 ;
        RECT 722.360 2.400 722.500 35.030 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1624.790 1211.660 1625.110 1211.720 ;
        RECT 1652.390 1211.660 1652.710 1211.720 ;
        RECT 1624.790 1211.520 1652.710 1211.660 ;
        RECT 1624.790 1211.460 1625.110 1211.520 ;
        RECT 1652.390 1211.460 1652.710 1211.520 ;
        RECT 1652.390 16.560 1652.710 16.620 ;
        RECT 1703.450 16.560 1703.770 16.620 ;
        RECT 1652.390 16.420 1703.770 16.560 ;
        RECT 1652.390 16.360 1652.710 16.420 ;
        RECT 1703.450 16.360 1703.770 16.420 ;
      LAYER via ;
        RECT 1624.820 1211.460 1625.080 1211.720 ;
        RECT 1652.420 1211.460 1652.680 1211.720 ;
        RECT 1652.420 16.360 1652.680 16.620 ;
        RECT 1703.480 16.360 1703.740 16.620 ;
      LAYER met2 ;
        RECT 1624.830 1219.680 1625.390 1228.680 ;
        RECT 1624.880 1211.750 1625.020 1219.680 ;
        RECT 1624.820 1211.430 1625.080 1211.750 ;
        RECT 1652.420 1211.430 1652.680 1211.750 ;
        RECT 1652.480 16.650 1652.620 1211.430 ;
        RECT 1652.420 16.330 1652.680 16.650 ;
        RECT 1703.480 16.330 1703.740 16.650 ;
        RECT 1703.540 2.400 1703.680 16.330 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1633.990 1212.000 1634.310 1212.060 ;
        RECT 1714.490 1212.000 1714.810 1212.060 ;
        RECT 1633.990 1211.860 1714.810 1212.000 ;
        RECT 1633.990 1211.800 1634.310 1211.860 ;
        RECT 1714.490 1211.800 1714.810 1211.860 ;
        RECT 1714.490 20.640 1714.810 20.700 ;
        RECT 1721.390 20.640 1721.710 20.700 ;
        RECT 1714.490 20.500 1721.710 20.640 ;
        RECT 1714.490 20.440 1714.810 20.500 ;
        RECT 1721.390 20.440 1721.710 20.500 ;
      LAYER via ;
        RECT 1634.020 1211.800 1634.280 1212.060 ;
        RECT 1714.520 1211.800 1714.780 1212.060 ;
        RECT 1714.520 20.440 1714.780 20.700 ;
        RECT 1721.420 20.440 1721.680 20.700 ;
      LAYER met2 ;
        RECT 1634.030 1219.680 1634.590 1228.680 ;
        RECT 1634.080 1212.090 1634.220 1219.680 ;
        RECT 1634.020 1211.770 1634.280 1212.090 ;
        RECT 1714.520 1211.770 1714.780 1212.090 ;
        RECT 1714.580 20.730 1714.720 1211.770 ;
        RECT 1714.520 20.410 1714.780 20.730 ;
        RECT 1721.420 20.410 1721.680 20.730 ;
        RECT 1721.480 2.400 1721.620 20.410 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1709.965 1212.185 1710.135 1213.375 ;
      LAYER mcon ;
        RECT 1709.965 1213.205 1710.135 1213.375 ;
      LAYER met1 ;
        RECT 1643.190 1213.360 1643.510 1213.420 ;
        RECT 1709.905 1213.360 1710.195 1213.405 ;
        RECT 1643.190 1213.220 1710.195 1213.360 ;
        RECT 1643.190 1213.160 1643.510 1213.220 ;
        RECT 1709.905 1213.175 1710.195 1213.220 ;
        RECT 1709.905 1212.340 1710.195 1212.385 ;
        RECT 1739.790 1212.340 1740.110 1212.400 ;
        RECT 1709.905 1212.200 1740.110 1212.340 ;
        RECT 1709.905 1212.155 1710.195 1212.200 ;
        RECT 1739.790 1212.140 1740.110 1212.200 ;
      LAYER via ;
        RECT 1643.220 1213.160 1643.480 1213.420 ;
        RECT 1739.820 1212.140 1740.080 1212.400 ;
      LAYER met2 ;
        RECT 1643.230 1219.680 1643.790 1228.680 ;
        RECT 1643.280 1213.450 1643.420 1219.680 ;
        RECT 1643.220 1213.130 1643.480 1213.450 ;
        RECT 1739.820 1212.110 1740.080 1212.430 ;
        RECT 1739.880 3.130 1740.020 1212.110 ;
        RECT 1739.420 2.990 1740.020 3.130 ;
        RECT 1739.420 2.400 1739.560 2.990 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1720.545 1208.445 1720.715 1209.635 ;
      LAYER mcon ;
        RECT 1720.545 1209.465 1720.715 1209.635 ;
      LAYER met1 ;
        RECT 1720.485 1209.620 1720.775 1209.665 ;
        RECT 1754.050 1209.620 1754.370 1209.680 ;
        RECT 1720.485 1209.480 1754.370 1209.620 ;
        RECT 1720.485 1209.435 1720.775 1209.480 ;
        RECT 1754.050 1209.420 1754.370 1209.480 ;
        RECT 1653.770 1208.600 1654.090 1208.660 ;
        RECT 1720.485 1208.600 1720.775 1208.645 ;
        RECT 1653.770 1208.460 1720.775 1208.600 ;
        RECT 1653.770 1208.400 1654.090 1208.460 ;
        RECT 1720.485 1208.415 1720.775 1208.460 ;
        RECT 1754.050 2.960 1754.370 3.020 ;
        RECT 1756.810 2.960 1757.130 3.020 ;
        RECT 1754.050 2.820 1757.130 2.960 ;
        RECT 1754.050 2.760 1754.370 2.820 ;
        RECT 1756.810 2.760 1757.130 2.820 ;
      LAYER via ;
        RECT 1754.080 1209.420 1754.340 1209.680 ;
        RECT 1653.800 1208.400 1654.060 1208.660 ;
        RECT 1754.080 2.760 1754.340 3.020 ;
        RECT 1756.840 2.760 1757.100 3.020 ;
      LAYER met2 ;
        RECT 1652.430 1220.330 1652.990 1228.680 ;
        RECT 1652.430 1220.190 1654.000 1220.330 ;
        RECT 1652.430 1219.680 1652.990 1220.190 ;
        RECT 1653.860 1208.690 1654.000 1220.190 ;
        RECT 1754.080 1209.390 1754.340 1209.710 ;
        RECT 1653.800 1208.370 1654.060 1208.690 ;
        RECT 1754.140 3.050 1754.280 1209.390 ;
        RECT 1754.080 2.730 1754.340 3.050 ;
        RECT 1756.840 2.730 1757.100 3.050 ;
        RECT 1756.900 2.400 1757.040 2.730 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1728.365 1210.825 1728.535 1212.695 ;
        RECT 1752.745 1208.445 1752.915 1212.695 ;
        RECT 1766.545 1207.425 1766.715 1208.615 ;
      LAYER mcon ;
        RECT 1728.365 1212.525 1728.535 1212.695 ;
        RECT 1752.745 1212.525 1752.915 1212.695 ;
        RECT 1766.545 1208.445 1766.715 1208.615 ;
      LAYER met1 ;
        RECT 1728.305 1212.680 1728.595 1212.725 ;
        RECT 1752.685 1212.680 1752.975 1212.725 ;
        RECT 1728.305 1212.540 1752.975 1212.680 ;
        RECT 1728.305 1212.495 1728.595 1212.540 ;
        RECT 1752.685 1212.495 1752.975 1212.540 ;
        RECT 1661.590 1210.980 1661.910 1211.040 ;
        RECT 1728.305 1210.980 1728.595 1211.025 ;
        RECT 1661.590 1210.840 1728.595 1210.980 ;
        RECT 1661.590 1210.780 1661.910 1210.840 ;
        RECT 1728.305 1210.795 1728.595 1210.840 ;
        RECT 1752.685 1208.600 1752.975 1208.645 ;
        RECT 1766.485 1208.600 1766.775 1208.645 ;
        RECT 1752.685 1208.460 1766.775 1208.600 ;
        RECT 1752.685 1208.415 1752.975 1208.460 ;
        RECT 1766.485 1208.415 1766.775 1208.460 ;
        RECT 1766.485 1207.580 1766.775 1207.625 ;
        RECT 1773.830 1207.580 1774.150 1207.640 ;
        RECT 1766.485 1207.440 1774.150 1207.580 ;
        RECT 1766.485 1207.395 1766.775 1207.440 ;
        RECT 1773.830 1207.380 1774.150 1207.440 ;
      LAYER via ;
        RECT 1661.620 1210.780 1661.880 1211.040 ;
        RECT 1773.860 1207.380 1774.120 1207.640 ;
      LAYER met2 ;
        RECT 1661.630 1219.680 1662.190 1228.680 ;
        RECT 1661.680 1211.070 1661.820 1219.680 ;
        RECT 1661.620 1210.750 1661.880 1211.070 ;
        RECT 1773.860 1207.350 1774.120 1207.670 ;
        RECT 1773.920 1206.730 1774.060 1207.350 ;
        RECT 1773.920 1206.590 1774.520 1206.730 ;
        RECT 1774.380 3.130 1774.520 1206.590 ;
        RECT 1774.380 2.990 1774.980 3.130 ;
        RECT 1774.840 2.400 1774.980 2.990 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1670.790 1208.940 1671.110 1209.000 ;
        RECT 1670.790 1208.800 1769.920 1208.940 ;
        RECT 1670.790 1208.740 1671.110 1208.800 ;
        RECT 1769.780 1208.600 1769.920 1208.800 ;
        RECT 1787.170 1208.600 1787.490 1208.660 ;
        RECT 1769.780 1208.460 1787.490 1208.600 ;
        RECT 1787.170 1208.400 1787.490 1208.460 ;
        RECT 1787.170 62.120 1787.490 62.180 ;
        RECT 1792.690 62.120 1793.010 62.180 ;
        RECT 1787.170 61.980 1793.010 62.120 ;
        RECT 1787.170 61.920 1787.490 61.980 ;
        RECT 1792.690 61.920 1793.010 61.980 ;
      LAYER via ;
        RECT 1670.820 1208.740 1671.080 1209.000 ;
        RECT 1787.200 1208.400 1787.460 1208.660 ;
        RECT 1787.200 61.920 1787.460 62.180 ;
        RECT 1792.720 61.920 1792.980 62.180 ;
      LAYER met2 ;
        RECT 1670.830 1219.680 1671.390 1228.680 ;
        RECT 1670.880 1209.030 1671.020 1219.680 ;
        RECT 1670.820 1208.710 1671.080 1209.030 ;
        RECT 1787.200 1208.370 1787.460 1208.690 ;
        RECT 1787.260 62.210 1787.400 1208.370 ;
        RECT 1787.200 61.890 1787.460 62.210 ;
        RECT 1792.720 61.890 1792.980 62.210 ;
        RECT 1792.780 2.400 1792.920 61.890 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1809.250 1212.340 1809.570 1212.400 ;
        RECT 1798.300 1212.200 1809.570 1212.340 ;
        RECT 1679.990 1211.660 1680.310 1211.720 ;
        RECT 1776.130 1211.660 1776.450 1211.720 ;
        RECT 1679.990 1211.520 1776.450 1211.660 ;
        RECT 1679.990 1211.460 1680.310 1211.520 ;
        RECT 1776.130 1211.460 1776.450 1211.520 ;
        RECT 1777.510 1211.660 1777.830 1211.720 ;
        RECT 1798.300 1211.660 1798.440 1212.200 ;
        RECT 1809.250 1212.140 1809.570 1212.200 ;
        RECT 1777.510 1211.520 1798.440 1211.660 ;
        RECT 1777.510 1211.460 1777.830 1211.520 ;
        RECT 1809.250 2.960 1809.570 3.020 ;
        RECT 1810.630 2.960 1810.950 3.020 ;
        RECT 1809.250 2.820 1810.950 2.960 ;
        RECT 1809.250 2.760 1809.570 2.820 ;
        RECT 1810.630 2.760 1810.950 2.820 ;
      LAYER via ;
        RECT 1680.020 1211.460 1680.280 1211.720 ;
        RECT 1776.160 1211.460 1776.420 1211.720 ;
        RECT 1777.540 1211.460 1777.800 1211.720 ;
        RECT 1809.280 1212.140 1809.540 1212.400 ;
        RECT 1809.280 2.760 1809.540 3.020 ;
        RECT 1810.660 2.760 1810.920 3.020 ;
      LAYER met2 ;
        RECT 1680.030 1219.680 1680.590 1228.680 ;
        RECT 1680.080 1211.750 1680.220 1219.680 ;
        RECT 1809.280 1212.110 1809.540 1212.430 ;
        RECT 1680.020 1211.430 1680.280 1211.750 ;
        RECT 1776.160 1211.490 1776.420 1211.750 ;
        RECT 1777.540 1211.490 1777.800 1211.750 ;
        RECT 1776.160 1211.430 1777.800 1211.490 ;
        RECT 1776.220 1211.350 1777.740 1211.430 ;
        RECT 1809.340 3.050 1809.480 1212.110 ;
        RECT 1809.280 2.730 1809.540 3.050 ;
        RECT 1810.660 2.730 1810.920 3.050 ;
        RECT 1810.720 2.400 1810.860 2.730 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1776.665 1208.785 1776.835 1211.335 ;
      LAYER mcon ;
        RECT 1776.665 1211.165 1776.835 1211.335 ;
      LAYER met1 ;
        RECT 1688.730 1211.320 1689.050 1211.380 ;
        RECT 1776.605 1211.320 1776.895 1211.365 ;
        RECT 1688.730 1211.180 1776.895 1211.320 ;
        RECT 1688.730 1211.120 1689.050 1211.180 ;
        RECT 1776.605 1211.135 1776.895 1211.180 ;
        RECT 1776.605 1208.940 1776.895 1208.985 ;
        RECT 1829.030 1208.940 1829.350 1209.000 ;
        RECT 1776.605 1208.800 1829.350 1208.940 ;
        RECT 1776.605 1208.755 1776.895 1208.800 ;
        RECT 1829.030 1208.740 1829.350 1208.800 ;
      LAYER via ;
        RECT 1688.760 1211.120 1689.020 1211.380 ;
        RECT 1829.060 1208.740 1829.320 1209.000 ;
      LAYER met2 ;
        RECT 1688.770 1219.680 1689.330 1228.680 ;
        RECT 1688.820 1211.410 1688.960 1219.680 ;
        RECT 1688.760 1211.090 1689.020 1211.410 ;
        RECT 1829.060 1208.710 1829.320 1209.030 ;
        RECT 1829.120 3.130 1829.260 1208.710 ;
        RECT 1828.660 2.990 1829.260 3.130 ;
        RECT 1828.660 2.400 1828.800 2.990 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.930 1209.280 1698.250 1209.340 ;
        RECT 1842.370 1209.280 1842.690 1209.340 ;
        RECT 1697.930 1209.140 1842.690 1209.280 ;
        RECT 1697.930 1209.080 1698.250 1209.140 ;
        RECT 1842.370 1209.080 1842.690 1209.140 ;
        RECT 1842.370 2.960 1842.690 3.020 ;
        RECT 1846.050 2.960 1846.370 3.020 ;
        RECT 1842.370 2.820 1846.370 2.960 ;
        RECT 1842.370 2.760 1842.690 2.820 ;
        RECT 1846.050 2.760 1846.370 2.820 ;
      LAYER via ;
        RECT 1697.960 1209.080 1698.220 1209.340 ;
        RECT 1842.400 1209.080 1842.660 1209.340 ;
        RECT 1842.400 2.760 1842.660 3.020 ;
        RECT 1846.080 2.760 1846.340 3.020 ;
      LAYER met2 ;
        RECT 1697.970 1219.680 1698.530 1228.680 ;
        RECT 1698.020 1209.370 1698.160 1219.680 ;
        RECT 1697.960 1209.050 1698.220 1209.370 ;
        RECT 1842.400 1209.050 1842.660 1209.370 ;
        RECT 1842.460 3.050 1842.600 1209.050 ;
        RECT 1842.400 2.730 1842.660 3.050 ;
        RECT 1846.080 2.730 1846.340 3.050 ;
        RECT 1846.140 2.400 1846.280 2.730 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1729.745 1209.805 1729.915 1214.395 ;
      LAYER mcon ;
        RECT 1729.745 1214.225 1729.915 1214.395 ;
      LAYER met1 ;
        RECT 1707.130 1214.380 1707.450 1214.440 ;
        RECT 1729.685 1214.380 1729.975 1214.425 ;
        RECT 1707.130 1214.240 1729.975 1214.380 ;
        RECT 1707.130 1214.180 1707.450 1214.240 ;
        RECT 1729.685 1214.195 1729.975 1214.240 ;
        RECT 1729.685 1209.960 1729.975 1210.005 ;
        RECT 1863.990 1209.960 1864.310 1210.020 ;
        RECT 1729.685 1209.820 1864.310 1209.960 ;
        RECT 1729.685 1209.775 1729.975 1209.820 ;
        RECT 1863.990 1209.760 1864.310 1209.820 ;
        RECT 1863.070 2.960 1863.390 3.020 ;
        RECT 1863.990 2.960 1864.310 3.020 ;
        RECT 1863.070 2.820 1864.310 2.960 ;
        RECT 1863.070 2.760 1863.390 2.820 ;
        RECT 1863.990 2.760 1864.310 2.820 ;
      LAYER via ;
        RECT 1707.160 1214.180 1707.420 1214.440 ;
        RECT 1864.020 1209.760 1864.280 1210.020 ;
        RECT 1863.100 2.760 1863.360 3.020 ;
        RECT 1864.020 2.760 1864.280 3.020 ;
      LAYER met2 ;
        RECT 1707.170 1219.680 1707.730 1228.680 ;
        RECT 1707.220 1214.470 1707.360 1219.680 ;
        RECT 1707.160 1214.150 1707.420 1214.470 ;
        RECT 1864.020 1209.730 1864.280 1210.050 ;
        RECT 1864.080 1206.730 1864.220 1209.730 ;
        RECT 1863.160 1206.590 1864.220 1206.730 ;
        RECT 1863.160 3.050 1863.300 1206.590 ;
        RECT 1863.100 2.730 1863.360 3.050 ;
        RECT 1864.020 2.730 1864.280 3.050 ;
        RECT 1864.080 2.400 1864.220 2.730 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1125.765 1104.065 1125.935 1111.035 ;
      LAYER mcon ;
        RECT 1125.765 1110.865 1125.935 1111.035 ;
      LAYER met1 ;
        RECT 1125.230 1159.300 1125.550 1159.360 ;
        RECT 1128.450 1159.300 1128.770 1159.360 ;
        RECT 1125.230 1159.160 1128.770 1159.300 ;
        RECT 1125.230 1159.100 1125.550 1159.160 ;
        RECT 1128.450 1159.100 1128.770 1159.160 ;
        RECT 1125.690 1111.020 1126.010 1111.080 ;
        RECT 1125.495 1110.880 1126.010 1111.020 ;
        RECT 1125.690 1110.820 1126.010 1110.880 ;
        RECT 1125.690 1104.220 1126.010 1104.280 ;
        RECT 1125.495 1104.080 1126.010 1104.220 ;
        RECT 1125.690 1104.020 1126.010 1104.080 ;
        RECT 1125.230 241.300 1125.550 241.360 ;
        RECT 1125.690 241.300 1126.010 241.360 ;
        RECT 1125.230 241.160 1126.010 241.300 ;
        RECT 1125.230 241.100 1125.550 241.160 ;
        RECT 1125.690 241.100 1126.010 241.160 ;
        RECT 740.210 34.920 740.530 34.980 ;
        RECT 1125.690 34.920 1126.010 34.980 ;
        RECT 740.210 34.780 1126.010 34.920 ;
        RECT 740.210 34.720 740.530 34.780 ;
        RECT 1125.690 34.720 1126.010 34.780 ;
      LAYER via ;
        RECT 1125.260 1159.100 1125.520 1159.360 ;
        RECT 1128.480 1159.100 1128.740 1159.360 ;
        RECT 1125.720 1110.820 1125.980 1111.080 ;
        RECT 1125.720 1104.020 1125.980 1104.280 ;
        RECT 1125.260 241.100 1125.520 241.360 ;
        RECT 1125.720 241.100 1125.980 241.360 ;
        RECT 740.240 34.720 740.500 34.980 ;
        RECT 1125.720 34.720 1125.980 34.980 ;
      LAYER met2 ;
        RECT 1129.870 1220.330 1130.430 1228.680 ;
        RECT 1128.540 1220.190 1130.430 1220.330 ;
        RECT 1128.540 1159.390 1128.680 1220.190 ;
        RECT 1129.870 1219.680 1130.430 1220.190 ;
        RECT 1125.260 1159.245 1125.520 1159.390 ;
        RECT 1125.250 1158.875 1125.530 1159.245 ;
        RECT 1126.170 1158.875 1126.450 1159.245 ;
        RECT 1128.480 1159.070 1128.740 1159.390 ;
        RECT 1126.240 1152.330 1126.380 1158.875 ;
        RECT 1125.780 1152.190 1126.380 1152.330 ;
        RECT 1125.780 1111.110 1125.920 1152.190 ;
        RECT 1125.720 1110.790 1125.980 1111.110 ;
        RECT 1125.720 1104.165 1125.980 1104.310 ;
        RECT 1125.710 1103.795 1125.990 1104.165 ;
        RECT 1126.630 1103.795 1126.910 1104.165 ;
        RECT 1126.700 1079.570 1126.840 1103.795 ;
        RECT 1125.780 1079.430 1126.840 1079.570 ;
        RECT 1125.780 980.290 1125.920 1079.430 ;
        RECT 1125.320 980.150 1125.920 980.290 ;
        RECT 1125.320 979.610 1125.460 980.150 ;
        RECT 1125.320 979.470 1125.920 979.610 ;
        RECT 1125.780 883.050 1125.920 979.470 ;
        RECT 1125.320 882.910 1125.920 883.050 ;
        RECT 1125.320 881.690 1125.460 882.910 ;
        RECT 1125.320 881.550 1125.920 881.690 ;
        RECT 1125.780 690.610 1125.920 881.550 ;
        RECT 1125.320 690.470 1125.920 690.610 ;
        RECT 1125.320 688.570 1125.460 690.470 ;
        RECT 1125.320 688.430 1125.920 688.570 ;
        RECT 1125.780 265.610 1125.920 688.430 ;
        RECT 1125.320 265.470 1125.920 265.610 ;
        RECT 1125.320 241.390 1125.460 265.470 ;
        RECT 1125.260 241.070 1125.520 241.390 ;
        RECT 1125.720 241.070 1125.980 241.390 ;
        RECT 1125.780 35.010 1125.920 241.070 ;
        RECT 740.240 34.690 740.500 35.010 ;
        RECT 1125.720 34.690 1125.980 35.010 ;
        RECT 740.300 2.400 740.440 34.690 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 1125.250 1158.920 1125.530 1159.200 ;
        RECT 1126.170 1158.920 1126.450 1159.200 ;
        RECT 1125.710 1103.840 1125.990 1104.120 ;
        RECT 1126.630 1103.840 1126.910 1104.120 ;
      LAYER met3 ;
        RECT 1125.225 1159.210 1125.555 1159.225 ;
        RECT 1126.145 1159.210 1126.475 1159.225 ;
        RECT 1125.225 1158.910 1126.475 1159.210 ;
        RECT 1125.225 1158.895 1125.555 1158.910 ;
        RECT 1126.145 1158.895 1126.475 1158.910 ;
        RECT 1125.685 1104.130 1126.015 1104.145 ;
        RECT 1126.605 1104.130 1126.935 1104.145 ;
        RECT 1125.685 1103.830 1126.935 1104.130 ;
        RECT 1125.685 1103.815 1126.015 1103.830 ;
        RECT 1126.605 1103.815 1126.935 1103.830 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1751.825 1213.885 1752.455 1214.055 ;
        RECT 1751.825 1213.545 1751.995 1213.885 ;
        RECT 1823.125 1212.185 1823.295 1214.055 ;
        RECT 1836.005 1207.765 1836.175 1212.355 ;
      LAYER mcon ;
        RECT 1752.285 1213.885 1752.455 1214.055 ;
        RECT 1823.125 1213.885 1823.295 1214.055 ;
        RECT 1836.005 1212.185 1836.175 1212.355 ;
      LAYER met1 ;
        RECT 1752.225 1214.040 1752.515 1214.085 ;
        RECT 1823.065 1214.040 1823.355 1214.085 ;
        RECT 1752.225 1213.900 1823.355 1214.040 ;
        RECT 1752.225 1213.855 1752.515 1213.900 ;
        RECT 1823.065 1213.855 1823.355 1213.900 ;
        RECT 1716.330 1213.700 1716.650 1213.760 ;
        RECT 1751.765 1213.700 1752.055 1213.745 ;
        RECT 1716.330 1213.560 1752.055 1213.700 ;
        RECT 1716.330 1213.500 1716.650 1213.560 ;
        RECT 1751.765 1213.515 1752.055 1213.560 ;
        RECT 1823.065 1212.340 1823.355 1212.385 ;
        RECT 1835.945 1212.340 1836.235 1212.385 ;
        RECT 1823.065 1212.200 1836.235 1212.340 ;
        RECT 1823.065 1212.155 1823.355 1212.200 ;
        RECT 1835.945 1212.155 1836.235 1212.200 ;
        RECT 1835.945 1207.920 1836.235 1207.965 ;
        RECT 1877.790 1207.920 1878.110 1207.980 ;
        RECT 1835.945 1207.780 1878.110 1207.920 ;
        RECT 1835.945 1207.735 1836.235 1207.780 ;
        RECT 1877.790 1207.720 1878.110 1207.780 ;
        RECT 1877.790 62.120 1878.110 62.180 ;
        RECT 1881.930 62.120 1882.250 62.180 ;
        RECT 1877.790 61.980 1882.250 62.120 ;
        RECT 1877.790 61.920 1878.110 61.980 ;
        RECT 1881.930 61.920 1882.250 61.980 ;
      LAYER via ;
        RECT 1716.360 1213.500 1716.620 1213.760 ;
        RECT 1877.820 1207.720 1878.080 1207.980 ;
        RECT 1877.820 61.920 1878.080 62.180 ;
        RECT 1881.960 61.920 1882.220 62.180 ;
      LAYER met2 ;
        RECT 1716.370 1219.680 1716.930 1228.680 ;
        RECT 1716.420 1213.790 1716.560 1219.680 ;
        RECT 1716.360 1213.470 1716.620 1213.790 ;
        RECT 1877.820 1207.690 1878.080 1208.010 ;
        RECT 1877.880 62.210 1878.020 1207.690 ;
        RECT 1877.820 61.890 1878.080 62.210 ;
        RECT 1881.960 61.890 1882.220 62.210 ;
        RECT 1882.020 2.400 1882.160 61.890 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.125 1212.865 1754.295 1214.735 ;
        RECT 1836.005 1212.865 1837.095 1213.035 ;
      LAYER mcon ;
        RECT 1754.125 1214.565 1754.295 1214.735 ;
        RECT 1836.925 1212.865 1837.095 1213.035 ;
      LAYER met1 ;
        RECT 1754.065 1214.720 1754.355 1214.765 ;
        RECT 1751.380 1214.580 1754.355 1214.720 ;
        RECT 1725.530 1214.040 1725.850 1214.100 ;
        RECT 1751.380 1214.040 1751.520 1214.580 ;
        RECT 1754.065 1214.535 1754.355 1214.580 ;
        RECT 1725.530 1213.900 1751.520 1214.040 ;
        RECT 1725.530 1213.840 1725.850 1213.900 ;
        RECT 1754.065 1213.020 1754.355 1213.065 ;
        RECT 1835.945 1213.020 1836.235 1213.065 ;
        RECT 1754.065 1212.880 1836.235 1213.020 ;
        RECT 1754.065 1212.835 1754.355 1212.880 ;
        RECT 1835.945 1212.835 1836.235 1212.880 ;
        RECT 1836.865 1213.020 1837.155 1213.065 ;
        RECT 1898.490 1213.020 1898.810 1213.080 ;
        RECT 1836.865 1212.880 1898.810 1213.020 ;
        RECT 1836.865 1212.835 1837.155 1212.880 ;
        RECT 1898.490 1212.820 1898.810 1212.880 ;
        RECT 1898.490 2.960 1898.810 3.020 ;
        RECT 1899.870 2.960 1900.190 3.020 ;
        RECT 1898.490 2.820 1900.190 2.960 ;
        RECT 1898.490 2.760 1898.810 2.820 ;
        RECT 1899.870 2.760 1900.190 2.820 ;
      LAYER via ;
        RECT 1725.560 1213.840 1725.820 1214.100 ;
        RECT 1898.520 1212.820 1898.780 1213.080 ;
        RECT 1898.520 2.760 1898.780 3.020 ;
        RECT 1899.900 2.760 1900.160 3.020 ;
      LAYER met2 ;
        RECT 1725.570 1219.680 1726.130 1228.680 ;
        RECT 1725.620 1214.130 1725.760 1219.680 ;
        RECT 1725.560 1213.810 1725.820 1214.130 ;
        RECT 1898.520 1212.790 1898.780 1213.110 ;
        RECT 1898.580 3.050 1898.720 1212.790 ;
        RECT 1898.520 2.730 1898.780 3.050 ;
        RECT 1899.900 2.730 1900.160 3.050 ;
        RECT 1899.960 2.400 1900.100 2.730 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1777.125 1211.165 1777.295 1216.095 ;
      LAYER mcon ;
        RECT 1777.125 1215.925 1777.295 1216.095 ;
      LAYER met1 ;
        RECT 1734.730 1216.080 1735.050 1216.140 ;
        RECT 1777.065 1216.080 1777.355 1216.125 ;
        RECT 1734.730 1215.940 1777.355 1216.080 ;
        RECT 1734.730 1215.880 1735.050 1215.940 ;
        RECT 1777.065 1215.895 1777.355 1215.940 ;
        RECT 1847.890 1212.000 1848.210 1212.060 ;
        RECT 1912.290 1212.000 1912.610 1212.060 ;
        RECT 1847.890 1211.860 1912.610 1212.000 ;
        RECT 1847.890 1211.800 1848.210 1211.860 ;
        RECT 1912.290 1211.800 1912.610 1211.860 ;
        RECT 1777.065 1211.320 1777.355 1211.365 ;
        RECT 1787.170 1211.320 1787.490 1211.380 ;
        RECT 1777.065 1211.180 1787.490 1211.320 ;
        RECT 1777.065 1211.135 1777.355 1211.180 ;
        RECT 1787.170 1211.120 1787.490 1211.180 ;
        RECT 1912.290 2.960 1912.610 3.020 ;
        RECT 1917.810 2.960 1918.130 3.020 ;
        RECT 1912.290 2.820 1918.130 2.960 ;
        RECT 1912.290 2.760 1912.610 2.820 ;
        RECT 1917.810 2.760 1918.130 2.820 ;
      LAYER via ;
        RECT 1734.760 1215.880 1735.020 1216.140 ;
        RECT 1847.920 1211.800 1848.180 1212.060 ;
        RECT 1912.320 1211.800 1912.580 1212.060 ;
        RECT 1787.200 1211.120 1787.460 1211.380 ;
        RECT 1912.320 2.760 1912.580 3.020 ;
        RECT 1917.840 2.760 1918.100 3.020 ;
      LAYER met2 ;
        RECT 1734.770 1219.680 1735.330 1228.680 ;
        RECT 1734.820 1216.170 1734.960 1219.680 ;
        RECT 1734.760 1215.850 1735.020 1216.170 ;
        RECT 1835.950 1212.000 1836.230 1212.285 ;
        RECT 1835.100 1211.915 1836.230 1212.000 ;
        RECT 1847.910 1211.915 1848.190 1212.285 ;
        RECT 1835.100 1211.860 1836.160 1211.915 ;
        RECT 1835.100 1211.605 1835.240 1211.860 ;
        RECT 1847.920 1211.770 1848.180 1211.915 ;
        RECT 1912.320 1211.770 1912.580 1212.090 ;
        RECT 1787.200 1211.090 1787.460 1211.410 ;
        RECT 1787.650 1211.235 1787.930 1211.605 ;
        RECT 1835.030 1211.235 1835.310 1211.605 ;
        RECT 1787.260 1210.810 1787.400 1211.090 ;
        RECT 1787.720 1210.810 1787.860 1211.235 ;
        RECT 1787.260 1210.670 1787.860 1210.810 ;
        RECT 1912.380 3.050 1912.520 1211.770 ;
        RECT 1912.320 2.730 1912.580 3.050 ;
        RECT 1917.840 2.730 1918.100 3.050 ;
        RECT 1917.900 2.400 1918.040 2.730 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
      LAYER via2 ;
        RECT 1835.950 1211.960 1836.230 1212.240 ;
        RECT 1847.910 1211.960 1848.190 1212.240 ;
        RECT 1787.650 1211.280 1787.930 1211.560 ;
        RECT 1835.030 1211.280 1835.310 1211.560 ;
      LAYER met3 ;
        RECT 1835.925 1212.250 1836.255 1212.265 ;
        RECT 1847.885 1212.250 1848.215 1212.265 ;
        RECT 1835.925 1211.950 1848.215 1212.250 ;
        RECT 1835.925 1211.935 1836.255 1211.950 ;
        RECT 1847.885 1211.935 1848.215 1211.950 ;
        RECT 1787.625 1211.570 1787.955 1211.585 ;
        RECT 1835.005 1211.570 1835.335 1211.585 ;
        RECT 1787.625 1211.270 1835.335 1211.570 ;
        RECT 1787.625 1211.255 1787.955 1211.270 ;
        RECT 1835.005 1211.255 1835.335 1211.270 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1897.645 1213.205 1898.275 1213.375 ;
        RECT 1897.645 1210.825 1897.815 1213.205 ;
      LAYER mcon ;
        RECT 1898.105 1213.205 1898.275 1213.375 ;
      LAYER met1 ;
        RECT 1898.045 1213.360 1898.335 1213.405 ;
        RECT 1928.390 1213.360 1928.710 1213.420 ;
        RECT 1898.045 1213.220 1928.710 1213.360 ;
        RECT 1898.045 1213.175 1898.335 1213.220 ;
        RECT 1928.390 1213.160 1928.710 1213.220 ;
        RECT 1743.930 1210.980 1744.250 1211.040 ;
        RECT 1897.585 1210.980 1897.875 1211.025 ;
        RECT 1743.930 1210.840 1897.875 1210.980 ;
        RECT 1743.930 1210.780 1744.250 1210.840 ;
        RECT 1897.585 1210.795 1897.875 1210.840 ;
        RECT 1928.390 20.640 1928.710 20.700 ;
        RECT 1935.290 20.640 1935.610 20.700 ;
        RECT 1928.390 20.500 1935.610 20.640 ;
        RECT 1928.390 20.440 1928.710 20.500 ;
        RECT 1935.290 20.440 1935.610 20.500 ;
      LAYER via ;
        RECT 1928.420 1213.160 1928.680 1213.420 ;
        RECT 1743.960 1210.780 1744.220 1211.040 ;
        RECT 1928.420 20.440 1928.680 20.700 ;
        RECT 1935.320 20.440 1935.580 20.700 ;
      LAYER met2 ;
        RECT 1743.970 1219.680 1744.530 1228.680 ;
        RECT 1744.020 1211.070 1744.160 1219.680 ;
        RECT 1928.420 1213.130 1928.680 1213.450 ;
        RECT 1743.960 1210.750 1744.220 1211.070 ;
        RECT 1928.480 20.730 1928.620 1213.130 ;
        RECT 1928.420 20.410 1928.680 20.730 ;
        RECT 1935.320 20.410 1935.580 20.730 ;
        RECT 1935.380 2.400 1935.520 20.410 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.970 1173.240 1755.290 1173.300 ;
        RECT 1758.650 1173.240 1758.970 1173.300 ;
        RECT 1754.970 1173.100 1758.970 1173.240 ;
        RECT 1754.970 1173.040 1755.290 1173.100 ;
        RECT 1758.650 1173.040 1758.970 1173.100 ;
        RECT 1758.650 22.000 1758.970 22.060 ;
        RECT 1953.230 22.000 1953.550 22.060 ;
        RECT 1758.650 21.860 1953.550 22.000 ;
        RECT 1758.650 21.800 1758.970 21.860 ;
        RECT 1953.230 21.800 1953.550 21.860 ;
      LAYER via ;
        RECT 1755.000 1173.040 1755.260 1173.300 ;
        RECT 1758.680 1173.040 1758.940 1173.300 ;
        RECT 1758.680 21.800 1758.940 22.060 ;
        RECT 1953.260 21.800 1953.520 22.060 ;
      LAYER met2 ;
        RECT 1753.170 1220.330 1753.730 1228.680 ;
        RECT 1753.170 1220.190 1755.200 1220.330 ;
        RECT 1753.170 1219.680 1753.730 1220.190 ;
        RECT 1755.060 1173.330 1755.200 1220.190 ;
        RECT 1755.000 1173.010 1755.260 1173.330 ;
        RECT 1758.680 1173.010 1758.940 1173.330 ;
        RECT 1758.740 22.090 1758.880 1173.010 ;
        RECT 1758.680 21.770 1758.940 22.090 ;
        RECT 1953.260 21.770 1953.520 22.090 ;
        RECT 1953.320 2.400 1953.460 21.770 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1762.330 1207.580 1762.650 1207.640 ;
        RECT 1766.010 1207.580 1766.330 1207.640 ;
        RECT 1762.330 1207.440 1766.330 1207.580 ;
        RECT 1762.330 1207.380 1762.650 1207.440 ;
        RECT 1766.010 1207.380 1766.330 1207.440 ;
        RECT 1766.010 23.020 1766.330 23.080 ;
        RECT 1971.170 23.020 1971.490 23.080 ;
        RECT 1766.010 22.880 1971.490 23.020 ;
        RECT 1766.010 22.820 1766.330 22.880 ;
        RECT 1971.170 22.820 1971.490 22.880 ;
      LAYER via ;
        RECT 1762.360 1207.380 1762.620 1207.640 ;
        RECT 1766.040 1207.380 1766.300 1207.640 ;
        RECT 1766.040 22.820 1766.300 23.080 ;
        RECT 1971.200 22.820 1971.460 23.080 ;
      LAYER met2 ;
        RECT 1762.370 1219.680 1762.930 1228.680 ;
        RECT 1762.420 1207.670 1762.560 1219.680 ;
        RECT 1762.360 1207.350 1762.620 1207.670 ;
        RECT 1766.040 1207.350 1766.300 1207.670 ;
        RECT 1766.100 23.110 1766.240 1207.350 ;
        RECT 1766.040 22.790 1766.300 23.110 ;
        RECT 1971.200 22.790 1971.460 23.110 ;
        RECT 1971.260 2.400 1971.400 22.790 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 23.360 1773.230 23.420 ;
        RECT 1989.110 23.360 1989.430 23.420 ;
        RECT 1772.910 23.220 1989.430 23.360 ;
        RECT 1772.910 23.160 1773.230 23.220 ;
        RECT 1989.110 23.160 1989.430 23.220 ;
      LAYER via ;
        RECT 1772.940 23.160 1773.200 23.420 ;
        RECT 1989.140 23.160 1989.400 23.420 ;
      LAYER met2 ;
        RECT 1771.570 1220.330 1772.130 1228.680 ;
        RECT 1771.570 1220.190 1773.140 1220.330 ;
        RECT 1771.570 1219.680 1772.130 1220.190 ;
        RECT 1773.000 23.450 1773.140 1220.190 ;
        RECT 1772.940 23.130 1773.200 23.450 ;
        RECT 1989.140 23.130 1989.400 23.450 ;
        RECT 1989.200 2.400 1989.340 23.130 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1786.325 786.505 1786.495 821.015 ;
        RECT 1786.325 689.605 1786.495 724.455 ;
        RECT 1786.325 593.045 1786.495 627.895 ;
        RECT 1786.325 496.485 1786.495 531.335 ;
        RECT 1786.325 386.325 1786.495 434.775 ;
        RECT 1786.325 338.045 1786.495 385.815 ;
        RECT 1786.325 241.485 1786.495 289.595 ;
        RECT 1786.325 158.525 1786.495 193.035 ;
      LAYER mcon ;
        RECT 1786.325 820.845 1786.495 821.015 ;
        RECT 1786.325 724.285 1786.495 724.455 ;
        RECT 1786.325 627.725 1786.495 627.895 ;
        RECT 1786.325 531.165 1786.495 531.335 ;
        RECT 1786.325 434.605 1786.495 434.775 ;
        RECT 1786.325 385.645 1786.495 385.815 ;
        RECT 1786.325 289.425 1786.495 289.595 ;
        RECT 1786.325 192.865 1786.495 193.035 ;
      LAYER met1 ;
        RECT 1780.730 1207.580 1781.050 1207.640 ;
        RECT 1786.710 1207.580 1787.030 1207.640 ;
        RECT 1780.730 1207.440 1787.030 1207.580 ;
        RECT 1780.730 1207.380 1781.050 1207.440 ;
        RECT 1786.710 1207.380 1787.030 1207.440 ;
        RECT 1785.790 1124.960 1786.110 1125.020 ;
        RECT 1786.710 1124.960 1787.030 1125.020 ;
        RECT 1785.790 1124.820 1787.030 1124.960 ;
        RECT 1785.790 1124.760 1786.110 1124.820 ;
        RECT 1786.710 1124.760 1787.030 1124.820 ;
        RECT 1785.790 1028.400 1786.110 1028.460 ;
        RECT 1786.710 1028.400 1787.030 1028.460 ;
        RECT 1785.790 1028.260 1787.030 1028.400 ;
        RECT 1785.790 1028.200 1786.110 1028.260 ;
        RECT 1786.710 1028.200 1787.030 1028.260 ;
        RECT 1785.790 931.840 1786.110 931.900 ;
        RECT 1786.710 931.840 1787.030 931.900 ;
        RECT 1785.790 931.700 1787.030 931.840 ;
        RECT 1785.790 931.640 1786.110 931.700 ;
        RECT 1786.710 931.640 1787.030 931.700 ;
        RECT 1785.330 869.620 1785.650 869.680 ;
        RECT 1786.710 869.620 1787.030 869.680 ;
        RECT 1785.330 869.480 1787.030 869.620 ;
        RECT 1785.330 869.420 1785.650 869.480 ;
        RECT 1786.710 869.420 1787.030 869.480 ;
        RECT 1785.790 835.280 1786.110 835.340 ;
        RECT 1786.710 835.280 1787.030 835.340 ;
        RECT 1785.790 835.140 1787.030 835.280 ;
        RECT 1785.790 835.080 1786.110 835.140 ;
        RECT 1786.710 835.080 1787.030 835.140 ;
        RECT 1786.250 821.000 1786.570 821.060 ;
        RECT 1786.055 820.860 1786.570 821.000 ;
        RECT 1786.250 820.800 1786.570 820.860 ;
        RECT 1786.250 786.660 1786.570 786.720 ;
        RECT 1786.055 786.520 1786.570 786.660 ;
        RECT 1786.250 786.460 1786.570 786.520 ;
        RECT 1785.790 738.380 1786.110 738.440 ;
        RECT 1786.710 738.380 1787.030 738.440 ;
        RECT 1785.790 738.240 1787.030 738.380 ;
        RECT 1785.790 738.180 1786.110 738.240 ;
        RECT 1786.710 738.180 1787.030 738.240 ;
        RECT 1786.250 724.440 1786.570 724.500 ;
        RECT 1786.055 724.300 1786.570 724.440 ;
        RECT 1786.250 724.240 1786.570 724.300 ;
        RECT 1786.250 689.760 1786.570 689.820 ;
        RECT 1786.055 689.620 1786.570 689.760 ;
        RECT 1786.250 689.560 1786.570 689.620 ;
        RECT 1785.790 641.820 1786.110 641.880 ;
        RECT 1786.710 641.820 1787.030 641.880 ;
        RECT 1785.790 641.680 1787.030 641.820 ;
        RECT 1785.790 641.620 1786.110 641.680 ;
        RECT 1786.710 641.620 1787.030 641.680 ;
        RECT 1786.250 627.880 1786.570 627.940 ;
        RECT 1786.055 627.740 1786.570 627.880 ;
        RECT 1786.250 627.680 1786.570 627.740 ;
        RECT 1786.250 593.200 1786.570 593.260 ;
        RECT 1786.055 593.060 1786.570 593.200 ;
        RECT 1786.250 593.000 1786.570 593.060 ;
        RECT 1785.790 545.260 1786.110 545.320 ;
        RECT 1786.710 545.260 1787.030 545.320 ;
        RECT 1785.790 545.120 1787.030 545.260 ;
        RECT 1785.790 545.060 1786.110 545.120 ;
        RECT 1786.710 545.060 1787.030 545.120 ;
        RECT 1786.250 531.320 1786.570 531.380 ;
        RECT 1786.055 531.180 1786.570 531.320 ;
        RECT 1786.250 531.120 1786.570 531.180 ;
        RECT 1786.250 496.640 1786.570 496.700 ;
        RECT 1786.055 496.500 1786.570 496.640 ;
        RECT 1786.250 496.440 1786.570 496.500 ;
        RECT 1785.790 448.700 1786.110 448.760 ;
        RECT 1786.710 448.700 1787.030 448.760 ;
        RECT 1785.790 448.560 1787.030 448.700 ;
        RECT 1785.790 448.500 1786.110 448.560 ;
        RECT 1786.710 448.500 1787.030 448.560 ;
        RECT 1786.250 434.760 1786.570 434.820 ;
        RECT 1786.055 434.620 1786.570 434.760 ;
        RECT 1786.250 434.560 1786.570 434.620 ;
        RECT 1786.265 386.480 1786.555 386.525 ;
        RECT 1786.710 386.480 1787.030 386.540 ;
        RECT 1786.265 386.340 1787.030 386.480 ;
        RECT 1786.265 386.295 1786.555 386.340 ;
        RECT 1786.710 386.280 1787.030 386.340 ;
        RECT 1786.265 385.800 1786.555 385.845 ;
        RECT 1786.710 385.800 1787.030 385.860 ;
        RECT 1786.265 385.660 1787.030 385.800 ;
        RECT 1786.265 385.615 1786.555 385.660 ;
        RECT 1786.710 385.600 1787.030 385.660 ;
        RECT 1786.250 338.200 1786.570 338.260 ;
        RECT 1786.055 338.060 1786.570 338.200 ;
        RECT 1786.250 338.000 1786.570 338.060 ;
        RECT 1786.265 289.580 1786.555 289.625 ;
        RECT 1786.710 289.580 1787.030 289.640 ;
        RECT 1786.265 289.440 1787.030 289.580 ;
        RECT 1786.265 289.395 1786.555 289.440 ;
        RECT 1786.710 289.380 1787.030 289.440 ;
        RECT 1786.250 241.640 1786.570 241.700 ;
        RECT 1786.055 241.500 1786.570 241.640 ;
        RECT 1786.250 241.440 1786.570 241.500 ;
        RECT 1786.265 193.020 1786.555 193.065 ;
        RECT 1786.710 193.020 1787.030 193.080 ;
        RECT 1786.265 192.880 1787.030 193.020 ;
        RECT 1786.265 192.835 1786.555 192.880 ;
        RECT 1786.710 192.820 1787.030 192.880 ;
        RECT 1786.250 158.680 1786.570 158.740 ;
        RECT 1786.055 158.540 1786.570 158.680 ;
        RECT 1786.250 158.480 1786.570 158.540 ;
        RECT 1785.790 22.680 1786.110 22.740 ;
        RECT 2006.590 22.680 2006.910 22.740 ;
        RECT 1785.790 22.540 2006.910 22.680 ;
        RECT 1785.790 22.480 1786.110 22.540 ;
        RECT 2006.590 22.480 2006.910 22.540 ;
      LAYER via ;
        RECT 1780.760 1207.380 1781.020 1207.640 ;
        RECT 1786.740 1207.380 1787.000 1207.640 ;
        RECT 1785.820 1124.760 1786.080 1125.020 ;
        RECT 1786.740 1124.760 1787.000 1125.020 ;
        RECT 1785.820 1028.200 1786.080 1028.460 ;
        RECT 1786.740 1028.200 1787.000 1028.460 ;
        RECT 1785.820 931.640 1786.080 931.900 ;
        RECT 1786.740 931.640 1787.000 931.900 ;
        RECT 1785.360 869.420 1785.620 869.680 ;
        RECT 1786.740 869.420 1787.000 869.680 ;
        RECT 1785.820 835.080 1786.080 835.340 ;
        RECT 1786.740 835.080 1787.000 835.340 ;
        RECT 1786.280 820.800 1786.540 821.060 ;
        RECT 1786.280 786.460 1786.540 786.720 ;
        RECT 1785.820 738.180 1786.080 738.440 ;
        RECT 1786.740 738.180 1787.000 738.440 ;
        RECT 1786.280 724.240 1786.540 724.500 ;
        RECT 1786.280 689.560 1786.540 689.820 ;
        RECT 1785.820 641.620 1786.080 641.880 ;
        RECT 1786.740 641.620 1787.000 641.880 ;
        RECT 1786.280 627.680 1786.540 627.940 ;
        RECT 1786.280 593.000 1786.540 593.260 ;
        RECT 1785.820 545.060 1786.080 545.320 ;
        RECT 1786.740 545.060 1787.000 545.320 ;
        RECT 1786.280 531.120 1786.540 531.380 ;
        RECT 1786.280 496.440 1786.540 496.700 ;
        RECT 1785.820 448.500 1786.080 448.760 ;
        RECT 1786.740 448.500 1787.000 448.760 ;
        RECT 1786.280 434.560 1786.540 434.820 ;
        RECT 1786.740 386.280 1787.000 386.540 ;
        RECT 1786.740 385.600 1787.000 385.860 ;
        RECT 1786.280 338.000 1786.540 338.260 ;
        RECT 1786.740 289.380 1787.000 289.640 ;
        RECT 1786.280 241.440 1786.540 241.700 ;
        RECT 1786.740 192.820 1787.000 193.080 ;
        RECT 1786.280 158.480 1786.540 158.740 ;
        RECT 1785.820 22.480 1786.080 22.740 ;
        RECT 2006.620 22.480 2006.880 22.740 ;
      LAYER met2 ;
        RECT 1780.770 1219.680 1781.330 1228.680 ;
        RECT 1780.820 1207.670 1780.960 1219.680 ;
        RECT 1780.760 1207.350 1781.020 1207.670 ;
        RECT 1786.740 1207.350 1787.000 1207.670 ;
        RECT 1786.800 1125.050 1786.940 1207.350 ;
        RECT 1785.820 1124.730 1786.080 1125.050 ;
        RECT 1786.740 1124.730 1787.000 1125.050 ;
        RECT 1785.880 1124.450 1786.020 1124.730 ;
        RECT 1785.880 1124.310 1786.480 1124.450 ;
        RECT 1786.340 1076.850 1786.480 1124.310 ;
        RECT 1786.340 1076.710 1786.940 1076.850 ;
        RECT 1786.800 1028.490 1786.940 1076.710 ;
        RECT 1785.820 1028.170 1786.080 1028.490 ;
        RECT 1786.740 1028.170 1787.000 1028.490 ;
        RECT 1785.880 1027.890 1786.020 1028.170 ;
        RECT 1785.880 1027.750 1786.480 1027.890 ;
        RECT 1786.340 980.290 1786.480 1027.750 ;
        RECT 1786.340 980.150 1786.940 980.290 ;
        RECT 1786.800 931.930 1786.940 980.150 ;
        RECT 1785.820 931.610 1786.080 931.930 ;
        RECT 1786.740 931.610 1787.000 931.930 ;
        RECT 1785.880 931.330 1786.020 931.610 ;
        RECT 1785.880 931.190 1786.480 931.330 ;
        RECT 1786.340 917.845 1786.480 931.190 ;
        RECT 1785.350 917.475 1785.630 917.845 ;
        RECT 1786.270 917.475 1786.550 917.845 ;
        RECT 1785.420 869.710 1785.560 917.475 ;
        RECT 1785.360 869.390 1785.620 869.710 ;
        RECT 1786.740 869.390 1787.000 869.710 ;
        RECT 1786.800 835.370 1786.940 869.390 ;
        RECT 1785.820 835.050 1786.080 835.370 ;
        RECT 1786.740 835.050 1787.000 835.370 ;
        RECT 1785.880 834.770 1786.020 835.050 ;
        RECT 1785.880 834.630 1786.480 834.770 ;
        RECT 1786.340 821.090 1786.480 834.630 ;
        RECT 1786.280 820.770 1786.540 821.090 ;
        RECT 1786.280 786.430 1786.540 786.750 ;
        RECT 1786.340 772.890 1786.480 786.430 ;
        RECT 1786.340 772.750 1786.940 772.890 ;
        RECT 1786.800 738.470 1786.940 772.750 ;
        RECT 1785.820 738.210 1786.080 738.470 ;
        RECT 1785.820 738.150 1786.480 738.210 ;
        RECT 1786.740 738.150 1787.000 738.470 ;
        RECT 1785.880 738.070 1786.480 738.150 ;
        RECT 1786.340 724.530 1786.480 738.070 ;
        RECT 1786.280 724.210 1786.540 724.530 ;
        RECT 1786.280 689.530 1786.540 689.850 ;
        RECT 1786.340 676.330 1786.480 689.530 ;
        RECT 1786.340 676.190 1786.940 676.330 ;
        RECT 1786.800 641.910 1786.940 676.190 ;
        RECT 1785.820 641.650 1786.080 641.910 ;
        RECT 1785.820 641.590 1786.480 641.650 ;
        RECT 1786.740 641.590 1787.000 641.910 ;
        RECT 1785.880 641.510 1786.480 641.590 ;
        RECT 1786.340 627.970 1786.480 641.510 ;
        RECT 1786.280 627.650 1786.540 627.970 ;
        RECT 1786.280 592.970 1786.540 593.290 ;
        RECT 1786.340 579.770 1786.480 592.970 ;
        RECT 1786.340 579.630 1786.940 579.770 ;
        RECT 1786.800 545.350 1786.940 579.630 ;
        RECT 1785.820 545.090 1786.080 545.350 ;
        RECT 1785.820 545.030 1786.480 545.090 ;
        RECT 1786.740 545.030 1787.000 545.350 ;
        RECT 1785.880 544.950 1786.480 545.030 ;
        RECT 1786.340 531.410 1786.480 544.950 ;
        RECT 1786.280 531.090 1786.540 531.410 ;
        RECT 1786.280 496.410 1786.540 496.730 ;
        RECT 1786.340 483.210 1786.480 496.410 ;
        RECT 1786.340 483.070 1786.940 483.210 ;
        RECT 1786.800 448.790 1786.940 483.070 ;
        RECT 1785.820 448.530 1786.080 448.790 ;
        RECT 1785.820 448.470 1786.480 448.530 ;
        RECT 1786.740 448.470 1787.000 448.790 ;
        RECT 1785.880 448.390 1786.480 448.470 ;
        RECT 1786.340 434.850 1786.480 448.390 ;
        RECT 1786.280 434.530 1786.540 434.850 ;
        RECT 1786.740 386.250 1787.000 386.570 ;
        RECT 1786.800 385.890 1786.940 386.250 ;
        RECT 1786.740 385.570 1787.000 385.890 ;
        RECT 1786.280 337.970 1786.540 338.290 ;
        RECT 1786.340 303.690 1786.480 337.970 ;
        RECT 1786.340 303.550 1786.940 303.690 ;
        RECT 1786.800 289.670 1786.940 303.550 ;
        RECT 1786.740 289.350 1787.000 289.670 ;
        RECT 1786.280 241.410 1786.540 241.730 ;
        RECT 1786.340 207.130 1786.480 241.410 ;
        RECT 1786.340 206.990 1786.940 207.130 ;
        RECT 1786.800 193.110 1786.940 206.990 ;
        RECT 1786.740 192.790 1787.000 193.110 ;
        RECT 1786.280 158.450 1786.540 158.770 ;
        RECT 1786.340 110.570 1786.480 158.450 ;
        RECT 1786.340 110.430 1786.940 110.570 ;
        RECT 1786.800 62.290 1786.940 110.430 ;
        RECT 1785.880 62.150 1786.940 62.290 ;
        RECT 1785.880 22.770 1786.020 62.150 ;
        RECT 1785.820 22.450 1786.080 22.770 ;
        RECT 2006.620 22.450 2006.880 22.770 ;
        RECT 2006.680 2.400 2006.820 22.450 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
      LAYER via2 ;
        RECT 1785.350 917.520 1785.630 917.800 ;
        RECT 1786.270 917.520 1786.550 917.800 ;
      LAYER met3 ;
        RECT 1785.325 917.810 1785.655 917.825 ;
        RECT 1786.245 917.810 1786.575 917.825 ;
        RECT 1785.325 917.510 1786.575 917.810 ;
        RECT 1785.325 917.495 1785.655 917.510 ;
        RECT 1786.245 917.495 1786.575 917.510 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1789.930 1207.580 1790.250 1207.640 ;
        RECT 1793.610 1207.580 1793.930 1207.640 ;
        RECT 1789.930 1207.440 1793.930 1207.580 ;
        RECT 1789.930 1207.380 1790.250 1207.440 ;
        RECT 1793.610 1207.380 1793.930 1207.440 ;
        RECT 2024.530 24.040 2024.850 24.100 ;
        RECT 2001.620 23.900 2024.850 24.040 ;
        RECT 1793.610 23.700 1793.930 23.760 ;
        RECT 2001.620 23.700 2001.760 23.900 ;
        RECT 2024.530 23.840 2024.850 23.900 ;
        RECT 1793.610 23.560 2001.760 23.700 ;
        RECT 1793.610 23.500 1793.930 23.560 ;
      LAYER via ;
        RECT 1789.960 1207.380 1790.220 1207.640 ;
        RECT 1793.640 1207.380 1793.900 1207.640 ;
        RECT 1793.640 23.500 1793.900 23.760 ;
        RECT 2024.560 23.840 2024.820 24.100 ;
      LAYER met2 ;
        RECT 1789.970 1219.680 1790.530 1228.680 ;
        RECT 1790.020 1207.670 1790.160 1219.680 ;
        RECT 1789.960 1207.350 1790.220 1207.670 ;
        RECT 1793.640 1207.350 1793.900 1207.670 ;
        RECT 1793.700 23.790 1793.840 1207.350 ;
        RECT 2024.560 23.810 2024.820 24.130 ;
        RECT 1793.640 23.470 1793.900 23.790 ;
        RECT 2024.620 2.400 2024.760 23.810 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.050 27.100 1800.370 27.160 ;
        RECT 2042.470 27.100 2042.790 27.160 ;
        RECT 1800.050 26.960 2042.790 27.100 ;
        RECT 1800.050 26.900 1800.370 26.960 ;
        RECT 2042.470 26.900 2042.790 26.960 ;
      LAYER via ;
        RECT 1800.080 26.900 1800.340 27.160 ;
        RECT 2042.500 26.900 2042.760 27.160 ;
      LAYER met2 ;
        RECT 1799.170 1220.330 1799.730 1228.680 ;
        RECT 1799.170 1220.190 1800.280 1220.330 ;
        RECT 1799.170 1219.680 1799.730 1220.190 ;
        RECT 1800.140 27.190 1800.280 1220.190 ;
        RECT 1800.080 26.870 1800.340 27.190 ;
        RECT 2042.500 26.870 2042.760 27.190 ;
        RECT 2042.560 2.400 2042.700 26.870 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 757.690 24.040 758.010 24.100 ;
        RECT 1139.490 24.040 1139.810 24.100 ;
        RECT 757.690 23.900 1139.810 24.040 ;
        RECT 757.690 23.840 758.010 23.900 ;
        RECT 1139.490 23.840 1139.810 23.900 ;
      LAYER via ;
        RECT 757.720 23.840 757.980 24.100 ;
        RECT 1139.520 23.840 1139.780 24.100 ;
      LAYER met2 ;
        RECT 1139.070 1220.330 1139.630 1228.680 ;
        RECT 1139.070 1219.680 1139.720 1220.330 ;
        RECT 1139.580 24.130 1139.720 1219.680 ;
        RECT 757.720 23.810 757.980 24.130 ;
        RECT 1139.520 23.810 1139.780 24.130 ;
        RECT 757.780 2.400 757.920 23.810 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.870 1207.580 1808.190 1207.640 ;
        RECT 1813.850 1207.580 1814.170 1207.640 ;
        RECT 1807.870 1207.440 1814.170 1207.580 ;
        RECT 1807.870 1207.380 1808.190 1207.440 ;
        RECT 1813.850 1207.380 1814.170 1207.440 ;
        RECT 1813.850 27.440 1814.170 27.500 ;
        RECT 2060.410 27.440 2060.730 27.500 ;
        RECT 1813.850 27.300 2060.730 27.440 ;
        RECT 1813.850 27.240 1814.170 27.300 ;
        RECT 2060.410 27.240 2060.730 27.300 ;
      LAYER via ;
        RECT 1807.900 1207.380 1808.160 1207.640 ;
        RECT 1813.880 1207.380 1814.140 1207.640 ;
        RECT 1813.880 27.240 1814.140 27.500 ;
        RECT 2060.440 27.240 2060.700 27.500 ;
      LAYER met2 ;
        RECT 1807.910 1219.680 1808.470 1228.680 ;
        RECT 1807.960 1207.670 1808.100 1219.680 ;
        RECT 1807.900 1207.350 1808.160 1207.670 ;
        RECT 1813.880 1207.350 1814.140 1207.670 ;
        RECT 1813.940 27.530 1814.080 1207.350 ;
        RECT 1813.880 27.210 1814.140 27.530 ;
        RECT 2060.440 27.210 2060.700 27.530 ;
        RECT 2060.500 2.400 2060.640 27.210 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1817.070 1207.580 1817.390 1207.640 ;
        RECT 1821.210 1207.580 1821.530 1207.640 ;
        RECT 1817.070 1207.440 1821.530 1207.580 ;
        RECT 1817.070 1207.380 1817.390 1207.440 ;
        RECT 1821.210 1207.380 1821.530 1207.440 ;
        RECT 1821.210 26.760 1821.530 26.820 ;
        RECT 2078.350 26.760 2078.670 26.820 ;
        RECT 1821.210 26.620 2078.670 26.760 ;
        RECT 1821.210 26.560 1821.530 26.620 ;
        RECT 2078.350 26.560 2078.670 26.620 ;
      LAYER via ;
        RECT 1817.100 1207.380 1817.360 1207.640 ;
        RECT 1821.240 1207.380 1821.500 1207.640 ;
        RECT 1821.240 26.560 1821.500 26.820 ;
        RECT 2078.380 26.560 2078.640 26.820 ;
      LAYER met2 ;
        RECT 1817.110 1219.680 1817.670 1228.680 ;
        RECT 1817.160 1207.670 1817.300 1219.680 ;
        RECT 1817.100 1207.350 1817.360 1207.670 ;
        RECT 1821.240 1207.350 1821.500 1207.670 ;
        RECT 1821.300 26.850 1821.440 1207.350 ;
        RECT 1821.240 26.530 1821.500 26.850 ;
        RECT 2078.380 26.530 2078.640 26.850 ;
        RECT 2078.440 2.400 2078.580 26.530 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.110 26.420 1828.430 26.480 ;
        RECT 2095.830 26.420 2096.150 26.480 ;
        RECT 1828.110 26.280 2096.150 26.420 ;
        RECT 1828.110 26.220 1828.430 26.280 ;
        RECT 2095.830 26.220 2096.150 26.280 ;
      LAYER via ;
        RECT 1828.140 26.220 1828.400 26.480 ;
        RECT 2095.860 26.220 2096.120 26.480 ;
      LAYER met2 ;
        RECT 1826.310 1220.330 1826.870 1228.680 ;
        RECT 1826.310 1220.190 1828.340 1220.330 ;
        RECT 1826.310 1219.680 1826.870 1220.190 ;
        RECT 1828.200 26.510 1828.340 1220.190 ;
        RECT 1828.140 26.190 1828.400 26.510 ;
        RECT 2095.860 26.190 2096.120 26.510 ;
        RECT 2095.920 2.400 2096.060 26.190 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1836.850 1208.940 1837.170 1209.000 ;
        RECT 1841.910 1208.940 1842.230 1209.000 ;
        RECT 1836.850 1208.800 1842.230 1208.940 ;
        RECT 1836.850 1208.740 1837.170 1208.800 ;
        RECT 1841.910 1208.740 1842.230 1208.800 ;
        RECT 1841.910 26.080 1842.230 26.140 ;
        RECT 2113.770 26.080 2114.090 26.140 ;
        RECT 1841.910 25.940 2114.090 26.080 ;
        RECT 1841.910 25.880 1842.230 25.940 ;
        RECT 2113.770 25.880 2114.090 25.940 ;
      LAYER via ;
        RECT 1836.880 1208.740 1837.140 1209.000 ;
        RECT 1841.940 1208.740 1842.200 1209.000 ;
        RECT 1841.940 25.880 1842.200 26.140 ;
        RECT 2113.800 25.880 2114.060 26.140 ;
      LAYER met2 ;
        RECT 1835.510 1220.330 1836.070 1228.680 ;
        RECT 1835.510 1220.190 1837.080 1220.330 ;
        RECT 1835.510 1219.680 1836.070 1220.190 ;
        RECT 1836.940 1209.030 1837.080 1220.190 ;
        RECT 1836.880 1208.710 1837.140 1209.030 ;
        RECT 1841.940 1208.710 1842.200 1209.030 ;
        RECT 1842.000 26.170 1842.140 1208.710 ;
        RECT 1841.940 25.850 1842.200 26.170 ;
        RECT 2113.800 25.850 2114.060 26.170 ;
        RECT 2113.860 2.400 2114.000 25.850 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2111.085 22.525 2111.255 25.755 ;
      LAYER mcon ;
        RECT 2111.085 25.585 2111.255 25.755 ;
      LAYER met1 ;
        RECT 1844.670 1215.400 1844.990 1215.460 ;
        RECT 1848.810 1215.400 1849.130 1215.460 ;
        RECT 1844.670 1215.260 1849.130 1215.400 ;
        RECT 1844.670 1215.200 1844.990 1215.260 ;
        RECT 1848.810 1215.200 1849.130 1215.260 ;
        RECT 1848.810 25.740 1849.130 25.800 ;
        RECT 2111.025 25.740 2111.315 25.785 ;
        RECT 1848.810 25.600 2111.315 25.740 ;
        RECT 1848.810 25.540 1849.130 25.600 ;
        RECT 2111.025 25.555 2111.315 25.600 ;
        RECT 2111.025 22.680 2111.315 22.725 ;
        RECT 2131.710 22.680 2132.030 22.740 ;
        RECT 2111.025 22.540 2132.030 22.680 ;
        RECT 2111.025 22.495 2111.315 22.540 ;
        RECT 2131.710 22.480 2132.030 22.540 ;
      LAYER via ;
        RECT 1844.700 1215.200 1844.960 1215.460 ;
        RECT 1848.840 1215.200 1849.100 1215.460 ;
        RECT 1848.840 25.540 1849.100 25.800 ;
        RECT 2131.740 22.480 2132.000 22.740 ;
      LAYER met2 ;
        RECT 1844.710 1219.680 1845.270 1228.680 ;
        RECT 1844.760 1215.490 1844.900 1219.680 ;
        RECT 1844.700 1215.170 1844.960 1215.490 ;
        RECT 1848.840 1215.170 1849.100 1215.490 ;
        RECT 1848.900 25.830 1849.040 1215.170 ;
        RECT 1848.840 25.510 1849.100 25.830 ;
        RECT 2131.740 22.450 2132.000 22.770 ;
        RECT 2131.800 2.400 2131.940 22.450 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2017.705 22.525 2017.875 25.415 ;
        RECT 2062.785 22.525 2062.955 25.415 ;
      LAYER mcon ;
        RECT 2017.705 25.245 2017.875 25.415 ;
        RECT 2062.785 25.245 2062.955 25.415 ;
      LAYER met1 ;
        RECT 2120.670 27.100 2120.990 27.160 ;
        RECT 2149.650 27.100 2149.970 27.160 ;
        RECT 2120.670 26.960 2149.970 27.100 ;
        RECT 2120.670 26.900 2120.990 26.960 ;
        RECT 2149.650 26.900 2149.970 26.960 ;
        RECT 1855.250 25.400 1855.570 25.460 ;
        RECT 2017.645 25.400 2017.935 25.445 ;
        RECT 1855.250 25.260 2017.935 25.400 ;
        RECT 1855.250 25.200 1855.570 25.260 ;
        RECT 2017.645 25.215 2017.935 25.260 ;
        RECT 2062.725 25.400 2063.015 25.445 ;
        RECT 2100.430 25.400 2100.750 25.460 ;
        RECT 2062.725 25.260 2100.750 25.400 ;
        RECT 2062.725 25.215 2063.015 25.260 ;
        RECT 2100.430 25.200 2100.750 25.260 ;
        RECT 2017.645 22.680 2017.935 22.725 ;
        RECT 2062.725 22.680 2063.015 22.725 ;
        RECT 2017.645 22.540 2063.015 22.680 ;
        RECT 2017.645 22.495 2017.935 22.540 ;
        RECT 2062.725 22.495 2063.015 22.540 ;
      LAYER via ;
        RECT 2120.700 26.900 2120.960 27.160 ;
        RECT 2149.680 26.900 2149.940 27.160 ;
        RECT 1855.280 25.200 1855.540 25.460 ;
        RECT 2100.460 25.200 2100.720 25.460 ;
      LAYER met2 ;
        RECT 1853.910 1220.330 1854.470 1228.680 ;
        RECT 1853.910 1220.190 1855.480 1220.330 ;
        RECT 1853.910 1219.680 1854.470 1220.190 ;
        RECT 1855.340 25.490 1855.480 1220.190 ;
        RECT 2120.700 26.870 2120.960 27.190 ;
        RECT 2149.680 26.870 2149.940 27.190 ;
        RECT 2120.760 26.365 2120.900 26.870 ;
        RECT 2100.450 25.995 2100.730 26.365 ;
        RECT 2120.690 25.995 2120.970 26.365 ;
        RECT 2100.520 25.490 2100.660 25.995 ;
        RECT 1855.280 25.170 1855.540 25.490 ;
        RECT 2100.460 25.170 2100.720 25.490 ;
        RECT 2149.740 2.400 2149.880 26.870 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
      LAYER via2 ;
        RECT 2100.450 26.040 2100.730 26.320 ;
        RECT 2120.690 26.040 2120.970 26.320 ;
      LAYER met3 ;
        RECT 2100.425 26.330 2100.755 26.345 ;
        RECT 2120.665 26.330 2120.995 26.345 ;
        RECT 2100.425 26.030 2120.995 26.330 ;
        RECT 2100.425 26.015 2100.755 26.030 ;
        RECT 2120.665 26.015 2120.995 26.030 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1863.070 1207.580 1863.390 1207.640 ;
        RECT 1869.050 1207.580 1869.370 1207.640 ;
        RECT 1863.070 1207.440 1869.370 1207.580 ;
        RECT 1863.070 1207.380 1863.390 1207.440 ;
        RECT 1869.050 1207.380 1869.370 1207.440 ;
        RECT 2115.700 26.280 2163.680 26.420 ;
        RECT 2115.700 25.740 2115.840 26.280 ;
        RECT 2115.240 25.600 2115.840 25.740 ;
        RECT 2163.540 25.740 2163.680 26.280 ;
        RECT 2167.590 25.740 2167.910 25.800 ;
        RECT 2163.540 25.600 2167.910 25.740 ;
        RECT 2018.090 25.400 2018.410 25.460 ;
        RECT 2018.090 25.260 2062.480 25.400 ;
        RECT 2018.090 25.200 2018.410 25.260 ;
        RECT 1869.050 25.060 1869.370 25.120 ;
        RECT 1896.650 25.060 1896.970 25.120 ;
        RECT 1869.050 24.920 1896.970 25.060 ;
        RECT 1869.050 24.860 1869.370 24.920 ;
        RECT 1896.650 24.860 1896.970 24.920 ;
        RECT 1897.570 25.060 1897.890 25.120 ;
        RECT 1993.710 25.060 1994.030 25.120 ;
        RECT 1897.570 24.920 1994.030 25.060 ;
        RECT 2062.340 25.060 2062.480 25.260 ;
        RECT 2115.240 25.060 2115.380 25.600 ;
        RECT 2167.590 25.540 2167.910 25.600 ;
        RECT 2062.340 24.920 2115.380 25.060 ;
        RECT 1897.570 24.860 1897.890 24.920 ;
        RECT 1993.710 24.860 1994.030 24.920 ;
      LAYER via ;
        RECT 1863.100 1207.380 1863.360 1207.640 ;
        RECT 1869.080 1207.380 1869.340 1207.640 ;
        RECT 2018.120 25.200 2018.380 25.460 ;
        RECT 1869.080 24.860 1869.340 25.120 ;
        RECT 1896.680 24.860 1896.940 25.120 ;
        RECT 1897.600 24.860 1897.860 25.120 ;
        RECT 1993.740 24.860 1994.000 25.120 ;
        RECT 2167.620 25.540 2167.880 25.800 ;
      LAYER met2 ;
        RECT 1863.110 1219.680 1863.670 1228.680 ;
        RECT 1863.160 1207.670 1863.300 1219.680 ;
        RECT 1863.100 1207.350 1863.360 1207.670 ;
        RECT 1869.080 1207.350 1869.340 1207.670 ;
        RECT 1869.140 25.150 1869.280 1207.350 ;
        RECT 2167.620 25.510 2167.880 25.830 ;
        RECT 2018.120 25.170 2018.380 25.490 ;
        RECT 1869.080 24.830 1869.340 25.150 ;
        RECT 1896.680 25.005 1896.940 25.150 ;
        RECT 1897.600 25.005 1897.860 25.150 ;
        RECT 1993.740 25.005 1994.000 25.150 ;
        RECT 2018.180 25.005 2018.320 25.170 ;
        RECT 1896.670 24.635 1896.950 25.005 ;
        RECT 1897.590 24.635 1897.870 25.005 ;
        RECT 1993.730 24.635 1994.010 25.005 ;
        RECT 2018.110 24.635 2018.390 25.005 ;
        RECT 2167.680 2.400 2167.820 25.510 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
      LAYER via2 ;
        RECT 1896.670 24.680 1896.950 24.960 ;
        RECT 1897.590 24.680 1897.870 24.960 ;
        RECT 1993.730 24.680 1994.010 24.960 ;
        RECT 2018.110 24.680 2018.390 24.960 ;
      LAYER met3 ;
        RECT 1896.645 24.970 1896.975 24.985 ;
        RECT 1897.565 24.970 1897.895 24.985 ;
        RECT 1896.645 24.670 1897.895 24.970 ;
        RECT 1896.645 24.655 1896.975 24.670 ;
        RECT 1897.565 24.655 1897.895 24.670 ;
        RECT 1993.705 24.970 1994.035 24.985 ;
        RECT 2018.085 24.970 2018.415 24.985 ;
        RECT 1993.705 24.670 2018.415 24.970 ;
        RECT 1993.705 24.655 1994.035 24.670 ;
        RECT 2018.085 24.655 2018.415 24.670 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1872.270 1207.580 1872.590 1207.640 ;
        RECT 1876.410 1207.580 1876.730 1207.640 ;
        RECT 1872.270 1207.440 1876.730 1207.580 ;
        RECT 1872.270 1207.380 1872.590 1207.440 ;
        RECT 1876.410 1207.380 1876.730 1207.440 ;
        RECT 2163.450 25.060 2163.770 25.120 ;
        RECT 2185.070 25.060 2185.390 25.120 ;
        RECT 2163.450 24.920 2185.390 25.060 ;
        RECT 2163.450 24.860 2163.770 24.920 ;
        RECT 2185.070 24.860 2185.390 24.920 ;
        RECT 1876.410 24.720 1876.730 24.780 ;
        RECT 1876.410 24.580 2115.380 24.720 ;
        RECT 1876.410 24.520 1876.730 24.580 ;
        RECT 2115.240 24.380 2115.380 24.580 ;
        RECT 2162.070 24.380 2162.390 24.440 ;
        RECT 2115.240 24.240 2162.390 24.380 ;
        RECT 2162.070 24.180 2162.390 24.240 ;
      LAYER via ;
        RECT 1872.300 1207.380 1872.560 1207.640 ;
        RECT 1876.440 1207.380 1876.700 1207.640 ;
        RECT 2163.480 24.860 2163.740 25.120 ;
        RECT 2185.100 24.860 2185.360 25.120 ;
        RECT 1876.440 24.520 1876.700 24.780 ;
        RECT 2162.100 24.180 2162.360 24.440 ;
      LAYER met2 ;
        RECT 1872.310 1219.680 1872.870 1228.680 ;
        RECT 1872.360 1207.670 1872.500 1219.680 ;
        RECT 1872.300 1207.350 1872.560 1207.670 ;
        RECT 1876.440 1207.350 1876.700 1207.670 ;
        RECT 1876.500 24.810 1876.640 1207.350 ;
        RECT 2163.480 24.890 2163.740 25.150 ;
        RECT 2162.160 24.830 2163.740 24.890 ;
        RECT 2185.100 24.830 2185.360 25.150 ;
        RECT 1876.440 24.490 1876.700 24.810 ;
        RECT 2162.160 24.750 2163.680 24.830 ;
        RECT 2162.160 24.470 2162.300 24.750 ;
        RECT 2162.100 24.150 2162.360 24.470 ;
        RECT 2185.160 2.400 2185.300 24.830 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2001.145 23.715 2001.315 24.055 ;
        RECT 2115.685 23.885 2115.855 25.075 ;
        RECT 2001.145 23.545 2002.235 23.715 ;
      LAYER mcon ;
        RECT 2115.685 24.905 2115.855 25.075 ;
        RECT 2001.145 23.885 2001.315 24.055 ;
        RECT 2002.065 23.545 2002.235 23.715 ;
      LAYER met1 ;
        RECT 2115.700 25.260 2163.220 25.400 ;
        RECT 2115.700 25.105 2115.840 25.260 ;
        RECT 2115.625 24.875 2115.915 25.105 ;
        RECT 2163.080 24.720 2163.220 25.260 ;
        RECT 2203.010 24.720 2203.330 24.780 ;
        RECT 2163.080 24.580 2203.330 24.720 ;
        RECT 2203.010 24.520 2203.330 24.580 ;
        RECT 1883.310 24.040 1883.630 24.100 ;
        RECT 2001.085 24.040 2001.375 24.085 ;
        RECT 2115.625 24.040 2115.915 24.085 ;
        RECT 1883.310 23.900 2001.375 24.040 ;
        RECT 1883.310 23.840 1883.630 23.900 ;
        RECT 2001.085 23.855 2001.375 23.900 ;
        RECT 2087.180 23.900 2115.915 24.040 ;
        RECT 2002.005 23.700 2002.295 23.745 ;
        RECT 2087.180 23.700 2087.320 23.900 ;
        RECT 2115.625 23.855 2115.915 23.900 ;
        RECT 2002.005 23.560 2087.320 23.700 ;
        RECT 2002.005 23.515 2002.295 23.560 ;
      LAYER via ;
        RECT 2203.040 24.520 2203.300 24.780 ;
        RECT 1883.340 23.840 1883.600 24.100 ;
      LAYER met2 ;
        RECT 1881.510 1220.330 1882.070 1228.680 ;
        RECT 1881.510 1220.190 1883.540 1220.330 ;
        RECT 1881.510 1219.680 1882.070 1220.190 ;
        RECT 1883.400 24.130 1883.540 1220.190 ;
        RECT 2203.040 24.490 2203.300 24.810 ;
        RECT 1883.340 23.810 1883.600 24.130 ;
        RECT 2203.100 2.400 2203.240 24.490 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2114.765 24.225 2114.935 27.455 ;
        RECT 2208.145 25.245 2209.695 25.415 ;
        RECT 2209.525 24.225 2209.695 25.245 ;
      LAYER mcon ;
        RECT 2114.765 27.285 2114.935 27.455 ;
      LAYER met1 ;
        RECT 1890.670 1213.700 1890.990 1213.760 ;
        RECT 1897.110 1213.700 1897.430 1213.760 ;
        RECT 1890.670 1213.560 1897.430 1213.700 ;
        RECT 1890.670 1213.500 1890.990 1213.560 ;
        RECT 1897.110 1213.500 1897.430 1213.560 ;
        RECT 2114.705 27.440 2114.995 27.485 ;
        RECT 2114.705 27.300 2162.760 27.440 ;
        RECT 2114.705 27.255 2114.995 27.300 ;
        RECT 2162.620 27.100 2162.760 27.300 ;
        RECT 2163.910 27.100 2164.230 27.160 ;
        RECT 2162.620 26.960 2164.230 27.100 ;
        RECT 2163.910 26.900 2164.230 26.960 ;
        RECT 2163.910 25.400 2164.230 25.460 ;
        RECT 2208.085 25.400 2208.375 25.445 ;
        RECT 2163.910 25.260 2208.375 25.400 ;
        RECT 2163.910 25.200 2164.230 25.260 ;
        RECT 2208.085 25.215 2208.375 25.260 ;
        RECT 1897.110 24.380 1897.430 24.440 ;
        RECT 1994.170 24.380 1994.490 24.440 ;
        RECT 2114.705 24.380 2114.995 24.425 ;
        RECT 1897.110 24.240 1994.490 24.380 ;
        RECT 1897.110 24.180 1897.430 24.240 ;
        RECT 1994.170 24.180 1994.490 24.240 ;
        RECT 2062.800 24.240 2114.995 24.380 ;
        RECT 2024.990 24.040 2025.310 24.100 ;
        RECT 2062.800 24.040 2062.940 24.240 ;
        RECT 2114.705 24.195 2114.995 24.240 ;
        RECT 2209.465 24.380 2209.755 24.425 ;
        RECT 2220.950 24.380 2221.270 24.440 ;
        RECT 2209.465 24.240 2221.270 24.380 ;
        RECT 2209.465 24.195 2209.755 24.240 ;
        RECT 2220.950 24.180 2221.270 24.240 ;
        RECT 2024.990 23.900 2062.940 24.040 ;
        RECT 2024.990 23.840 2025.310 23.900 ;
      LAYER via ;
        RECT 1890.700 1213.500 1890.960 1213.760 ;
        RECT 1897.140 1213.500 1897.400 1213.760 ;
        RECT 2163.940 26.900 2164.200 27.160 ;
        RECT 2163.940 25.200 2164.200 25.460 ;
        RECT 1897.140 24.180 1897.400 24.440 ;
        RECT 1994.200 24.180 1994.460 24.440 ;
        RECT 2025.020 23.840 2025.280 24.100 ;
        RECT 2220.980 24.180 2221.240 24.440 ;
      LAYER met2 ;
        RECT 1890.710 1219.680 1891.270 1228.680 ;
        RECT 1890.760 1213.790 1890.900 1219.680 ;
        RECT 1890.700 1213.470 1890.960 1213.790 ;
        RECT 1897.140 1213.470 1897.400 1213.790 ;
        RECT 1897.200 24.470 1897.340 1213.470 ;
        RECT 2163.940 26.870 2164.200 27.190 ;
        RECT 2164.000 25.490 2164.140 26.870 ;
        RECT 2163.940 25.170 2164.200 25.490 ;
        RECT 1897.140 24.150 1897.400 24.470 ;
        RECT 1994.200 24.210 1994.460 24.470 ;
        RECT 1994.200 24.150 1994.860 24.210 ;
        RECT 2220.980 24.150 2221.240 24.470 ;
        RECT 1994.260 24.070 1994.860 24.150 ;
        RECT 1994.720 23.645 1994.860 24.070 ;
        RECT 2025.020 23.810 2025.280 24.130 ;
        RECT 2025.080 23.645 2025.220 23.810 ;
        RECT 1994.650 23.275 1994.930 23.645 ;
        RECT 2025.010 23.275 2025.290 23.645 ;
        RECT 2221.040 2.400 2221.180 24.150 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
      LAYER via2 ;
        RECT 1994.650 23.320 1994.930 23.600 ;
        RECT 2025.010 23.320 2025.290 23.600 ;
      LAYER met3 ;
        RECT 1994.625 23.610 1994.955 23.625 ;
        RECT 2024.985 23.610 2025.315 23.625 ;
        RECT 1994.625 23.310 2025.315 23.610 ;
        RECT 1994.625 23.295 1994.955 23.310 ;
        RECT 2024.985 23.295 2025.315 23.310 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 776.090 24.720 776.410 24.780 ;
        RECT 1145.470 24.720 1145.790 24.780 ;
        RECT 776.090 24.580 1145.790 24.720 ;
        RECT 776.090 24.520 776.410 24.580 ;
        RECT 1145.470 24.520 1145.790 24.580 ;
      LAYER via ;
        RECT 776.120 24.520 776.380 24.780 ;
        RECT 1145.500 24.520 1145.760 24.780 ;
      LAYER met2 ;
        RECT 1148.270 1221.010 1148.830 1228.680 ;
        RECT 1146.020 1220.870 1148.830 1221.010 ;
        RECT 1146.020 1196.530 1146.160 1220.870 ;
        RECT 1148.270 1219.680 1148.830 1220.870 ;
        RECT 1145.560 1196.390 1146.160 1196.530 ;
        RECT 1145.560 24.810 1145.700 1196.390 ;
        RECT 776.120 24.490 776.380 24.810 ;
        RECT 1145.500 24.490 1145.760 24.810 ;
        RECT 776.180 12.650 776.320 24.490 ;
        RECT 775.720 12.510 776.320 12.650 ;
        RECT 775.720 2.400 775.860 12.510 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.870 1207.580 1900.190 1207.640 ;
        RECT 1904.010 1207.580 1904.330 1207.640 ;
        RECT 1899.870 1207.440 1904.330 1207.580 ;
        RECT 1899.870 1207.380 1900.190 1207.440 ;
        RECT 1904.010 1207.380 1904.330 1207.440 ;
      LAYER via ;
        RECT 1899.900 1207.380 1900.160 1207.640 ;
        RECT 1904.040 1207.380 1904.300 1207.640 ;
      LAYER met2 ;
        RECT 1899.910 1219.680 1900.470 1228.680 ;
        RECT 1899.960 1207.670 1900.100 1219.680 ;
        RECT 1899.900 1207.350 1900.160 1207.670 ;
        RECT 1904.040 1207.350 1904.300 1207.670 ;
        RECT 1904.100 24.325 1904.240 1207.350 ;
        RECT 1904.030 23.955 1904.310 24.325 ;
        RECT 2238.910 23.955 2239.190 24.325 ;
        RECT 2238.980 2.400 2239.120 23.955 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
      LAYER via2 ;
        RECT 1904.030 24.000 1904.310 24.280 ;
        RECT 2238.910 24.000 2239.190 24.280 ;
      LAYER met3 ;
        RECT 1904.005 24.290 1904.335 24.305 ;
        RECT 2238.885 24.290 2239.215 24.305 ;
        RECT 1904.005 23.990 2239.215 24.290 ;
        RECT 1904.005 23.975 1904.335 23.990 ;
        RECT 2238.885 23.975 2239.215 23.990 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1923.880 21.180 1942.420 21.320 ;
        RECT 1910.910 20.980 1911.230 21.040 ;
        RECT 1910.910 20.840 1922.180 20.980 ;
        RECT 1910.910 20.780 1911.230 20.840 ;
        RECT 1922.040 20.640 1922.180 20.840 ;
        RECT 1923.880 20.640 1924.020 21.180 ;
        RECT 1942.280 20.980 1942.420 21.180 ;
        RECT 2256.370 20.980 2256.690 21.040 ;
        RECT 1942.280 20.840 2256.690 20.980 ;
        RECT 2256.370 20.780 2256.690 20.840 ;
        RECT 1922.040 20.500 1924.020 20.640 ;
      LAYER via ;
        RECT 1910.940 20.780 1911.200 21.040 ;
        RECT 2256.400 20.780 2256.660 21.040 ;
      LAYER met2 ;
        RECT 1909.110 1220.330 1909.670 1228.680 ;
        RECT 1909.110 1220.190 1911.140 1220.330 ;
        RECT 1909.110 1219.680 1909.670 1220.190 ;
        RECT 1911.000 21.070 1911.140 1220.190 ;
        RECT 1910.940 20.750 1911.200 21.070 ;
        RECT 2256.400 20.750 2256.660 21.070 ;
        RECT 2256.460 2.400 2256.600 20.750 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1918.270 1207.580 1918.590 1207.640 ;
        RECT 1924.710 1207.580 1925.030 1207.640 ;
        RECT 1918.270 1207.440 1925.030 1207.580 ;
        RECT 1918.270 1207.380 1918.590 1207.440 ;
        RECT 1924.710 1207.380 1925.030 1207.440 ;
        RECT 1924.710 27.780 1925.030 27.840 ;
        RECT 2274.310 27.780 2274.630 27.840 ;
        RECT 1924.710 27.640 2274.630 27.780 ;
        RECT 1924.710 27.580 1925.030 27.640 ;
        RECT 2274.310 27.580 2274.630 27.640 ;
      LAYER via ;
        RECT 1918.300 1207.380 1918.560 1207.640 ;
        RECT 1924.740 1207.380 1925.000 1207.640 ;
        RECT 1924.740 27.580 1925.000 27.840 ;
        RECT 2274.340 27.580 2274.600 27.840 ;
      LAYER met2 ;
        RECT 1918.310 1219.680 1918.870 1228.680 ;
        RECT 1918.360 1207.670 1918.500 1219.680 ;
        RECT 1918.300 1207.350 1918.560 1207.670 ;
        RECT 1924.740 1207.350 1925.000 1207.670 ;
        RECT 1924.800 27.870 1924.940 1207.350 ;
        RECT 1924.740 27.550 1925.000 27.870 ;
        RECT 2274.340 27.550 2274.600 27.870 ;
        RECT 2274.400 2.400 2274.540 27.550 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1927.010 1207.580 1927.330 1207.640 ;
        RECT 1931.610 1207.580 1931.930 1207.640 ;
        RECT 1927.010 1207.440 1931.930 1207.580 ;
        RECT 1927.010 1207.380 1927.330 1207.440 ;
        RECT 1931.610 1207.380 1931.930 1207.440 ;
        RECT 1931.610 28.120 1931.930 28.180 ;
        RECT 2292.250 28.120 2292.570 28.180 ;
        RECT 1931.610 27.980 2292.570 28.120 ;
        RECT 1931.610 27.920 1931.930 27.980 ;
        RECT 2292.250 27.920 2292.570 27.980 ;
      LAYER via ;
        RECT 1927.040 1207.380 1927.300 1207.640 ;
        RECT 1931.640 1207.380 1931.900 1207.640 ;
        RECT 1931.640 27.920 1931.900 28.180 ;
        RECT 2292.280 27.920 2292.540 28.180 ;
      LAYER met2 ;
        RECT 1927.050 1219.680 1927.610 1228.680 ;
        RECT 1927.100 1207.670 1927.240 1219.680 ;
        RECT 1927.040 1207.350 1927.300 1207.670 ;
        RECT 1931.640 1207.350 1931.900 1207.670 ;
        RECT 1931.700 28.210 1931.840 1207.350 ;
        RECT 1931.640 27.890 1931.900 28.210 ;
        RECT 2292.280 27.890 2292.540 28.210 ;
        RECT 2292.340 2.400 2292.480 27.890 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 28.460 1938.830 28.520 ;
        RECT 2310.190 28.460 2310.510 28.520 ;
        RECT 1938.510 28.320 2310.510 28.460 ;
        RECT 1938.510 28.260 1938.830 28.320 ;
        RECT 2310.190 28.260 2310.510 28.320 ;
      LAYER via ;
        RECT 1938.540 28.260 1938.800 28.520 ;
        RECT 2310.220 28.260 2310.480 28.520 ;
      LAYER met2 ;
        RECT 1936.250 1220.330 1936.810 1228.680 ;
        RECT 1936.250 1220.190 1938.740 1220.330 ;
        RECT 1936.250 1219.680 1936.810 1220.190 ;
        RECT 1938.600 28.550 1938.740 1220.190 ;
        RECT 1938.540 28.230 1938.800 28.550 ;
        RECT 2310.220 28.230 2310.480 28.550 ;
        RECT 2310.280 2.400 2310.420 28.230 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1945.410 28.800 1945.730 28.860 ;
        RECT 2328.130 28.800 2328.450 28.860 ;
        RECT 1945.410 28.660 2328.450 28.800 ;
        RECT 1945.410 28.600 1945.730 28.660 ;
        RECT 2328.130 28.600 2328.450 28.660 ;
      LAYER via ;
        RECT 1945.440 28.600 1945.700 28.860 ;
        RECT 2328.160 28.600 2328.420 28.860 ;
      LAYER met2 ;
        RECT 1945.450 1219.680 1946.010 1228.680 ;
        RECT 1945.500 28.890 1945.640 1219.680 ;
        RECT 1945.440 28.570 1945.700 28.890 ;
        RECT 2328.160 28.570 2328.420 28.890 ;
        RECT 2328.220 2.400 2328.360 28.570 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1954.610 1207.580 1954.930 1207.640 ;
        RECT 1959.210 1207.580 1959.530 1207.640 ;
        RECT 1954.610 1207.440 1959.530 1207.580 ;
        RECT 1954.610 1207.380 1954.930 1207.440 ;
        RECT 1959.210 1207.380 1959.530 1207.440 ;
        RECT 1959.210 29.140 1959.530 29.200 ;
        RECT 2345.610 29.140 2345.930 29.200 ;
        RECT 1959.210 29.000 2345.930 29.140 ;
        RECT 1959.210 28.940 1959.530 29.000 ;
        RECT 2345.610 28.940 2345.930 29.000 ;
      LAYER via ;
        RECT 1954.640 1207.380 1954.900 1207.640 ;
        RECT 1959.240 1207.380 1959.500 1207.640 ;
        RECT 1959.240 28.940 1959.500 29.200 ;
        RECT 2345.640 28.940 2345.900 29.200 ;
      LAYER met2 ;
        RECT 1954.650 1219.680 1955.210 1228.680 ;
        RECT 1954.700 1207.670 1954.840 1219.680 ;
        RECT 1954.640 1207.350 1954.900 1207.670 ;
        RECT 1959.240 1207.350 1959.500 1207.670 ;
        RECT 1959.300 29.230 1959.440 1207.350 ;
        RECT 1959.240 28.910 1959.500 29.230 ;
        RECT 2345.640 28.910 2345.900 29.230 ;
        RECT 2345.700 2.400 2345.840 28.910 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 29.480 1966.430 29.540 ;
        RECT 2363.550 29.480 2363.870 29.540 ;
        RECT 1966.110 29.340 2363.870 29.480 ;
        RECT 1966.110 29.280 1966.430 29.340 ;
        RECT 2363.550 29.280 2363.870 29.340 ;
      LAYER via ;
        RECT 1966.140 29.280 1966.400 29.540 ;
        RECT 2363.580 29.280 2363.840 29.540 ;
      LAYER met2 ;
        RECT 1963.850 1220.330 1964.410 1228.680 ;
        RECT 1963.850 1220.190 1966.340 1220.330 ;
        RECT 1963.850 1219.680 1964.410 1220.190 ;
        RECT 1966.200 29.570 1966.340 1220.190 ;
        RECT 1966.140 29.250 1966.400 29.570 ;
        RECT 2363.580 29.250 2363.840 29.570 ;
        RECT 2363.640 2.400 2363.780 29.250 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.010 29.820 1973.330 29.880 ;
        RECT 2381.490 29.820 2381.810 29.880 ;
        RECT 1973.010 29.680 2381.810 29.820 ;
        RECT 1973.010 29.620 1973.330 29.680 ;
        RECT 2381.490 29.620 2381.810 29.680 ;
      LAYER via ;
        RECT 1973.040 29.620 1973.300 29.880 ;
        RECT 2381.520 29.620 2381.780 29.880 ;
      LAYER met2 ;
        RECT 1973.050 1219.680 1973.610 1228.680 ;
        RECT 1973.100 29.910 1973.240 1219.680 ;
        RECT 1973.040 29.590 1973.300 29.910 ;
        RECT 2381.520 29.590 2381.780 29.910 ;
        RECT 2381.580 2.400 2381.720 29.590 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1982.210 1207.580 1982.530 1207.640 ;
        RECT 1986.810 1207.580 1987.130 1207.640 ;
        RECT 1982.210 1207.440 1987.130 1207.580 ;
        RECT 1982.210 1207.380 1982.530 1207.440 ;
        RECT 1986.810 1207.380 1987.130 1207.440 ;
        RECT 1986.810 30.160 1987.130 30.220 ;
        RECT 2399.430 30.160 2399.750 30.220 ;
        RECT 1986.810 30.020 2399.750 30.160 ;
        RECT 1986.810 29.960 1987.130 30.020 ;
        RECT 2399.430 29.960 2399.750 30.020 ;
      LAYER via ;
        RECT 1982.240 1207.380 1982.500 1207.640 ;
        RECT 1986.840 1207.380 1987.100 1207.640 ;
        RECT 1986.840 29.960 1987.100 30.220 ;
        RECT 2399.460 29.960 2399.720 30.220 ;
      LAYER met2 ;
        RECT 1982.250 1219.680 1982.810 1228.680 ;
        RECT 1982.300 1207.670 1982.440 1219.680 ;
        RECT 1982.240 1207.350 1982.500 1207.670 ;
        RECT 1986.840 1207.350 1987.100 1207.670 ;
        RECT 1986.900 30.250 1987.040 1207.350 ;
        RECT 1986.840 29.930 1987.100 30.250 ;
        RECT 2399.460 29.930 2399.720 30.250 ;
        RECT 2399.520 2.400 2399.660 29.930 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.370 1196.700 1152.690 1196.760 ;
        RECT 1155.590 1196.700 1155.910 1196.760 ;
        RECT 1152.370 1196.560 1155.910 1196.700 ;
        RECT 1152.370 1196.500 1152.690 1196.560 ;
        RECT 1155.590 1196.500 1155.910 1196.560 ;
        RECT 794.950 25.060 795.270 25.120 ;
        RECT 1152.370 25.060 1152.690 25.120 ;
        RECT 794.950 24.920 1152.690 25.060 ;
        RECT 794.950 24.860 795.270 24.920 ;
        RECT 1152.370 24.860 1152.690 24.920 ;
      LAYER via ;
        RECT 1152.400 1196.500 1152.660 1196.760 ;
        RECT 1155.620 1196.500 1155.880 1196.760 ;
        RECT 794.980 24.860 795.240 25.120 ;
        RECT 1152.400 24.860 1152.660 25.120 ;
      LAYER met2 ;
        RECT 1157.470 1220.330 1158.030 1228.680 ;
        RECT 1155.680 1220.190 1158.030 1220.330 ;
        RECT 1155.680 1196.790 1155.820 1220.190 ;
        RECT 1157.470 1219.680 1158.030 1220.190 ;
        RECT 1152.400 1196.470 1152.660 1196.790 ;
        RECT 1155.620 1196.470 1155.880 1196.790 ;
        RECT 1152.460 25.150 1152.600 1196.470 ;
        RECT 794.980 24.830 795.240 25.150 ;
        RECT 1152.400 24.830 1152.660 25.150 ;
        RECT 795.040 12.650 795.180 24.830 ;
        RECT 793.660 12.510 795.180 12.650 ;
        RECT 793.660 2.400 793.800 12.510 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 37.300 639.330 37.360 ;
        RECT 1076.930 37.300 1077.250 37.360 ;
        RECT 639.010 37.160 1077.250 37.300 ;
        RECT 639.010 37.100 639.330 37.160 ;
        RECT 1076.930 37.100 1077.250 37.160 ;
      LAYER via ;
        RECT 639.040 37.100 639.300 37.360 ;
        RECT 1076.960 37.100 1077.220 37.360 ;
      LAYER met2 ;
        RECT 1077.890 1220.330 1078.450 1228.680 ;
        RECT 1077.020 1220.190 1078.450 1220.330 ;
        RECT 1077.020 37.390 1077.160 1220.190 ;
        RECT 1077.890 1219.680 1078.450 1220.190 ;
        RECT 639.040 37.070 639.300 37.390 ;
        RECT 1076.960 37.070 1077.220 37.390 ;
        RECT 639.100 2.400 639.240 37.070 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1994.630 1207.580 1994.950 1207.640 ;
        RECT 2000.610 1207.580 2000.930 1207.640 ;
        RECT 1994.630 1207.440 2000.930 1207.580 ;
        RECT 1994.630 1207.380 1994.950 1207.440 ;
        RECT 2000.610 1207.380 2000.930 1207.440 ;
        RECT 2000.610 30.500 2000.930 30.560 ;
        RECT 2422.890 30.500 2423.210 30.560 ;
        RECT 2000.610 30.360 2423.210 30.500 ;
        RECT 2000.610 30.300 2000.930 30.360 ;
        RECT 2422.890 30.300 2423.210 30.360 ;
      LAYER via ;
        RECT 1994.660 1207.380 1994.920 1207.640 ;
        RECT 2000.640 1207.380 2000.900 1207.640 ;
        RECT 2000.640 30.300 2000.900 30.560 ;
        RECT 2422.920 30.300 2423.180 30.560 ;
      LAYER met2 ;
        RECT 1994.670 1219.680 1995.230 1228.680 ;
        RECT 1994.720 1207.670 1994.860 1219.680 ;
        RECT 1994.660 1207.350 1994.920 1207.670 ;
        RECT 2000.640 1207.350 2000.900 1207.670 ;
        RECT 2000.700 30.590 2000.840 1207.350 ;
        RECT 2000.640 30.270 2000.900 30.590 ;
        RECT 2422.920 30.270 2423.180 30.590 ;
        RECT 2422.980 2.400 2423.120 30.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2003.830 1207.580 2004.150 1207.640 ;
        RECT 2007.510 1207.580 2007.830 1207.640 ;
        RECT 2003.830 1207.440 2007.830 1207.580 ;
        RECT 2003.830 1207.380 2004.150 1207.440 ;
        RECT 2007.510 1207.380 2007.830 1207.440 ;
        RECT 2007.510 33.900 2007.830 33.960 ;
        RECT 2440.830 33.900 2441.150 33.960 ;
        RECT 2007.510 33.760 2441.150 33.900 ;
        RECT 2007.510 33.700 2007.830 33.760 ;
        RECT 2440.830 33.700 2441.150 33.760 ;
      LAYER via ;
        RECT 2003.860 1207.380 2004.120 1207.640 ;
        RECT 2007.540 1207.380 2007.800 1207.640 ;
        RECT 2007.540 33.700 2007.800 33.960 ;
        RECT 2440.860 33.700 2441.120 33.960 ;
      LAYER met2 ;
        RECT 2003.870 1219.680 2004.430 1228.680 ;
        RECT 2003.920 1207.670 2004.060 1219.680 ;
        RECT 2003.860 1207.350 2004.120 1207.670 ;
        RECT 2007.540 1207.350 2007.800 1207.670 ;
        RECT 2007.600 33.990 2007.740 1207.350 ;
        RECT 2007.540 33.670 2007.800 33.990 ;
        RECT 2440.860 33.670 2441.120 33.990 ;
        RECT 2440.920 2.400 2441.060 33.670 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2014.410 33.560 2014.730 33.620 ;
        RECT 2458.770 33.560 2459.090 33.620 ;
        RECT 2014.410 33.420 2459.090 33.560 ;
        RECT 2014.410 33.360 2014.730 33.420 ;
        RECT 2458.770 33.360 2459.090 33.420 ;
      LAYER via ;
        RECT 2014.440 33.360 2014.700 33.620 ;
        RECT 2458.800 33.360 2459.060 33.620 ;
      LAYER met2 ;
        RECT 2012.610 1220.330 2013.170 1228.680 ;
        RECT 2012.610 1220.190 2014.640 1220.330 ;
        RECT 2012.610 1219.680 2013.170 1220.190 ;
        RECT 2014.500 33.650 2014.640 1220.190 ;
        RECT 2014.440 33.330 2014.700 33.650 ;
        RECT 2458.800 33.330 2459.060 33.650 ;
        RECT 2458.860 2.400 2459.000 33.330 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2021.770 1207.580 2022.090 1207.640 ;
        RECT 2028.210 1207.580 2028.530 1207.640 ;
        RECT 2021.770 1207.440 2028.530 1207.580 ;
        RECT 2021.770 1207.380 2022.090 1207.440 ;
        RECT 2028.210 1207.380 2028.530 1207.440 ;
        RECT 2028.210 33.220 2028.530 33.280 ;
        RECT 2476.710 33.220 2477.030 33.280 ;
        RECT 2028.210 33.080 2477.030 33.220 ;
        RECT 2028.210 33.020 2028.530 33.080 ;
        RECT 2476.710 33.020 2477.030 33.080 ;
      LAYER via ;
        RECT 2021.800 1207.380 2022.060 1207.640 ;
        RECT 2028.240 1207.380 2028.500 1207.640 ;
        RECT 2028.240 33.020 2028.500 33.280 ;
        RECT 2476.740 33.020 2477.000 33.280 ;
      LAYER met2 ;
        RECT 2021.810 1219.680 2022.370 1228.680 ;
        RECT 2021.860 1207.670 2022.000 1219.680 ;
        RECT 2021.800 1207.350 2022.060 1207.670 ;
        RECT 2028.240 1207.350 2028.500 1207.670 ;
        RECT 2028.300 33.310 2028.440 1207.350 ;
        RECT 2028.240 32.990 2028.500 33.310 ;
        RECT 2476.740 32.990 2477.000 33.310 ;
        RECT 2476.800 2.400 2476.940 32.990 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2030.970 1207.580 2031.290 1207.640 ;
        RECT 2035.110 1207.580 2035.430 1207.640 ;
        RECT 2030.970 1207.440 2035.430 1207.580 ;
        RECT 2030.970 1207.380 2031.290 1207.440 ;
        RECT 2035.110 1207.380 2035.430 1207.440 ;
        RECT 2035.110 32.880 2035.430 32.940 ;
        RECT 2494.650 32.880 2494.970 32.940 ;
        RECT 2035.110 32.740 2494.970 32.880 ;
        RECT 2035.110 32.680 2035.430 32.740 ;
        RECT 2494.650 32.680 2494.970 32.740 ;
      LAYER via ;
        RECT 2031.000 1207.380 2031.260 1207.640 ;
        RECT 2035.140 1207.380 2035.400 1207.640 ;
        RECT 2035.140 32.680 2035.400 32.940 ;
        RECT 2494.680 32.680 2494.940 32.940 ;
      LAYER met2 ;
        RECT 2031.010 1219.680 2031.570 1228.680 ;
        RECT 2031.060 1207.670 2031.200 1219.680 ;
        RECT 2031.000 1207.350 2031.260 1207.670 ;
        RECT 2035.140 1207.350 2035.400 1207.670 ;
        RECT 2035.200 32.970 2035.340 1207.350 ;
        RECT 2035.140 32.650 2035.400 32.970 ;
        RECT 2494.680 32.650 2494.940 32.970 ;
        RECT 2494.740 2.400 2494.880 32.650 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2042.010 32.540 2042.330 32.600 ;
        RECT 2512.130 32.540 2512.450 32.600 ;
        RECT 2042.010 32.400 2512.450 32.540 ;
        RECT 2042.010 32.340 2042.330 32.400 ;
        RECT 2512.130 32.340 2512.450 32.400 ;
      LAYER via ;
        RECT 2042.040 32.340 2042.300 32.600 ;
        RECT 2512.160 32.340 2512.420 32.600 ;
      LAYER met2 ;
        RECT 2040.210 1220.330 2040.770 1228.680 ;
        RECT 2040.210 1220.190 2042.240 1220.330 ;
        RECT 2040.210 1219.680 2040.770 1220.190 ;
        RECT 2042.100 32.630 2042.240 1220.190 ;
        RECT 2042.040 32.310 2042.300 32.630 ;
        RECT 2512.160 32.310 2512.420 32.630 ;
        RECT 2512.220 2.400 2512.360 32.310 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2049.370 1207.580 2049.690 1207.640 ;
        RECT 2055.810 1207.580 2056.130 1207.640 ;
        RECT 2049.370 1207.440 2056.130 1207.580 ;
        RECT 2049.370 1207.380 2049.690 1207.440 ;
        RECT 2055.810 1207.380 2056.130 1207.440 ;
        RECT 2055.810 32.200 2056.130 32.260 ;
        RECT 2530.070 32.200 2530.390 32.260 ;
        RECT 2055.810 32.060 2530.390 32.200 ;
        RECT 2055.810 32.000 2056.130 32.060 ;
        RECT 2530.070 32.000 2530.390 32.060 ;
      LAYER via ;
        RECT 2049.400 1207.380 2049.660 1207.640 ;
        RECT 2055.840 1207.380 2056.100 1207.640 ;
        RECT 2055.840 32.000 2056.100 32.260 ;
        RECT 2530.100 32.000 2530.360 32.260 ;
      LAYER met2 ;
        RECT 2049.410 1219.680 2049.970 1228.680 ;
        RECT 2049.460 1207.670 2049.600 1219.680 ;
        RECT 2049.400 1207.350 2049.660 1207.670 ;
        RECT 2055.840 1207.350 2056.100 1207.670 ;
        RECT 2055.900 32.290 2056.040 1207.350 ;
        RECT 2055.840 31.970 2056.100 32.290 ;
        RECT 2530.100 31.970 2530.360 32.290 ;
        RECT 2530.160 2.400 2530.300 31.970 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2058.570 1211.320 2058.890 1211.380 ;
        RECT 2062.710 1211.320 2063.030 1211.380 ;
        RECT 2058.570 1211.180 2063.030 1211.320 ;
        RECT 2058.570 1211.120 2058.890 1211.180 ;
        RECT 2062.710 1211.120 2063.030 1211.180 ;
        RECT 2062.710 31.860 2063.030 31.920 ;
        RECT 2548.010 31.860 2548.330 31.920 ;
        RECT 2062.710 31.720 2548.330 31.860 ;
        RECT 2062.710 31.660 2063.030 31.720 ;
        RECT 2548.010 31.660 2548.330 31.720 ;
      LAYER via ;
        RECT 2058.600 1211.120 2058.860 1211.380 ;
        RECT 2062.740 1211.120 2063.000 1211.380 ;
        RECT 2062.740 31.660 2063.000 31.920 ;
        RECT 2548.040 31.660 2548.300 31.920 ;
      LAYER met2 ;
        RECT 2058.610 1219.680 2059.170 1228.680 ;
        RECT 2058.660 1211.410 2058.800 1219.680 ;
        RECT 2058.600 1211.090 2058.860 1211.410 ;
        RECT 2062.740 1211.090 2063.000 1211.410 ;
        RECT 2062.800 31.950 2062.940 1211.090 ;
        RECT 2062.740 31.630 2063.000 31.950 ;
        RECT 2548.040 31.630 2548.300 31.950 ;
        RECT 2548.100 2.400 2548.240 31.630 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2069.150 31.520 2069.470 31.580 ;
        RECT 2565.950 31.520 2566.270 31.580 ;
        RECT 2069.150 31.380 2566.270 31.520 ;
        RECT 2069.150 31.320 2069.470 31.380 ;
        RECT 2565.950 31.320 2566.270 31.380 ;
      LAYER via ;
        RECT 2069.180 31.320 2069.440 31.580 ;
        RECT 2565.980 31.320 2566.240 31.580 ;
      LAYER met2 ;
        RECT 2067.810 1220.330 2068.370 1228.680 ;
        RECT 2067.810 1220.190 2069.380 1220.330 ;
        RECT 2067.810 1219.680 2068.370 1220.190 ;
        RECT 2069.240 31.610 2069.380 1220.190 ;
        RECT 2069.180 31.290 2069.440 31.610 ;
        RECT 2565.980 31.290 2566.240 31.610 ;
        RECT 2566.040 2.400 2566.180 31.290 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2076.970 1210.640 2077.290 1210.700 ;
        RECT 2082.490 1210.640 2082.810 1210.700 ;
        RECT 2076.970 1210.500 2082.810 1210.640 ;
        RECT 2076.970 1210.440 2077.290 1210.500 ;
        RECT 2082.490 1210.440 2082.810 1210.500 ;
        RECT 2082.490 31.180 2082.810 31.240 ;
        RECT 2583.890 31.180 2584.210 31.240 ;
        RECT 2082.490 31.040 2584.210 31.180 ;
        RECT 2082.490 30.980 2082.810 31.040 ;
        RECT 2583.890 30.980 2584.210 31.040 ;
      LAYER via ;
        RECT 2077.000 1210.440 2077.260 1210.700 ;
        RECT 2082.520 1210.440 2082.780 1210.700 ;
        RECT 2082.520 30.980 2082.780 31.240 ;
        RECT 2583.920 30.980 2584.180 31.240 ;
      LAYER met2 ;
        RECT 2077.010 1219.680 2077.570 1228.680 ;
        RECT 2077.060 1210.730 2077.200 1219.680 ;
        RECT 2077.000 1210.410 2077.260 1210.730 ;
        RECT 2082.520 1210.410 2082.780 1210.730 ;
        RECT 2082.580 31.270 2082.720 1210.410 ;
        RECT 2082.520 30.950 2082.780 31.270 ;
        RECT 2583.920 30.950 2584.180 31.270 ;
        RECT 2583.980 2.400 2584.120 30.950 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1166.170 1183.440 1166.490 1183.500 ;
        RECT 1167.550 1183.440 1167.870 1183.500 ;
        RECT 1166.170 1183.300 1167.870 1183.440 ;
        RECT 1166.170 1183.240 1166.490 1183.300 ;
        RECT 1167.550 1183.240 1167.870 1183.300 ;
        RECT 817.490 25.400 817.810 25.460 ;
        RECT 1166.170 25.400 1166.490 25.460 ;
        RECT 817.490 25.260 1166.490 25.400 ;
        RECT 817.490 25.200 817.810 25.260 ;
        RECT 1166.170 25.200 1166.490 25.260 ;
      LAYER via ;
        RECT 1166.200 1183.240 1166.460 1183.500 ;
        RECT 1167.580 1183.240 1167.840 1183.500 ;
        RECT 817.520 25.200 817.780 25.460 ;
        RECT 1166.200 25.200 1166.460 25.460 ;
      LAYER met2 ;
        RECT 1169.430 1220.330 1169.990 1228.680 ;
        RECT 1167.640 1220.190 1169.990 1220.330 ;
        RECT 1167.640 1183.530 1167.780 1220.190 ;
        RECT 1169.430 1219.680 1169.990 1220.190 ;
        RECT 1166.200 1183.210 1166.460 1183.530 ;
        RECT 1167.580 1183.210 1167.840 1183.530 ;
        RECT 1166.260 25.490 1166.400 1183.210 ;
        RECT 817.520 25.170 817.780 25.490 ;
        RECT 1166.200 25.170 1166.460 25.490 ;
        RECT 817.580 2.400 817.720 25.170 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2086.170 1210.640 2086.490 1210.700 ;
        RECT 2090.310 1210.640 2090.630 1210.700 ;
        RECT 2086.170 1210.500 2090.630 1210.640 ;
        RECT 2086.170 1210.440 2086.490 1210.500 ;
        RECT 2090.310 1210.440 2090.630 1210.500 ;
        RECT 2090.310 30.840 2090.630 30.900 ;
        RECT 2601.370 30.840 2601.690 30.900 ;
        RECT 2090.310 30.700 2601.690 30.840 ;
        RECT 2090.310 30.640 2090.630 30.700 ;
        RECT 2601.370 30.640 2601.690 30.700 ;
      LAYER via ;
        RECT 2086.200 1210.440 2086.460 1210.700 ;
        RECT 2090.340 1210.440 2090.600 1210.700 ;
        RECT 2090.340 30.640 2090.600 30.900 ;
        RECT 2601.400 30.640 2601.660 30.900 ;
      LAYER met2 ;
        RECT 2086.210 1219.680 2086.770 1228.680 ;
        RECT 2086.260 1210.730 2086.400 1219.680 ;
        RECT 2086.200 1210.410 2086.460 1210.730 ;
        RECT 2090.340 1210.410 2090.600 1210.730 ;
        RECT 2090.400 30.930 2090.540 1210.410 ;
        RECT 2090.340 30.610 2090.600 30.930 ;
        RECT 2601.400 30.610 2601.660 30.930 ;
        RECT 2601.460 2.400 2601.600 30.610 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2096.750 37.640 2097.070 37.700 ;
        RECT 2619.310 37.640 2619.630 37.700 ;
        RECT 2096.750 37.500 2619.630 37.640 ;
        RECT 2096.750 37.440 2097.070 37.500 ;
        RECT 2619.310 37.440 2619.630 37.500 ;
      LAYER via ;
        RECT 2096.780 37.440 2097.040 37.700 ;
        RECT 2619.340 37.440 2619.600 37.700 ;
      LAYER met2 ;
        RECT 2095.410 1220.330 2095.970 1228.680 ;
        RECT 2095.410 1220.190 2096.980 1220.330 ;
        RECT 2095.410 1219.680 2095.970 1220.190 ;
        RECT 2096.840 37.730 2096.980 1220.190 ;
        RECT 2096.780 37.410 2097.040 37.730 ;
        RECT 2619.340 37.410 2619.600 37.730 ;
        RECT 2619.400 2.400 2619.540 37.410 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2104.570 1207.580 2104.890 1207.640 ;
        RECT 2110.550 1207.580 2110.870 1207.640 ;
        RECT 2104.570 1207.440 2110.870 1207.580 ;
        RECT 2104.570 1207.380 2104.890 1207.440 ;
        RECT 2110.550 1207.380 2110.870 1207.440 ;
        RECT 2110.550 41.380 2110.870 41.440 ;
        RECT 2637.250 41.380 2637.570 41.440 ;
        RECT 2110.550 41.240 2637.570 41.380 ;
        RECT 2110.550 41.180 2110.870 41.240 ;
        RECT 2637.250 41.180 2637.570 41.240 ;
      LAYER via ;
        RECT 2104.600 1207.380 2104.860 1207.640 ;
        RECT 2110.580 1207.380 2110.840 1207.640 ;
        RECT 2110.580 41.180 2110.840 41.440 ;
        RECT 2637.280 41.180 2637.540 41.440 ;
      LAYER met2 ;
        RECT 2104.610 1219.680 2105.170 1228.680 ;
        RECT 2104.660 1207.670 2104.800 1219.680 ;
        RECT 2104.600 1207.350 2104.860 1207.670 ;
        RECT 2110.580 1207.350 2110.840 1207.670 ;
        RECT 2110.640 41.470 2110.780 1207.350 ;
        RECT 2110.580 41.150 2110.840 41.470 ;
        RECT 2637.280 41.150 2637.540 41.470 ;
        RECT 2637.340 2.400 2637.480 41.150 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2116.145 1196.205 2116.315 1207.255 ;
        RECT 2116.145 1110.865 2116.315 1124.975 ;
        RECT 2116.145 1014.305 2116.315 1028.415 ;
        RECT 2116.145 966.365 2116.315 1013.795 ;
        RECT 2115.685 917.745 2115.855 931.855 ;
        RECT 2116.145 814.385 2116.315 862.495 ;
        RECT 2116.145 717.825 2116.315 765.935 ;
        RECT 2116.145 565.845 2116.315 613.955 ;
        RECT 2115.225 524.365 2115.395 548.675 ;
      LAYER mcon ;
        RECT 2116.145 1207.085 2116.315 1207.255 ;
        RECT 2116.145 1124.805 2116.315 1124.975 ;
        RECT 2116.145 1028.245 2116.315 1028.415 ;
        RECT 2116.145 1013.625 2116.315 1013.795 ;
        RECT 2115.685 931.685 2115.855 931.855 ;
        RECT 2116.145 862.325 2116.315 862.495 ;
        RECT 2116.145 765.765 2116.315 765.935 ;
        RECT 2116.145 613.785 2116.315 613.955 ;
        RECT 2115.225 548.505 2115.395 548.675 ;
      LAYER met1 ;
        RECT 2116.070 1207.240 2116.390 1207.300 ;
        RECT 2115.875 1207.100 2116.390 1207.240 ;
        RECT 2116.070 1207.040 2116.390 1207.100 ;
        RECT 2116.085 1196.360 2116.375 1196.405 ;
        RECT 2116.530 1196.360 2116.850 1196.420 ;
        RECT 2116.085 1196.220 2116.850 1196.360 ;
        RECT 2116.085 1196.175 2116.375 1196.220 ;
        RECT 2116.530 1196.160 2116.850 1196.220 ;
        RECT 2116.070 1124.960 2116.390 1125.020 ;
        RECT 2115.875 1124.820 2116.390 1124.960 ;
        RECT 2116.070 1124.760 2116.390 1124.820 ;
        RECT 2116.070 1111.020 2116.390 1111.080 ;
        RECT 2115.875 1110.880 2116.390 1111.020 ;
        RECT 2116.070 1110.820 2116.390 1110.880 ;
        RECT 2116.070 1076.820 2116.390 1077.080 ;
        RECT 2116.160 1076.400 2116.300 1076.820 ;
        RECT 2116.070 1076.140 2116.390 1076.400 ;
        RECT 2116.070 1028.400 2116.390 1028.460 ;
        RECT 2115.875 1028.260 2116.390 1028.400 ;
        RECT 2116.070 1028.200 2116.390 1028.260 ;
        RECT 2116.070 1014.460 2116.390 1014.520 ;
        RECT 2115.875 1014.320 2116.390 1014.460 ;
        RECT 2116.070 1014.260 2116.390 1014.320 ;
        RECT 2116.070 1013.780 2116.390 1013.840 ;
        RECT 2115.875 1013.640 2116.390 1013.780 ;
        RECT 2116.070 1013.580 2116.390 1013.640 ;
        RECT 2116.085 966.520 2116.375 966.565 ;
        RECT 2116.530 966.520 2116.850 966.580 ;
        RECT 2116.085 966.380 2116.850 966.520 ;
        RECT 2116.085 966.335 2116.375 966.380 ;
        RECT 2116.530 966.320 2116.850 966.380 ;
        RECT 2115.625 931.840 2115.915 931.885 ;
        RECT 2116.070 931.840 2116.390 931.900 ;
        RECT 2115.625 931.700 2116.390 931.840 ;
        RECT 2115.625 931.655 2115.915 931.700 ;
        RECT 2116.070 931.640 2116.390 931.700 ;
        RECT 2115.610 917.900 2115.930 917.960 ;
        RECT 2115.415 917.760 2115.930 917.900 ;
        RECT 2115.610 917.700 2115.930 917.760 ;
        RECT 2115.610 910.760 2115.930 910.820 ;
        RECT 2116.070 910.760 2116.390 910.820 ;
        RECT 2115.610 910.620 2116.390 910.760 ;
        RECT 2115.610 910.560 2115.930 910.620 ;
        RECT 2116.070 910.560 2116.390 910.620 ;
        RECT 2116.085 862.480 2116.375 862.525 ;
        RECT 2116.530 862.480 2116.850 862.540 ;
        RECT 2116.085 862.340 2116.850 862.480 ;
        RECT 2116.085 862.295 2116.375 862.340 ;
        RECT 2116.530 862.280 2116.850 862.340 ;
        RECT 2116.070 814.540 2116.390 814.600 ;
        RECT 2115.875 814.400 2116.390 814.540 ;
        RECT 2116.070 814.340 2116.390 814.400 ;
        RECT 2116.070 786.800 2116.390 787.060 ;
        RECT 2116.160 786.320 2116.300 786.800 ;
        RECT 2116.530 786.320 2116.850 786.380 ;
        RECT 2116.160 786.180 2116.850 786.320 ;
        RECT 2116.530 786.120 2116.850 786.180 ;
        RECT 2116.085 765.920 2116.375 765.965 ;
        RECT 2116.530 765.920 2116.850 765.980 ;
        RECT 2116.085 765.780 2116.850 765.920 ;
        RECT 2116.085 765.735 2116.375 765.780 ;
        RECT 2116.530 765.720 2116.850 765.780 ;
        RECT 2116.070 717.980 2116.390 718.040 ;
        RECT 2115.875 717.840 2116.390 717.980 ;
        RECT 2116.070 717.780 2116.390 717.840 ;
        RECT 2116.070 689.900 2116.390 690.160 ;
        RECT 2116.160 689.760 2116.300 689.900 ;
        RECT 2116.530 689.760 2116.850 689.820 ;
        RECT 2116.160 689.620 2116.850 689.760 ;
        RECT 2116.530 689.560 2116.850 689.620 ;
        RECT 2116.530 645.220 2116.850 645.280 ;
        RECT 2117.450 645.220 2117.770 645.280 ;
        RECT 2116.530 645.080 2117.770 645.220 ;
        RECT 2116.530 645.020 2116.850 645.080 ;
        RECT 2117.450 645.020 2117.770 645.080 ;
        RECT 2116.070 613.940 2116.390 614.000 ;
        RECT 2115.875 613.800 2116.390 613.940 ;
        RECT 2116.070 613.740 2116.390 613.800 ;
        RECT 2116.085 566.000 2116.375 566.045 ;
        RECT 2116.530 566.000 2116.850 566.060 ;
        RECT 2116.085 565.860 2116.850 566.000 ;
        RECT 2116.085 565.815 2116.375 565.860 ;
        RECT 2116.530 565.800 2116.850 565.860 ;
        RECT 2115.165 548.660 2115.455 548.705 ;
        RECT 2116.530 548.660 2116.850 548.720 ;
        RECT 2115.165 548.520 2116.850 548.660 ;
        RECT 2115.165 548.475 2115.455 548.520 ;
        RECT 2116.530 548.460 2116.850 548.520 ;
        RECT 2115.150 524.520 2115.470 524.580 ;
        RECT 2114.955 524.380 2115.470 524.520 ;
        RECT 2115.150 524.320 2115.470 524.380 ;
        RECT 2115.150 483.040 2115.470 483.100 ;
        RECT 2115.610 483.040 2115.930 483.100 ;
        RECT 2115.150 482.900 2115.930 483.040 ;
        RECT 2115.150 482.840 2115.470 482.900 ;
        RECT 2115.610 482.840 2115.930 482.900 ;
        RECT 2116.070 434.760 2116.390 434.820 ;
        RECT 2116.990 434.760 2117.310 434.820 ;
        RECT 2116.070 434.620 2117.310 434.760 ;
        RECT 2116.070 434.560 2116.390 434.620 ;
        RECT 2116.990 434.560 2117.310 434.620 ;
        RECT 2116.070 338.200 2116.390 338.260 ;
        RECT 2116.530 338.200 2116.850 338.260 ;
        RECT 2116.070 338.060 2116.850 338.200 ;
        RECT 2116.070 338.000 2116.390 338.060 ;
        RECT 2116.530 338.000 2116.850 338.060 ;
        RECT 2116.070 290.260 2116.390 290.320 ;
        RECT 2117.450 290.260 2117.770 290.320 ;
        RECT 2116.070 290.120 2117.770 290.260 ;
        RECT 2116.070 290.060 2116.390 290.120 ;
        RECT 2117.450 290.060 2117.770 290.120 ;
        RECT 2116.530 193.700 2116.850 193.760 ;
        RECT 2117.450 193.700 2117.770 193.760 ;
        RECT 2116.530 193.560 2117.770 193.700 ;
        RECT 2116.530 193.500 2116.850 193.560 ;
        RECT 2117.450 193.500 2117.770 193.560 ;
        RECT 2116.530 158.820 2116.850 159.080 ;
        RECT 2116.620 158.340 2116.760 158.820 ;
        RECT 2116.990 158.340 2117.310 158.400 ;
        RECT 2116.620 158.200 2117.310 158.340 ;
        RECT 2116.990 158.140 2117.310 158.200 ;
        RECT 2116.990 41.040 2117.310 41.100 ;
        RECT 2655.190 41.040 2655.510 41.100 ;
        RECT 2116.990 40.900 2655.510 41.040 ;
        RECT 2116.990 40.840 2117.310 40.900 ;
        RECT 2655.190 40.840 2655.510 40.900 ;
      LAYER via ;
        RECT 2116.100 1207.040 2116.360 1207.300 ;
        RECT 2116.560 1196.160 2116.820 1196.420 ;
        RECT 2116.100 1124.760 2116.360 1125.020 ;
        RECT 2116.100 1110.820 2116.360 1111.080 ;
        RECT 2116.100 1076.820 2116.360 1077.080 ;
        RECT 2116.100 1076.140 2116.360 1076.400 ;
        RECT 2116.100 1028.200 2116.360 1028.460 ;
        RECT 2116.100 1014.260 2116.360 1014.520 ;
        RECT 2116.100 1013.580 2116.360 1013.840 ;
        RECT 2116.560 966.320 2116.820 966.580 ;
        RECT 2116.100 931.640 2116.360 931.900 ;
        RECT 2115.640 917.700 2115.900 917.960 ;
        RECT 2115.640 910.560 2115.900 910.820 ;
        RECT 2116.100 910.560 2116.360 910.820 ;
        RECT 2116.560 862.280 2116.820 862.540 ;
        RECT 2116.100 814.340 2116.360 814.600 ;
        RECT 2116.100 786.800 2116.360 787.060 ;
        RECT 2116.560 786.120 2116.820 786.380 ;
        RECT 2116.560 765.720 2116.820 765.980 ;
        RECT 2116.100 717.780 2116.360 718.040 ;
        RECT 2116.100 689.900 2116.360 690.160 ;
        RECT 2116.560 689.560 2116.820 689.820 ;
        RECT 2116.560 645.020 2116.820 645.280 ;
        RECT 2117.480 645.020 2117.740 645.280 ;
        RECT 2116.100 613.740 2116.360 614.000 ;
        RECT 2116.560 565.800 2116.820 566.060 ;
        RECT 2116.560 548.460 2116.820 548.720 ;
        RECT 2115.180 524.320 2115.440 524.580 ;
        RECT 2115.180 482.840 2115.440 483.100 ;
        RECT 2115.640 482.840 2115.900 483.100 ;
        RECT 2116.100 434.560 2116.360 434.820 ;
        RECT 2117.020 434.560 2117.280 434.820 ;
        RECT 2116.100 338.000 2116.360 338.260 ;
        RECT 2116.560 338.000 2116.820 338.260 ;
        RECT 2116.100 290.060 2116.360 290.320 ;
        RECT 2117.480 290.060 2117.740 290.320 ;
        RECT 2116.560 193.500 2116.820 193.760 ;
        RECT 2117.480 193.500 2117.740 193.760 ;
        RECT 2116.560 158.820 2116.820 159.080 ;
        RECT 2117.020 158.140 2117.280 158.400 ;
        RECT 2117.020 40.840 2117.280 41.100 ;
        RECT 2655.220 40.840 2655.480 41.100 ;
      LAYER met2 ;
        RECT 2113.810 1221.010 2114.370 1228.680 ;
        RECT 2113.810 1220.870 2116.300 1221.010 ;
        RECT 2113.810 1219.680 2114.370 1220.870 ;
        RECT 2116.160 1207.330 2116.300 1220.870 ;
        RECT 2116.100 1207.010 2116.360 1207.330 ;
        RECT 2116.560 1196.130 2116.820 1196.450 ;
        RECT 2116.620 1159.130 2116.760 1196.130 ;
        RECT 2116.160 1158.990 2116.760 1159.130 ;
        RECT 2116.160 1125.050 2116.300 1158.990 ;
        RECT 2116.100 1124.730 2116.360 1125.050 ;
        RECT 2116.100 1110.790 2116.360 1111.110 ;
        RECT 2116.160 1077.110 2116.300 1110.790 ;
        RECT 2116.100 1076.790 2116.360 1077.110 ;
        RECT 2116.100 1076.110 2116.360 1076.430 ;
        RECT 2116.160 1028.490 2116.300 1076.110 ;
        RECT 2116.100 1028.170 2116.360 1028.490 ;
        RECT 2116.100 1014.230 2116.360 1014.550 ;
        RECT 2116.160 1013.870 2116.300 1014.230 ;
        RECT 2116.100 1013.550 2116.360 1013.870 ;
        RECT 2116.560 966.290 2116.820 966.610 ;
        RECT 2116.620 966.010 2116.760 966.290 ;
        RECT 2116.160 965.870 2116.760 966.010 ;
        RECT 2116.160 931.930 2116.300 965.870 ;
        RECT 2116.100 931.610 2116.360 931.930 ;
        RECT 2115.640 917.670 2115.900 917.990 ;
        RECT 2115.700 910.850 2115.840 917.670 ;
        RECT 2115.640 910.530 2115.900 910.850 ;
        RECT 2116.100 910.530 2116.360 910.850 ;
        RECT 2116.160 868.770 2116.300 910.530 ;
        RECT 2116.160 868.630 2116.760 868.770 ;
        RECT 2116.620 862.570 2116.760 868.630 ;
        RECT 2116.560 862.250 2116.820 862.570 ;
        RECT 2116.100 814.310 2116.360 814.630 ;
        RECT 2116.160 787.090 2116.300 814.310 ;
        RECT 2116.100 786.770 2116.360 787.090 ;
        RECT 2116.560 786.090 2116.820 786.410 ;
        RECT 2116.620 766.010 2116.760 786.090 ;
        RECT 2116.560 765.690 2116.820 766.010 ;
        RECT 2116.100 717.750 2116.360 718.070 ;
        RECT 2116.160 690.190 2116.300 717.750 ;
        RECT 2116.100 689.870 2116.360 690.190 ;
        RECT 2116.560 689.530 2116.820 689.850 ;
        RECT 2116.620 645.310 2116.760 689.530 ;
        RECT 2116.560 644.990 2116.820 645.310 ;
        RECT 2117.480 644.990 2117.740 645.310 ;
        RECT 2117.540 621.365 2117.680 644.990 ;
        RECT 2116.550 621.250 2116.830 621.365 ;
        RECT 2116.160 621.110 2116.830 621.250 ;
        RECT 2116.160 614.030 2116.300 621.110 ;
        RECT 2116.550 620.995 2116.830 621.110 ;
        RECT 2117.470 620.995 2117.750 621.365 ;
        RECT 2116.100 613.710 2116.360 614.030 ;
        RECT 2116.560 565.770 2116.820 566.090 ;
        RECT 2116.620 548.750 2116.760 565.770 ;
        RECT 2116.560 548.430 2116.820 548.750 ;
        RECT 2115.180 524.290 2115.440 524.610 ;
        RECT 2115.240 483.130 2115.380 524.290 ;
        RECT 2115.180 482.810 2115.440 483.130 ;
        RECT 2115.640 482.810 2115.900 483.130 ;
        RECT 2115.700 434.930 2115.840 482.810 ;
        RECT 2115.700 434.850 2116.300 434.930 ;
        RECT 2115.700 434.790 2116.360 434.850 ;
        RECT 2116.100 434.530 2116.360 434.790 ;
        RECT 2117.020 434.530 2117.280 434.850 ;
        RECT 2117.080 399.570 2117.220 434.530 ;
        RECT 2116.620 399.430 2117.220 399.570 ;
        RECT 2116.620 338.290 2116.760 399.430 ;
        RECT 2116.100 337.970 2116.360 338.290 ;
        RECT 2116.560 337.970 2116.820 338.290 ;
        RECT 2116.160 290.350 2116.300 337.970 ;
        RECT 2116.100 290.030 2116.360 290.350 ;
        RECT 2117.480 290.030 2117.740 290.350 ;
        RECT 2117.540 193.790 2117.680 290.030 ;
        RECT 2116.560 193.470 2116.820 193.790 ;
        RECT 2117.480 193.470 2117.740 193.790 ;
        RECT 2116.620 159.110 2116.760 193.470 ;
        RECT 2116.560 158.790 2116.820 159.110 ;
        RECT 2117.020 158.110 2117.280 158.430 ;
        RECT 2117.080 144.570 2117.220 158.110 ;
        RECT 2117.080 144.430 2117.680 144.570 ;
        RECT 2117.540 62.290 2117.680 144.430 ;
        RECT 2117.080 62.150 2117.680 62.290 ;
        RECT 2117.080 41.130 2117.220 62.150 ;
        RECT 2117.020 40.810 2117.280 41.130 ;
        RECT 2655.220 40.810 2655.480 41.130 ;
        RECT 2655.280 2.400 2655.420 40.810 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
      LAYER via2 ;
        RECT 2116.550 621.040 2116.830 621.320 ;
        RECT 2117.470 621.040 2117.750 621.320 ;
      LAYER met3 ;
        RECT 2116.525 621.330 2116.855 621.345 ;
        RECT 2117.445 621.330 2117.775 621.345 ;
        RECT 2116.525 621.030 2117.775 621.330 ;
        RECT 2116.525 621.015 2116.855 621.030 ;
        RECT 2117.445 621.015 2117.775 621.030 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.350 40.700 2124.670 40.760 ;
        RECT 2672.670 40.700 2672.990 40.760 ;
        RECT 2124.350 40.560 2672.990 40.700 ;
        RECT 2124.350 40.500 2124.670 40.560 ;
        RECT 2672.670 40.500 2672.990 40.560 ;
      LAYER via ;
        RECT 2124.380 40.500 2124.640 40.760 ;
        RECT 2672.700 40.500 2672.960 40.760 ;
      LAYER met2 ;
        RECT 2123.010 1220.330 2123.570 1228.680 ;
        RECT 2123.010 1220.190 2124.580 1220.330 ;
        RECT 2123.010 1219.680 2123.570 1220.190 ;
        RECT 2124.440 40.790 2124.580 1220.190 ;
        RECT 2124.380 40.470 2124.640 40.790 ;
        RECT 2672.700 40.470 2672.960 40.790 ;
        RECT 2672.760 2.400 2672.900 40.470 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2131.250 40.360 2131.570 40.420 ;
        RECT 2690.610 40.360 2690.930 40.420 ;
        RECT 2131.250 40.220 2690.930 40.360 ;
        RECT 2131.250 40.160 2131.570 40.220 ;
        RECT 2690.610 40.160 2690.930 40.220 ;
      LAYER via ;
        RECT 2131.280 40.160 2131.540 40.420 ;
        RECT 2690.640 40.160 2690.900 40.420 ;
      LAYER met2 ;
        RECT 2131.750 1220.330 2132.310 1228.680 ;
        RECT 2131.340 1220.190 2132.310 1220.330 ;
        RECT 2131.340 40.450 2131.480 1220.190 ;
        RECT 2131.750 1219.680 2132.310 1220.190 ;
        RECT 2131.280 40.130 2131.540 40.450 ;
        RECT 2690.640 40.130 2690.900 40.450 ;
        RECT 2690.700 2.400 2690.840 40.130 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2140.910 1207.580 2141.230 1207.640 ;
        RECT 2145.510 1207.580 2145.830 1207.640 ;
        RECT 2140.910 1207.440 2145.830 1207.580 ;
        RECT 2140.910 1207.380 2141.230 1207.440 ;
        RECT 2145.510 1207.380 2145.830 1207.440 ;
        RECT 2145.510 40.020 2145.830 40.080 ;
        RECT 2708.550 40.020 2708.870 40.080 ;
        RECT 2145.510 39.880 2708.870 40.020 ;
        RECT 2145.510 39.820 2145.830 39.880 ;
        RECT 2708.550 39.820 2708.870 39.880 ;
      LAYER via ;
        RECT 2140.940 1207.380 2141.200 1207.640 ;
        RECT 2145.540 1207.380 2145.800 1207.640 ;
        RECT 2145.540 39.820 2145.800 40.080 ;
        RECT 2708.580 39.820 2708.840 40.080 ;
      LAYER met2 ;
        RECT 2140.950 1219.680 2141.510 1228.680 ;
        RECT 2141.000 1207.670 2141.140 1219.680 ;
        RECT 2140.940 1207.350 2141.200 1207.670 ;
        RECT 2145.540 1207.350 2145.800 1207.670 ;
        RECT 2145.600 40.110 2145.740 1207.350 ;
        RECT 2145.540 39.790 2145.800 40.110 ;
        RECT 2708.580 39.790 2708.840 40.110 ;
        RECT 2708.640 2.400 2708.780 39.790 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2151.950 39.680 2152.270 39.740 ;
        RECT 2726.490 39.680 2726.810 39.740 ;
        RECT 2151.950 39.540 2726.810 39.680 ;
        RECT 2151.950 39.480 2152.270 39.540 ;
        RECT 2726.490 39.480 2726.810 39.540 ;
      LAYER via ;
        RECT 2151.980 39.480 2152.240 39.740 ;
        RECT 2726.520 39.480 2726.780 39.740 ;
      LAYER met2 ;
        RECT 2150.150 1220.330 2150.710 1228.680 ;
        RECT 2150.150 1220.190 2152.180 1220.330 ;
        RECT 2150.150 1219.680 2150.710 1220.190 ;
        RECT 2152.040 39.770 2152.180 1220.190 ;
        RECT 2151.980 39.450 2152.240 39.770 ;
        RECT 2726.520 39.450 2726.780 39.770 ;
        RECT 2726.580 2.400 2726.720 39.450 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2158.390 1207.580 2158.710 1207.640 ;
        RECT 2159.310 1207.580 2159.630 1207.640 ;
        RECT 2158.390 1207.440 2159.630 1207.580 ;
        RECT 2158.390 1207.380 2158.710 1207.440 ;
        RECT 2159.310 1207.380 2159.630 1207.440 ;
        RECT 2158.390 39.340 2158.710 39.400 ;
        RECT 2744.430 39.340 2744.750 39.400 ;
        RECT 2158.390 39.200 2744.750 39.340 ;
        RECT 2158.390 39.140 2158.710 39.200 ;
        RECT 2744.430 39.140 2744.750 39.200 ;
      LAYER via ;
        RECT 2158.420 1207.380 2158.680 1207.640 ;
        RECT 2159.340 1207.380 2159.600 1207.640 ;
        RECT 2158.420 39.140 2158.680 39.400 ;
        RECT 2744.460 39.140 2744.720 39.400 ;
      LAYER met2 ;
        RECT 2159.350 1219.680 2159.910 1228.680 ;
        RECT 2159.400 1207.670 2159.540 1219.680 ;
        RECT 2158.420 1207.350 2158.680 1207.670 ;
        RECT 2159.340 1207.350 2159.600 1207.670 ;
        RECT 2158.480 39.430 2158.620 1207.350 ;
        RECT 2158.420 39.110 2158.680 39.430 ;
        RECT 2744.460 39.110 2744.720 39.430 ;
        RECT 2744.520 2.400 2744.660 39.110 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2168.510 1207.580 2168.830 1207.640 ;
        RECT 2172.650 1207.580 2172.970 1207.640 ;
        RECT 2168.510 1207.440 2172.970 1207.580 ;
        RECT 2168.510 1207.380 2168.830 1207.440 ;
        RECT 2172.650 1207.380 2172.970 1207.440 ;
        RECT 2172.650 39.000 2172.970 39.060 ;
        RECT 2761.910 39.000 2762.230 39.060 ;
        RECT 2172.650 38.860 2762.230 39.000 ;
        RECT 2172.650 38.800 2172.970 38.860 ;
        RECT 2761.910 38.800 2762.230 38.860 ;
      LAYER via ;
        RECT 2168.540 1207.380 2168.800 1207.640 ;
        RECT 2172.680 1207.380 2172.940 1207.640 ;
        RECT 2172.680 38.800 2172.940 39.060 ;
        RECT 2761.940 38.800 2762.200 39.060 ;
      LAYER met2 ;
        RECT 2168.550 1219.680 2169.110 1228.680 ;
        RECT 2168.600 1207.670 2168.740 1219.680 ;
        RECT 2168.540 1207.350 2168.800 1207.670 ;
        RECT 2172.680 1207.350 2172.940 1207.670 ;
        RECT 2172.740 39.090 2172.880 1207.350 ;
        RECT 2172.680 38.770 2172.940 39.090 ;
        RECT 2761.940 38.770 2762.200 39.090 ;
        RECT 2762.000 2.400 2762.140 38.770 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1174.065 621.265 1174.235 669.375 ;
        RECT 1174.065 572.645 1174.235 620.755 ;
        RECT 1174.065 193.205 1174.235 241.315 ;
      LAYER mcon ;
        RECT 1174.065 669.205 1174.235 669.375 ;
        RECT 1174.065 620.585 1174.235 620.755 ;
        RECT 1174.065 241.145 1174.235 241.315 ;
      LAYER met1 ;
        RECT 1174.450 1159.300 1174.770 1159.360 ;
        RECT 1177.210 1159.300 1177.530 1159.360 ;
        RECT 1174.450 1159.160 1177.530 1159.300 ;
        RECT 1174.450 1159.100 1174.770 1159.160 ;
        RECT 1177.210 1159.100 1177.530 1159.160 ;
        RECT 1174.450 966.520 1174.770 966.580 ;
        RECT 1174.080 966.380 1174.770 966.520 ;
        RECT 1174.080 966.240 1174.220 966.380 ;
        RECT 1174.450 966.320 1174.770 966.380 ;
        RECT 1173.990 965.980 1174.310 966.240 ;
        RECT 1174.450 724.440 1174.770 724.500 ;
        RECT 1174.910 724.440 1175.230 724.500 ;
        RECT 1174.450 724.300 1175.230 724.440 ;
        RECT 1174.450 724.240 1174.770 724.300 ;
        RECT 1174.910 724.240 1175.230 724.300 ;
        RECT 1173.990 676.160 1174.310 676.220 ;
        RECT 1174.910 676.160 1175.230 676.220 ;
        RECT 1173.990 676.020 1175.230 676.160 ;
        RECT 1173.990 675.960 1174.310 676.020 ;
        RECT 1174.910 675.960 1175.230 676.020 ;
        RECT 1174.005 669.360 1174.295 669.405 ;
        RECT 1174.910 669.360 1175.230 669.420 ;
        RECT 1174.005 669.220 1175.230 669.360 ;
        RECT 1174.005 669.175 1174.295 669.220 ;
        RECT 1174.910 669.160 1175.230 669.220 ;
        RECT 1173.990 621.420 1174.310 621.480 ;
        RECT 1173.795 621.280 1174.310 621.420 ;
        RECT 1173.990 621.220 1174.310 621.280 ;
        RECT 1173.990 620.740 1174.310 620.800 ;
        RECT 1173.795 620.600 1174.310 620.740 ;
        RECT 1173.990 620.540 1174.310 620.600 ;
        RECT 1173.990 572.800 1174.310 572.860 ;
        RECT 1173.795 572.660 1174.310 572.800 ;
        RECT 1173.990 572.600 1174.310 572.660 ;
        RECT 1173.530 386.480 1173.850 386.540 ;
        RECT 1173.990 386.480 1174.310 386.540 ;
        RECT 1173.530 386.340 1174.310 386.480 ;
        RECT 1173.530 386.280 1173.850 386.340 ;
        RECT 1173.990 386.280 1174.310 386.340 ;
        RECT 1174.005 241.300 1174.295 241.345 ;
        RECT 1174.450 241.300 1174.770 241.360 ;
        RECT 1174.005 241.160 1174.770 241.300 ;
        RECT 1174.005 241.115 1174.295 241.160 ;
        RECT 1174.450 241.100 1174.770 241.160 ;
        RECT 1173.990 193.360 1174.310 193.420 ;
        RECT 1173.795 193.220 1174.310 193.360 ;
        RECT 1173.990 193.160 1174.310 193.220 ;
        RECT 1173.530 96.800 1173.850 96.860 ;
        RECT 1173.990 96.800 1174.310 96.860 ;
        RECT 1173.530 96.660 1174.310 96.800 ;
        RECT 1173.530 96.600 1173.850 96.660 ;
        RECT 1173.990 96.600 1174.310 96.660 ;
        RECT 835.890 25.740 836.210 25.800 ;
        RECT 1173.990 25.740 1174.310 25.800 ;
        RECT 835.890 25.600 1174.310 25.740 ;
        RECT 835.890 25.540 836.210 25.600 ;
        RECT 1173.990 25.540 1174.310 25.600 ;
      LAYER via ;
        RECT 1174.480 1159.100 1174.740 1159.360 ;
        RECT 1177.240 1159.100 1177.500 1159.360 ;
        RECT 1174.480 966.320 1174.740 966.580 ;
        RECT 1174.020 965.980 1174.280 966.240 ;
        RECT 1174.480 724.240 1174.740 724.500 ;
        RECT 1174.940 724.240 1175.200 724.500 ;
        RECT 1174.020 675.960 1174.280 676.220 ;
        RECT 1174.940 675.960 1175.200 676.220 ;
        RECT 1174.940 669.160 1175.200 669.420 ;
        RECT 1174.020 621.220 1174.280 621.480 ;
        RECT 1174.020 620.540 1174.280 620.800 ;
        RECT 1174.020 572.600 1174.280 572.860 ;
        RECT 1173.560 386.280 1173.820 386.540 ;
        RECT 1174.020 386.280 1174.280 386.540 ;
        RECT 1174.480 241.100 1174.740 241.360 ;
        RECT 1174.020 193.160 1174.280 193.420 ;
        RECT 1173.560 96.600 1173.820 96.860 ;
        RECT 1174.020 96.600 1174.280 96.860 ;
        RECT 835.920 25.540 836.180 25.800 ;
        RECT 1174.020 25.540 1174.280 25.800 ;
      LAYER met2 ;
        RECT 1178.630 1220.330 1179.190 1228.680 ;
        RECT 1177.300 1220.190 1179.190 1220.330 ;
        RECT 1177.300 1159.390 1177.440 1220.190 ;
        RECT 1178.630 1219.680 1179.190 1220.190 ;
        RECT 1174.480 1159.070 1174.740 1159.390 ;
        RECT 1177.240 1159.070 1177.500 1159.390 ;
        RECT 1174.540 1076.850 1174.680 1159.070 ;
        RECT 1174.080 1076.710 1174.680 1076.850 ;
        RECT 1174.080 1038.770 1174.220 1076.710 ;
        RECT 1174.080 1038.630 1174.680 1038.770 ;
        RECT 1174.540 966.610 1174.680 1038.630 ;
        RECT 1174.480 966.290 1174.740 966.610 ;
        RECT 1174.020 966.125 1174.280 966.270 ;
        RECT 1174.010 965.755 1174.290 966.125 ;
        RECT 1174.930 965.755 1175.210 966.125 ;
        RECT 1175.000 814.485 1175.140 965.755 ;
        RECT 1174.010 814.115 1174.290 814.485 ;
        RECT 1174.930 814.115 1175.210 814.485 ;
        RECT 1174.080 737.530 1174.220 814.115 ;
        RECT 1174.080 737.390 1174.680 737.530 ;
        RECT 1174.540 724.530 1174.680 737.390 ;
        RECT 1174.480 724.210 1174.740 724.530 ;
        RECT 1174.940 724.210 1175.200 724.530 ;
        RECT 1175.000 676.445 1175.140 724.210 ;
        RECT 1174.010 676.075 1174.290 676.445 ;
        RECT 1174.930 676.075 1175.210 676.445 ;
        RECT 1174.020 675.930 1174.280 676.075 ;
        RECT 1174.940 675.930 1175.200 676.075 ;
        RECT 1175.000 669.450 1175.140 675.930 ;
        RECT 1174.940 669.130 1175.200 669.450 ;
        RECT 1174.020 621.190 1174.280 621.510 ;
        RECT 1174.080 620.830 1174.220 621.190 ;
        RECT 1174.020 620.510 1174.280 620.830 ;
        RECT 1174.020 572.570 1174.280 572.890 ;
        RECT 1174.080 531.490 1174.220 572.570 ;
        RECT 1174.080 531.350 1174.680 531.490 ;
        RECT 1174.540 507.010 1174.680 531.350 ;
        RECT 1174.080 506.870 1174.680 507.010 ;
        RECT 1174.080 435.725 1174.220 506.870 ;
        RECT 1174.010 435.355 1174.290 435.725 ;
        RECT 1173.550 434.675 1173.830 435.045 ;
        RECT 1173.620 386.570 1173.760 434.675 ;
        RECT 1173.560 386.250 1173.820 386.570 ;
        RECT 1174.020 386.250 1174.280 386.570 ;
        RECT 1174.080 254.730 1174.220 386.250 ;
        RECT 1174.080 254.590 1174.680 254.730 ;
        RECT 1174.540 241.390 1174.680 254.590 ;
        RECT 1174.480 241.070 1174.740 241.390 ;
        RECT 1174.020 193.130 1174.280 193.450 ;
        RECT 1174.080 169.050 1174.220 193.130 ;
        RECT 1173.620 168.910 1174.220 169.050 ;
        RECT 1173.620 96.890 1173.760 168.910 ;
        RECT 1173.560 96.570 1173.820 96.890 ;
        RECT 1174.020 96.570 1174.280 96.890 ;
        RECT 1174.080 25.830 1174.220 96.570 ;
        RECT 835.920 25.510 836.180 25.830 ;
        RECT 1174.020 25.510 1174.280 25.830 ;
        RECT 835.980 7.210 836.120 25.510 ;
        RECT 835.520 7.070 836.120 7.210 ;
        RECT 835.520 2.400 835.660 7.070 ;
        RECT 835.310 -4.800 835.870 2.400 ;
      LAYER via2 ;
        RECT 1174.010 965.800 1174.290 966.080 ;
        RECT 1174.930 965.800 1175.210 966.080 ;
        RECT 1174.010 814.160 1174.290 814.440 ;
        RECT 1174.930 814.160 1175.210 814.440 ;
        RECT 1174.010 676.120 1174.290 676.400 ;
        RECT 1174.930 676.120 1175.210 676.400 ;
        RECT 1174.010 435.400 1174.290 435.680 ;
        RECT 1173.550 434.720 1173.830 435.000 ;
      LAYER met3 ;
        RECT 1173.985 966.090 1174.315 966.105 ;
        RECT 1174.905 966.090 1175.235 966.105 ;
        RECT 1173.985 965.790 1175.235 966.090 ;
        RECT 1173.985 965.775 1174.315 965.790 ;
        RECT 1174.905 965.775 1175.235 965.790 ;
        RECT 1173.985 814.450 1174.315 814.465 ;
        RECT 1174.905 814.450 1175.235 814.465 ;
        RECT 1173.985 814.150 1175.235 814.450 ;
        RECT 1173.985 814.135 1174.315 814.150 ;
        RECT 1174.905 814.135 1175.235 814.150 ;
        RECT 1173.985 676.410 1174.315 676.425 ;
        RECT 1174.905 676.410 1175.235 676.425 ;
        RECT 1173.985 676.110 1175.235 676.410 ;
        RECT 1173.985 676.095 1174.315 676.110 ;
        RECT 1174.905 676.095 1175.235 676.110 ;
        RECT 1173.985 435.690 1174.315 435.705 ;
        RECT 1173.310 435.390 1174.315 435.690 ;
        RECT 1173.310 435.025 1173.610 435.390 ;
        RECT 1173.985 435.375 1174.315 435.390 ;
        RECT 1173.310 434.710 1173.855 435.025 ;
        RECT 1173.525 434.695 1173.855 434.710 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2179.550 38.660 2179.870 38.720 ;
        RECT 2779.850 38.660 2780.170 38.720 ;
        RECT 2179.550 38.520 2780.170 38.660 ;
        RECT 2179.550 38.460 2179.870 38.520 ;
        RECT 2779.850 38.460 2780.170 38.520 ;
      LAYER via ;
        RECT 2179.580 38.460 2179.840 38.720 ;
        RECT 2779.880 38.460 2780.140 38.720 ;
      LAYER met2 ;
        RECT 2177.750 1220.330 2178.310 1228.680 ;
        RECT 2177.750 1220.190 2179.780 1220.330 ;
        RECT 2177.750 1219.680 2178.310 1220.190 ;
        RECT 2179.640 38.750 2179.780 1220.190 ;
        RECT 2179.580 38.430 2179.840 38.750 ;
        RECT 2779.880 38.430 2780.140 38.750 ;
        RECT 2779.940 2.400 2780.080 38.430 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2186.450 38.320 2186.770 38.380 ;
        RECT 2797.790 38.320 2798.110 38.380 ;
        RECT 2186.450 38.180 2798.110 38.320 ;
        RECT 2186.450 38.120 2186.770 38.180 ;
        RECT 2797.790 38.120 2798.110 38.180 ;
      LAYER via ;
        RECT 2186.480 38.120 2186.740 38.380 ;
        RECT 2797.820 38.120 2798.080 38.380 ;
      LAYER met2 ;
        RECT 2186.950 1220.330 2187.510 1228.680 ;
        RECT 2186.540 1220.190 2187.510 1220.330 ;
        RECT 2186.540 38.410 2186.680 1220.190 ;
        RECT 2186.950 1219.680 2187.510 1220.190 ;
        RECT 2186.480 38.090 2186.740 38.410 ;
        RECT 2797.820 38.090 2798.080 38.410 ;
        RECT 2797.880 2.400 2798.020 38.090 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2196.110 1207.580 2196.430 1207.640 ;
        RECT 2200.710 1207.580 2201.030 1207.640 ;
        RECT 2196.110 1207.440 2201.030 1207.580 ;
        RECT 2196.110 1207.380 2196.430 1207.440 ;
        RECT 2200.710 1207.380 2201.030 1207.440 ;
      LAYER via ;
        RECT 2196.140 1207.380 2196.400 1207.640 ;
        RECT 2200.740 1207.380 2201.000 1207.640 ;
      LAYER met2 ;
        RECT 2196.150 1219.680 2196.710 1228.680 ;
        RECT 2196.200 1207.670 2196.340 1219.680 ;
        RECT 2196.140 1207.350 2196.400 1207.670 ;
        RECT 2200.740 1207.350 2201.000 1207.670 ;
        RECT 2200.800 31.125 2200.940 1207.350 ;
        RECT 2200.730 30.755 2201.010 31.125 ;
        RECT 2815.750 30.755 2816.030 31.125 ;
        RECT 2815.820 2.400 2815.960 30.755 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 2200.730 30.800 2201.010 31.080 ;
        RECT 2815.750 30.800 2816.030 31.080 ;
      LAYER met3 ;
        RECT 2200.705 31.090 2201.035 31.105 ;
        RECT 2815.725 31.090 2816.055 31.105 ;
        RECT 2200.705 30.790 2816.055 31.090 ;
        RECT 2200.705 30.775 2201.035 30.790 ;
        RECT 2815.725 30.775 2816.055 30.790 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2207.150 37.980 2207.470 38.040 ;
        RECT 2833.670 37.980 2833.990 38.040 ;
        RECT 2207.150 37.840 2833.990 37.980 ;
        RECT 2207.150 37.780 2207.470 37.840 ;
        RECT 2833.670 37.780 2833.990 37.840 ;
      LAYER via ;
        RECT 2207.180 37.780 2207.440 38.040 ;
        RECT 2833.700 37.780 2833.960 38.040 ;
      LAYER met2 ;
        RECT 2205.350 1220.330 2205.910 1228.680 ;
        RECT 2205.350 1220.190 2207.380 1220.330 ;
        RECT 2205.350 1219.680 2205.910 1220.190 ;
        RECT 2207.240 38.070 2207.380 1220.190 ;
        RECT 2207.180 37.750 2207.440 38.070 ;
        RECT 2833.700 37.750 2833.960 38.070 ;
        RECT 2833.760 2.400 2833.900 37.750 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2213.590 1210.300 2213.910 1210.360 ;
        RECT 2214.510 1210.300 2214.830 1210.360 ;
        RECT 2213.590 1210.160 2214.830 1210.300 ;
        RECT 2213.590 1210.100 2213.910 1210.160 ;
        RECT 2214.510 1210.100 2214.830 1210.160 ;
      LAYER via ;
        RECT 2213.620 1210.100 2213.880 1210.360 ;
        RECT 2214.540 1210.100 2214.800 1210.360 ;
      LAYER met2 ;
        RECT 2214.550 1219.680 2215.110 1228.680 ;
        RECT 2214.600 1210.390 2214.740 1219.680 ;
        RECT 2213.620 1210.070 2213.880 1210.390 ;
        RECT 2214.540 1210.070 2214.800 1210.390 ;
        RECT 2213.680 37.925 2213.820 1210.070 ;
        RECT 2213.610 37.555 2213.890 37.925 ;
        RECT 2851.170 37.555 2851.450 37.925 ;
        RECT 2851.240 2.400 2851.380 37.555 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
      LAYER via2 ;
        RECT 2213.610 37.600 2213.890 37.880 ;
        RECT 2851.170 37.600 2851.450 37.880 ;
      LAYER met3 ;
        RECT 2213.585 37.890 2213.915 37.905 ;
        RECT 2851.145 37.890 2851.475 37.905 ;
        RECT 2213.585 37.590 2851.475 37.890 ;
        RECT 2213.585 37.575 2213.915 37.590 ;
        RECT 2851.145 37.575 2851.475 37.590 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2223.710 1210.300 2224.030 1210.360 ;
        RECT 2227.850 1210.300 2228.170 1210.360 ;
        RECT 2223.710 1210.160 2228.170 1210.300 ;
        RECT 2223.710 1210.100 2224.030 1210.160 ;
        RECT 2227.850 1210.100 2228.170 1210.160 ;
        RECT 2227.850 45.460 2228.170 45.520 ;
        RECT 2869.090 45.460 2869.410 45.520 ;
        RECT 2227.850 45.320 2869.410 45.460 ;
        RECT 2227.850 45.260 2228.170 45.320 ;
        RECT 2869.090 45.260 2869.410 45.320 ;
      LAYER via ;
        RECT 2223.740 1210.100 2224.000 1210.360 ;
        RECT 2227.880 1210.100 2228.140 1210.360 ;
        RECT 2227.880 45.260 2228.140 45.520 ;
        RECT 2869.120 45.260 2869.380 45.520 ;
      LAYER met2 ;
        RECT 2223.750 1219.680 2224.310 1228.680 ;
        RECT 2223.800 1210.390 2223.940 1219.680 ;
        RECT 2223.740 1210.070 2224.000 1210.390 ;
        RECT 2227.880 1210.070 2228.140 1210.390 ;
        RECT 2227.940 45.550 2228.080 1210.070 ;
        RECT 2227.880 45.230 2228.140 45.550 ;
        RECT 2869.120 45.230 2869.380 45.550 ;
        RECT 2869.180 2.400 2869.320 45.230 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2234.750 45.120 2235.070 45.180 ;
        RECT 2887.030 45.120 2887.350 45.180 ;
        RECT 2234.750 44.980 2887.350 45.120 ;
        RECT 2234.750 44.920 2235.070 44.980 ;
        RECT 2887.030 44.920 2887.350 44.980 ;
      LAYER via ;
        RECT 2234.780 44.920 2235.040 45.180 ;
        RECT 2887.060 44.920 2887.320 45.180 ;
      LAYER met2 ;
        RECT 2232.950 1220.330 2233.510 1228.680 ;
        RECT 2232.950 1220.190 2234.980 1220.330 ;
        RECT 2232.950 1219.680 2233.510 1220.190 ;
        RECT 2234.840 45.210 2234.980 1220.190 ;
        RECT 2234.780 44.890 2235.040 45.210 ;
        RECT 2887.060 44.890 2887.320 45.210 ;
        RECT 2887.120 2.400 2887.260 44.890 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2241.650 44.780 2241.970 44.840 ;
        RECT 2904.970 44.780 2905.290 44.840 ;
        RECT 2241.650 44.640 2905.290 44.780 ;
        RECT 2241.650 44.580 2241.970 44.640 ;
        RECT 2904.970 44.580 2905.290 44.640 ;
      LAYER via ;
        RECT 2241.680 44.580 2241.940 44.840 ;
        RECT 2905.000 44.580 2905.260 44.840 ;
      LAYER met2 ;
        RECT 2242.150 1220.330 2242.710 1228.680 ;
        RECT 2241.740 1220.190 2242.710 1220.330 ;
        RECT 2241.740 44.870 2241.880 1220.190 ;
        RECT 2242.150 1219.680 2242.710 1220.190 ;
        RECT 2241.680 44.550 2241.940 44.870 ;
        RECT 2905.000 44.550 2905.260 44.870 ;
        RECT 2905.060 2.400 2905.200 44.550 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 852.910 26.080 853.230 26.140 ;
        RECT 1186.870 26.080 1187.190 26.140 ;
        RECT 852.910 25.940 1187.190 26.080 ;
        RECT 852.910 25.880 853.230 25.940 ;
        RECT 1186.870 25.880 1187.190 25.940 ;
      LAYER via ;
        RECT 852.940 25.880 853.200 26.140 ;
        RECT 1186.900 25.880 1187.160 26.140 ;
      LAYER met2 ;
        RECT 1187.830 1220.330 1188.390 1228.680 ;
        RECT 1186.960 1220.190 1188.390 1220.330 ;
        RECT 1186.960 26.170 1187.100 1220.190 ;
        RECT 1187.830 1219.680 1188.390 1220.190 ;
        RECT 852.940 25.850 853.200 26.170 ;
        RECT 1186.900 25.850 1187.160 26.170 ;
        RECT 853.000 2.400 853.140 25.850 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 907.265 26.265 907.435 27.115 ;
      LAYER mcon ;
        RECT 907.265 26.945 907.435 27.115 ;
      LAYER met1 ;
        RECT 870.850 27.100 871.170 27.160 ;
        RECT 907.205 27.100 907.495 27.145 ;
        RECT 870.850 26.960 907.495 27.100 ;
        RECT 870.850 26.900 871.170 26.960 ;
        RECT 907.205 26.915 907.495 26.960 ;
        RECT 907.205 26.420 907.495 26.465 ;
        RECT 1194.230 26.420 1194.550 26.480 ;
        RECT 907.205 26.280 1194.550 26.420 ;
        RECT 907.205 26.235 907.495 26.280 ;
        RECT 1194.230 26.220 1194.550 26.280 ;
      LAYER via ;
        RECT 870.880 26.900 871.140 27.160 ;
        RECT 1194.260 26.220 1194.520 26.480 ;
      LAYER met2 ;
        RECT 1197.030 1220.330 1197.590 1228.680 ;
        RECT 1195.700 1220.190 1197.590 1220.330 ;
        RECT 1195.700 1197.210 1195.840 1220.190 ;
        RECT 1197.030 1219.680 1197.590 1220.190 ;
        RECT 1194.320 1197.070 1195.840 1197.210 ;
        RECT 870.880 26.870 871.140 27.190 ;
        RECT 870.940 2.400 871.080 26.870 ;
        RECT 1194.320 26.510 1194.460 1197.070 ;
        RECT 1194.260 26.190 1194.520 26.510 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1024.490 1209.280 1024.810 1209.340 ;
        RECT 1206.190 1209.280 1206.510 1209.340 ;
        RECT 1024.490 1209.140 1206.510 1209.280 ;
        RECT 1024.490 1209.080 1024.810 1209.140 ;
        RECT 1206.190 1209.080 1206.510 1209.140 ;
        RECT 888.790 19.620 889.110 19.680 ;
        RECT 888.790 19.480 908.340 19.620 ;
        RECT 888.790 19.420 889.110 19.480 ;
        RECT 908.200 19.280 908.340 19.480 ;
        RECT 1024.490 19.280 1024.810 19.340 ;
        RECT 908.200 19.140 1024.810 19.280 ;
        RECT 1024.490 19.080 1024.810 19.140 ;
      LAYER via ;
        RECT 1024.520 1209.080 1024.780 1209.340 ;
        RECT 1206.220 1209.080 1206.480 1209.340 ;
        RECT 888.820 19.420 889.080 19.680 ;
        RECT 1024.520 19.080 1024.780 19.340 ;
      LAYER met2 ;
        RECT 1206.230 1219.680 1206.790 1228.680 ;
        RECT 1206.280 1209.370 1206.420 1219.680 ;
        RECT 1024.520 1209.050 1024.780 1209.370 ;
        RECT 1206.220 1209.050 1206.480 1209.370 ;
        RECT 888.820 19.390 889.080 19.710 ;
        RECT 888.880 2.400 889.020 19.390 ;
        RECT 1024.580 19.370 1024.720 1209.050 ;
        RECT 1024.520 19.050 1024.780 19.370 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 907.650 27.100 907.970 27.160 ;
        RECT 907.650 26.960 908.340 27.100 ;
        RECT 907.650 26.900 907.970 26.960 ;
        RECT 908.200 26.760 908.340 26.960 ;
        RECT 1214.930 26.760 1215.250 26.820 ;
        RECT 908.200 26.620 1215.250 26.760 ;
        RECT 1214.930 26.560 1215.250 26.620 ;
      LAYER via ;
        RECT 907.680 26.900 907.940 27.160 ;
        RECT 1214.960 26.560 1215.220 26.820 ;
      LAYER met2 ;
        RECT 1215.430 1220.330 1215.990 1228.680 ;
        RECT 1215.020 1220.190 1215.990 1220.330 ;
        RECT 907.680 26.870 907.940 27.190 ;
        RECT 907.740 14.010 907.880 26.870 ;
        RECT 1215.020 26.850 1215.160 1220.190 ;
        RECT 1215.430 1219.680 1215.990 1220.190 ;
        RECT 1214.960 26.530 1215.220 26.850 ;
        RECT 906.820 13.870 907.880 14.010 ;
        RECT 906.820 2.400 906.960 13.870 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 955.565 23.205 955.735 27.115 ;
      LAYER mcon ;
        RECT 955.565 26.945 955.735 27.115 ;
      LAYER met1 ;
        RECT 1221.830 1196.700 1222.150 1196.760 ;
        RECT 1222.750 1196.700 1223.070 1196.760 ;
        RECT 1221.830 1196.560 1223.070 1196.700 ;
        RECT 1221.830 1196.500 1222.150 1196.560 ;
        RECT 1222.750 1196.500 1223.070 1196.560 ;
        RECT 955.505 27.100 955.795 27.145 ;
        RECT 1221.830 27.100 1222.150 27.160 ;
        RECT 955.505 26.960 1222.150 27.100 ;
        RECT 955.505 26.915 955.795 26.960 ;
        RECT 1221.830 26.900 1222.150 26.960 ;
        RECT 924.210 23.360 924.530 23.420 ;
        RECT 955.505 23.360 955.795 23.405 ;
        RECT 924.210 23.220 955.795 23.360 ;
        RECT 924.210 23.160 924.530 23.220 ;
        RECT 955.505 23.175 955.795 23.220 ;
      LAYER via ;
        RECT 1221.860 1196.500 1222.120 1196.760 ;
        RECT 1222.780 1196.500 1223.040 1196.760 ;
        RECT 1221.860 26.900 1222.120 27.160 ;
        RECT 924.240 23.160 924.500 23.420 ;
      LAYER met2 ;
        RECT 1224.630 1220.330 1225.190 1228.680 ;
        RECT 1222.840 1220.190 1225.190 1220.330 ;
        RECT 1222.840 1196.790 1222.980 1220.190 ;
        RECT 1224.630 1219.680 1225.190 1220.190 ;
        RECT 1221.860 1196.470 1222.120 1196.790 ;
        RECT 1222.780 1196.470 1223.040 1196.790 ;
        RECT 1221.920 27.190 1222.060 1196.470 ;
        RECT 1221.860 26.870 1222.120 27.190 ;
        RECT 924.240 23.130 924.500 23.450 ;
        RECT 924.300 2.400 924.440 23.130 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1228.805 620.925 1228.975 669.375 ;
        RECT 1228.805 524.365 1228.975 548.675 ;
        RECT 1228.805 415.905 1228.975 452.115 ;
        RECT 1230.185 324.445 1230.355 372.555 ;
        RECT 1228.805 138.125 1228.975 227.715 ;
        RECT 1229.265 96.645 1229.435 136.255 ;
      LAYER mcon ;
        RECT 1228.805 669.205 1228.975 669.375 ;
        RECT 1228.805 548.505 1228.975 548.675 ;
        RECT 1228.805 451.945 1228.975 452.115 ;
        RECT 1230.185 372.385 1230.355 372.555 ;
        RECT 1228.805 227.545 1228.975 227.715 ;
        RECT 1229.265 136.085 1229.435 136.255 ;
      LAYER met1 ;
        RECT 1229.650 1173.240 1229.970 1173.300 ;
        RECT 1232.410 1173.240 1232.730 1173.300 ;
        RECT 1229.650 1173.100 1232.730 1173.240 ;
        RECT 1229.650 1173.040 1229.970 1173.100 ;
        RECT 1232.410 1173.040 1232.730 1173.100 ;
        RECT 1229.650 1125.300 1229.970 1125.360 ;
        RECT 1229.280 1125.160 1229.970 1125.300 ;
        RECT 1229.280 1124.680 1229.420 1125.160 ;
        RECT 1229.650 1125.100 1229.970 1125.160 ;
        RECT 1229.190 1124.420 1229.510 1124.680 ;
        RECT 1229.190 1110.480 1229.510 1110.740 ;
        RECT 1229.280 1110.000 1229.420 1110.480 ;
        RECT 1229.650 1110.000 1229.970 1110.060 ;
        RECT 1229.280 1109.860 1229.970 1110.000 ;
        RECT 1229.650 1109.800 1229.970 1109.860 ;
        RECT 1229.650 966.180 1229.970 966.240 ;
        RECT 1230.570 966.180 1230.890 966.240 ;
        RECT 1229.650 966.040 1230.890 966.180 ;
        RECT 1229.650 965.980 1229.970 966.040 ;
        RECT 1230.570 965.980 1230.890 966.040 ;
        RECT 1229.650 869.620 1229.970 869.680 ;
        RECT 1230.570 869.620 1230.890 869.680 ;
        RECT 1229.650 869.480 1230.890 869.620 ;
        RECT 1229.650 869.420 1229.970 869.480 ;
        RECT 1230.570 869.420 1230.890 869.480 ;
        RECT 1228.730 717.440 1229.050 717.700 ;
        RECT 1228.820 717.300 1228.960 717.440 ;
        RECT 1229.650 717.300 1229.970 717.360 ;
        RECT 1228.820 717.160 1229.970 717.300 ;
        RECT 1229.650 717.100 1229.970 717.160 ;
        RECT 1228.745 669.360 1229.035 669.405 ;
        RECT 1229.650 669.360 1229.970 669.420 ;
        RECT 1228.745 669.220 1229.970 669.360 ;
        RECT 1228.745 669.175 1229.035 669.220 ;
        RECT 1229.650 669.160 1229.970 669.220 ;
        RECT 1228.730 621.080 1229.050 621.140 ;
        RECT 1228.535 620.940 1229.050 621.080 ;
        RECT 1228.730 620.880 1229.050 620.940 ;
        RECT 1228.745 548.660 1229.035 548.705 ;
        RECT 1229.650 548.660 1229.970 548.720 ;
        RECT 1228.745 548.520 1229.970 548.660 ;
        RECT 1228.745 548.475 1229.035 548.520 ;
        RECT 1229.650 548.460 1229.970 548.520 ;
        RECT 1228.730 524.520 1229.050 524.580 ;
        RECT 1228.535 524.380 1229.050 524.520 ;
        RECT 1228.730 524.320 1229.050 524.380 ;
        RECT 1228.745 452.100 1229.035 452.145 ;
        RECT 1229.650 452.100 1229.970 452.160 ;
        RECT 1228.745 451.960 1229.970 452.100 ;
        RECT 1228.745 451.915 1229.035 451.960 ;
        RECT 1229.650 451.900 1229.970 451.960 ;
        RECT 1228.745 416.060 1229.035 416.105 ;
        RECT 1231.030 416.060 1231.350 416.120 ;
        RECT 1228.745 415.920 1231.350 416.060 ;
        RECT 1228.745 415.875 1229.035 415.920 ;
        RECT 1231.030 415.860 1231.350 415.920 ;
        RECT 1230.125 372.540 1230.415 372.585 ;
        RECT 1231.030 372.540 1231.350 372.600 ;
        RECT 1230.125 372.400 1231.350 372.540 ;
        RECT 1230.125 372.355 1230.415 372.400 ;
        RECT 1231.030 372.340 1231.350 372.400 ;
        RECT 1230.110 324.600 1230.430 324.660 ;
        RECT 1229.915 324.460 1230.430 324.600 ;
        RECT 1230.110 324.400 1230.430 324.460 ;
        RECT 1230.110 283.460 1230.430 283.520 ;
        RECT 1229.280 283.320 1230.430 283.460 ;
        RECT 1229.280 282.840 1229.420 283.320 ;
        RECT 1230.110 283.260 1230.430 283.320 ;
        RECT 1229.190 282.580 1229.510 282.840 ;
        RECT 1229.190 234.300 1229.510 234.560 ;
        RECT 1228.730 234.160 1229.050 234.220 ;
        RECT 1229.280 234.160 1229.420 234.300 ;
        RECT 1228.730 234.020 1229.420 234.160 ;
        RECT 1228.730 233.960 1229.050 234.020 ;
        RECT 1228.730 227.700 1229.050 227.760 ;
        RECT 1228.535 227.560 1229.050 227.700 ;
        RECT 1228.730 227.500 1229.050 227.560 ;
        RECT 1228.745 138.280 1229.035 138.325 ;
        RECT 1229.190 138.280 1229.510 138.340 ;
        RECT 1228.745 138.140 1229.510 138.280 ;
        RECT 1228.745 138.095 1229.035 138.140 ;
        RECT 1229.190 138.080 1229.510 138.140 ;
        RECT 1229.190 136.240 1229.510 136.300 ;
        RECT 1228.995 136.100 1229.510 136.240 ;
        RECT 1229.190 136.040 1229.510 136.100 ;
        RECT 1229.205 96.800 1229.495 96.845 ;
        RECT 1229.650 96.800 1229.970 96.860 ;
        RECT 1229.205 96.660 1229.970 96.800 ;
        RECT 1229.205 96.615 1229.495 96.660 ;
        RECT 1229.650 96.600 1229.970 96.660 ;
        RECT 942.150 23.700 942.470 23.760 ;
        RECT 1229.650 23.700 1229.970 23.760 ;
        RECT 942.150 23.560 1229.970 23.700 ;
        RECT 942.150 23.500 942.470 23.560 ;
        RECT 1229.650 23.500 1229.970 23.560 ;
      LAYER via ;
        RECT 1229.680 1173.040 1229.940 1173.300 ;
        RECT 1232.440 1173.040 1232.700 1173.300 ;
        RECT 1229.680 1125.100 1229.940 1125.360 ;
        RECT 1229.220 1124.420 1229.480 1124.680 ;
        RECT 1229.220 1110.480 1229.480 1110.740 ;
        RECT 1229.680 1109.800 1229.940 1110.060 ;
        RECT 1229.680 965.980 1229.940 966.240 ;
        RECT 1230.600 965.980 1230.860 966.240 ;
        RECT 1229.680 869.420 1229.940 869.680 ;
        RECT 1230.600 869.420 1230.860 869.680 ;
        RECT 1228.760 717.440 1229.020 717.700 ;
        RECT 1229.680 717.100 1229.940 717.360 ;
        RECT 1229.680 669.160 1229.940 669.420 ;
        RECT 1228.760 620.880 1229.020 621.140 ;
        RECT 1229.680 548.460 1229.940 548.720 ;
        RECT 1228.760 524.320 1229.020 524.580 ;
        RECT 1229.680 451.900 1229.940 452.160 ;
        RECT 1231.060 415.860 1231.320 416.120 ;
        RECT 1231.060 372.340 1231.320 372.600 ;
        RECT 1230.140 324.400 1230.400 324.660 ;
        RECT 1230.140 283.260 1230.400 283.520 ;
        RECT 1229.220 282.580 1229.480 282.840 ;
        RECT 1229.220 234.300 1229.480 234.560 ;
        RECT 1228.760 233.960 1229.020 234.220 ;
        RECT 1228.760 227.500 1229.020 227.760 ;
        RECT 1229.220 138.080 1229.480 138.340 ;
        RECT 1229.220 136.040 1229.480 136.300 ;
        RECT 1229.680 96.600 1229.940 96.860 ;
        RECT 942.180 23.500 942.440 23.760 ;
        RECT 1229.680 23.500 1229.940 23.760 ;
      LAYER met2 ;
        RECT 1233.830 1220.330 1234.390 1228.680 ;
        RECT 1232.500 1220.190 1234.390 1220.330 ;
        RECT 1232.500 1173.330 1232.640 1220.190 ;
        RECT 1233.830 1219.680 1234.390 1220.190 ;
        RECT 1229.680 1173.010 1229.940 1173.330 ;
        RECT 1232.440 1173.010 1232.700 1173.330 ;
        RECT 1229.740 1125.390 1229.880 1173.010 ;
        RECT 1229.680 1125.070 1229.940 1125.390 ;
        RECT 1229.220 1124.390 1229.480 1124.710 ;
        RECT 1229.280 1110.770 1229.420 1124.390 ;
        RECT 1229.220 1110.450 1229.480 1110.770 ;
        RECT 1229.680 1109.770 1229.940 1110.090 ;
        RECT 1229.740 1027.890 1229.880 1109.770 ;
        RECT 1229.280 1027.750 1229.880 1027.890 ;
        RECT 1229.280 1014.405 1229.420 1027.750 ;
        RECT 1229.210 1014.035 1229.490 1014.405 ;
        RECT 1230.590 1014.035 1230.870 1014.405 ;
        RECT 1230.660 966.270 1230.800 1014.035 ;
        RECT 1229.680 965.950 1229.940 966.270 ;
        RECT 1230.600 965.950 1230.860 966.270 ;
        RECT 1229.740 931.330 1229.880 965.950 ;
        RECT 1229.280 931.190 1229.880 931.330 ;
        RECT 1229.280 917.845 1229.420 931.190 ;
        RECT 1229.210 917.475 1229.490 917.845 ;
        RECT 1230.590 917.475 1230.870 917.845 ;
        RECT 1230.660 869.710 1230.800 917.475 ;
        RECT 1229.680 869.390 1229.940 869.710 ;
        RECT 1230.600 869.390 1230.860 869.710 ;
        RECT 1229.740 834.770 1229.880 869.390 ;
        RECT 1229.280 834.630 1229.880 834.770 ;
        RECT 1229.280 772.210 1229.420 834.630 ;
        RECT 1228.820 772.070 1229.420 772.210 ;
        RECT 1228.820 717.730 1228.960 772.070 ;
        RECT 1228.760 717.410 1229.020 717.730 ;
        RECT 1229.680 717.070 1229.940 717.390 ;
        RECT 1229.740 692.650 1229.880 717.070 ;
        RECT 1229.280 692.510 1229.880 692.650 ;
        RECT 1229.280 669.530 1229.420 692.510 ;
        RECT 1229.280 669.450 1229.880 669.530 ;
        RECT 1229.280 669.390 1229.940 669.450 ;
        RECT 1229.680 669.130 1229.940 669.390 ;
        RECT 1229.740 668.975 1229.880 669.130 ;
        RECT 1228.760 620.850 1229.020 621.170 ;
        RECT 1228.820 573.765 1228.960 620.850 ;
        RECT 1228.750 573.395 1229.030 573.765 ;
        RECT 1229.670 572.715 1229.950 573.085 ;
        RECT 1229.740 548.750 1229.880 572.715 ;
        RECT 1229.680 548.430 1229.940 548.750 ;
        RECT 1228.760 524.290 1229.020 524.610 ;
        RECT 1228.820 477.205 1228.960 524.290 ;
        RECT 1228.750 476.835 1229.030 477.205 ;
        RECT 1229.670 476.155 1229.950 476.525 ;
        RECT 1229.740 452.190 1229.880 476.155 ;
        RECT 1229.680 451.870 1229.940 452.190 ;
        RECT 1231.060 415.830 1231.320 416.150 ;
        RECT 1231.120 372.630 1231.260 415.830 ;
        RECT 1231.060 372.310 1231.320 372.630 ;
        RECT 1230.140 324.370 1230.400 324.690 ;
        RECT 1230.200 283.550 1230.340 324.370 ;
        RECT 1230.140 283.230 1230.400 283.550 ;
        RECT 1229.220 282.550 1229.480 282.870 ;
        RECT 1229.280 234.590 1229.420 282.550 ;
        RECT 1229.220 234.270 1229.480 234.590 ;
        RECT 1228.760 233.930 1229.020 234.250 ;
        RECT 1228.820 227.790 1228.960 233.930 ;
        RECT 1228.760 227.470 1229.020 227.790 ;
        RECT 1229.220 138.050 1229.480 138.370 ;
        RECT 1229.280 136.330 1229.420 138.050 ;
        RECT 1229.220 136.010 1229.480 136.330 ;
        RECT 1229.680 96.570 1229.940 96.890 ;
        RECT 1229.740 23.790 1229.880 96.570 ;
        RECT 942.180 23.470 942.440 23.790 ;
        RECT 1229.680 23.470 1229.940 23.790 ;
        RECT 942.240 2.400 942.380 23.470 ;
        RECT 942.030 -4.800 942.590 2.400 ;
      LAYER via2 ;
        RECT 1229.210 1014.080 1229.490 1014.360 ;
        RECT 1230.590 1014.080 1230.870 1014.360 ;
        RECT 1229.210 917.520 1229.490 917.800 ;
        RECT 1230.590 917.520 1230.870 917.800 ;
        RECT 1228.750 573.440 1229.030 573.720 ;
        RECT 1229.670 572.760 1229.950 573.040 ;
        RECT 1228.750 476.880 1229.030 477.160 ;
        RECT 1229.670 476.200 1229.950 476.480 ;
      LAYER met3 ;
        RECT 1229.185 1014.370 1229.515 1014.385 ;
        RECT 1230.565 1014.370 1230.895 1014.385 ;
        RECT 1229.185 1014.070 1230.895 1014.370 ;
        RECT 1229.185 1014.055 1229.515 1014.070 ;
        RECT 1230.565 1014.055 1230.895 1014.070 ;
        RECT 1229.185 917.810 1229.515 917.825 ;
        RECT 1230.565 917.810 1230.895 917.825 ;
        RECT 1229.185 917.510 1230.895 917.810 ;
        RECT 1229.185 917.495 1229.515 917.510 ;
        RECT 1230.565 917.495 1230.895 917.510 ;
        RECT 1228.725 573.730 1229.055 573.745 ;
        RECT 1228.725 573.430 1230.650 573.730 ;
        RECT 1228.725 573.415 1229.055 573.430 ;
        RECT 1229.645 573.050 1229.975 573.065 ;
        RECT 1230.350 573.050 1230.650 573.430 ;
        RECT 1229.645 572.750 1230.650 573.050 ;
        RECT 1229.645 572.735 1229.975 572.750 ;
        RECT 1228.725 477.170 1229.055 477.185 ;
        RECT 1228.725 476.870 1230.650 477.170 ;
        RECT 1228.725 476.855 1229.055 476.870 ;
        RECT 1229.645 476.490 1229.975 476.505 ;
        RECT 1230.350 476.490 1230.650 476.870 ;
        RECT 1229.645 476.190 1230.650 476.490 ;
        RECT 1229.645 476.175 1229.975 476.190 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 23.020 960.410 23.080 ;
        RECT 1242.530 23.020 1242.850 23.080 ;
        RECT 960.090 22.880 1242.850 23.020 ;
        RECT 960.090 22.820 960.410 22.880 ;
        RECT 1242.530 22.820 1242.850 22.880 ;
      LAYER via ;
        RECT 960.120 22.820 960.380 23.080 ;
        RECT 1242.560 22.820 1242.820 23.080 ;
      LAYER met2 ;
        RECT 1243.030 1220.330 1243.590 1228.680 ;
        RECT 1242.620 1220.190 1243.590 1220.330 ;
        RECT 1242.620 23.110 1242.760 1220.190 ;
        RECT 1243.030 1219.680 1243.590 1220.190 ;
        RECT 960.120 22.790 960.380 23.110 ;
        RECT 1242.560 22.790 1242.820 23.110 ;
        RECT 960.180 2.400 960.320 22.790 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1249.430 1196.700 1249.750 1196.760 ;
        RECT 1250.350 1196.700 1250.670 1196.760 ;
        RECT 1249.430 1196.560 1250.670 1196.700 ;
        RECT 1249.430 1196.500 1249.750 1196.560 ;
        RECT 1250.350 1196.500 1250.670 1196.560 ;
        RECT 978.030 22.340 978.350 22.400 ;
        RECT 1249.430 22.340 1249.750 22.400 ;
        RECT 978.030 22.200 1249.750 22.340 ;
        RECT 978.030 22.140 978.350 22.200 ;
        RECT 1249.430 22.140 1249.750 22.200 ;
      LAYER via ;
        RECT 1249.460 1196.500 1249.720 1196.760 ;
        RECT 1250.380 1196.500 1250.640 1196.760 ;
        RECT 978.060 22.140 978.320 22.400 ;
        RECT 1249.460 22.140 1249.720 22.400 ;
      LAYER met2 ;
        RECT 1252.230 1220.330 1252.790 1228.680 ;
        RECT 1250.440 1220.190 1252.790 1220.330 ;
        RECT 1250.440 1196.790 1250.580 1220.190 ;
        RECT 1252.230 1219.680 1252.790 1220.190 ;
        RECT 1249.460 1196.470 1249.720 1196.790 ;
        RECT 1250.380 1196.470 1250.640 1196.790 ;
        RECT 1249.520 22.430 1249.660 1196.470 ;
        RECT 978.060 22.110 978.320 22.430 ;
        RECT 1249.460 22.110 1249.720 22.430 ;
        RECT 978.120 2.400 978.260 22.110 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1084.825 1055.445 1084.995 1097.095 ;
        RECT 1083.905 758.965 1084.075 807.075 ;
        RECT 1083.905 648.465 1084.075 676.175 ;
        RECT 1084.365 427.805 1084.535 475.915 ;
        RECT 1084.825 227.885 1084.995 275.995 ;
      LAYER mcon ;
        RECT 1084.825 1096.925 1084.995 1097.095 ;
        RECT 1083.905 806.905 1084.075 807.075 ;
        RECT 1083.905 676.005 1084.075 676.175 ;
        RECT 1084.365 475.745 1084.535 475.915 ;
        RECT 1084.825 275.825 1084.995 275.995 ;
      LAYER met1 ;
        RECT 1083.830 1104.560 1084.150 1104.620 ;
        RECT 1084.290 1104.560 1084.610 1104.620 ;
        RECT 1083.830 1104.420 1084.610 1104.560 ;
        RECT 1083.830 1104.360 1084.150 1104.420 ;
        RECT 1084.290 1104.360 1084.610 1104.420 ;
        RECT 1083.830 1103.880 1084.150 1103.940 ;
        RECT 1084.750 1103.880 1085.070 1103.940 ;
        RECT 1083.830 1103.740 1085.070 1103.880 ;
        RECT 1083.830 1103.680 1084.150 1103.740 ;
        RECT 1084.750 1103.680 1085.070 1103.740 ;
        RECT 1084.750 1097.080 1085.070 1097.140 ;
        RECT 1084.555 1096.940 1085.070 1097.080 ;
        RECT 1084.750 1096.880 1085.070 1096.940 ;
        RECT 1084.750 1055.600 1085.070 1055.660 ;
        RECT 1084.555 1055.460 1085.070 1055.600 ;
        RECT 1084.750 1055.400 1085.070 1055.460 ;
        RECT 1082.910 895.120 1083.230 895.180 ;
        RECT 1084.290 895.120 1084.610 895.180 ;
        RECT 1082.910 894.980 1084.610 895.120 ;
        RECT 1082.910 894.920 1083.230 894.980 ;
        RECT 1084.290 894.920 1084.610 894.980 ;
        RECT 1083.830 807.060 1084.150 807.120 ;
        RECT 1083.635 806.920 1084.150 807.060 ;
        RECT 1083.830 806.860 1084.150 806.920 ;
        RECT 1083.845 759.120 1084.135 759.165 ;
        RECT 1084.290 759.120 1084.610 759.180 ;
        RECT 1083.845 758.980 1084.610 759.120 ;
        RECT 1083.845 758.935 1084.135 758.980 ;
        RECT 1084.290 758.920 1084.610 758.980 ;
        RECT 1083.845 676.160 1084.135 676.205 ;
        RECT 1084.290 676.160 1084.610 676.220 ;
        RECT 1083.845 676.020 1084.610 676.160 ;
        RECT 1083.845 675.975 1084.135 676.020 ;
        RECT 1084.290 675.960 1084.610 676.020 ;
        RECT 1083.830 648.620 1084.150 648.680 ;
        RECT 1083.635 648.480 1084.150 648.620 ;
        RECT 1083.830 648.420 1084.150 648.480 ;
        RECT 1083.830 627.880 1084.150 627.940 ;
        RECT 1084.750 627.880 1085.070 627.940 ;
        RECT 1083.830 627.740 1085.070 627.880 ;
        RECT 1083.830 627.680 1084.150 627.740 ;
        RECT 1084.750 627.680 1085.070 627.740 ;
        RECT 1084.750 573.140 1085.070 573.200 ;
        RECT 1084.380 573.000 1085.070 573.140 ;
        RECT 1084.380 572.860 1084.520 573.000 ;
        RECT 1084.750 572.940 1085.070 573.000 ;
        RECT 1084.290 572.600 1084.610 572.860 ;
        RECT 1084.290 475.900 1084.610 475.960 ;
        RECT 1084.095 475.760 1084.610 475.900 ;
        RECT 1084.290 475.700 1084.610 475.760 ;
        RECT 1084.290 427.960 1084.610 428.020 ;
        RECT 1084.095 427.820 1084.610 427.960 ;
        RECT 1084.290 427.760 1084.610 427.820 ;
        RECT 1084.290 352.480 1084.610 352.540 ;
        RECT 1083.920 352.340 1084.610 352.480 ;
        RECT 1083.920 351.860 1084.060 352.340 ;
        RECT 1084.290 352.280 1084.610 352.340 ;
        RECT 1083.830 351.600 1084.150 351.860 ;
        RECT 1084.290 282.780 1084.610 282.840 ;
        RECT 1084.750 282.780 1085.070 282.840 ;
        RECT 1084.290 282.640 1085.070 282.780 ;
        RECT 1084.290 282.580 1084.610 282.640 ;
        RECT 1084.750 282.580 1085.070 282.640 ;
        RECT 1084.750 275.980 1085.070 276.040 ;
        RECT 1084.555 275.840 1085.070 275.980 ;
        RECT 1084.750 275.780 1085.070 275.840 ;
        RECT 1084.750 228.040 1085.070 228.100 ;
        RECT 1084.555 227.900 1085.070 228.040 ;
        RECT 1084.750 227.840 1085.070 227.900 ;
        RECT 1084.290 62.460 1084.610 62.520 ;
        RECT 1083.920 62.320 1084.610 62.460 ;
        RECT 1083.920 62.180 1084.060 62.320 ;
        RECT 1084.290 62.260 1084.610 62.320 ;
        RECT 1083.830 61.920 1084.150 62.180 ;
        RECT 656.950 43.420 657.270 43.480 ;
        RECT 1083.830 43.420 1084.150 43.480 ;
        RECT 656.950 43.280 1084.150 43.420 ;
        RECT 656.950 43.220 657.270 43.280 ;
        RECT 1083.830 43.220 1084.150 43.280 ;
      LAYER via ;
        RECT 1083.860 1104.360 1084.120 1104.620 ;
        RECT 1084.320 1104.360 1084.580 1104.620 ;
        RECT 1083.860 1103.680 1084.120 1103.940 ;
        RECT 1084.780 1103.680 1085.040 1103.940 ;
        RECT 1084.780 1096.880 1085.040 1097.140 ;
        RECT 1084.780 1055.400 1085.040 1055.660 ;
        RECT 1082.940 894.920 1083.200 895.180 ;
        RECT 1084.320 894.920 1084.580 895.180 ;
        RECT 1083.860 806.860 1084.120 807.120 ;
        RECT 1084.320 758.920 1084.580 759.180 ;
        RECT 1084.320 675.960 1084.580 676.220 ;
        RECT 1083.860 648.420 1084.120 648.680 ;
        RECT 1083.860 627.680 1084.120 627.940 ;
        RECT 1084.780 627.680 1085.040 627.940 ;
        RECT 1084.780 572.940 1085.040 573.200 ;
        RECT 1084.320 572.600 1084.580 572.860 ;
        RECT 1084.320 475.700 1084.580 475.960 ;
        RECT 1084.320 427.760 1084.580 428.020 ;
        RECT 1084.320 352.280 1084.580 352.540 ;
        RECT 1083.860 351.600 1084.120 351.860 ;
        RECT 1084.320 282.580 1084.580 282.840 ;
        RECT 1084.780 282.580 1085.040 282.840 ;
        RECT 1084.780 275.780 1085.040 276.040 ;
        RECT 1084.780 227.840 1085.040 228.100 ;
        RECT 1084.320 62.260 1084.580 62.520 ;
        RECT 1083.860 61.920 1084.120 62.180 ;
        RECT 656.980 43.220 657.240 43.480 ;
        RECT 1083.860 43.220 1084.120 43.480 ;
      LAYER met2 ;
        RECT 1087.090 1220.330 1087.650 1228.680 ;
        RECT 1085.760 1220.190 1087.650 1220.330 ;
        RECT 1085.760 1196.700 1085.900 1220.190 ;
        RECT 1087.090 1219.680 1087.650 1220.190 ;
        RECT 1084.380 1196.560 1085.900 1196.700 ;
        RECT 1084.380 1104.650 1084.520 1196.560 ;
        RECT 1083.860 1104.330 1084.120 1104.650 ;
        RECT 1084.320 1104.330 1084.580 1104.650 ;
        RECT 1083.920 1103.970 1084.060 1104.330 ;
        RECT 1083.860 1103.650 1084.120 1103.970 ;
        RECT 1084.780 1103.650 1085.040 1103.970 ;
        RECT 1084.840 1097.170 1084.980 1103.650 ;
        RECT 1084.780 1096.850 1085.040 1097.170 ;
        RECT 1084.780 1055.370 1085.040 1055.690 ;
        RECT 1084.840 1031.290 1084.980 1055.370 ;
        RECT 1084.840 1031.150 1085.900 1031.290 ;
        RECT 1085.760 982.330 1085.900 1031.150 ;
        RECT 1084.380 982.190 1085.900 982.330 ;
        RECT 1084.380 942.210 1084.520 982.190 ;
        RECT 1083.920 942.070 1084.520 942.210 ;
        RECT 1083.920 917.845 1084.060 942.070 ;
        RECT 1082.930 917.475 1083.210 917.845 ;
        RECT 1083.850 917.475 1084.130 917.845 ;
        RECT 1083.000 895.210 1083.140 917.475 ;
        RECT 1082.940 894.890 1083.200 895.210 ;
        RECT 1084.320 894.890 1084.580 895.210 ;
        RECT 1084.380 815.165 1084.520 894.890 ;
        RECT 1084.310 814.795 1084.590 815.165 ;
        RECT 1083.850 814.115 1084.130 814.485 ;
        RECT 1083.920 807.150 1084.060 814.115 ;
        RECT 1083.860 806.830 1084.120 807.150 ;
        RECT 1084.320 758.890 1084.580 759.210 ;
        RECT 1084.380 741.610 1084.520 758.890 ;
        RECT 1084.380 741.470 1084.980 741.610 ;
        RECT 1084.840 689.250 1084.980 741.470 ;
        RECT 1084.380 689.110 1084.980 689.250 ;
        RECT 1084.380 676.250 1084.520 689.110 ;
        RECT 1084.320 675.930 1084.580 676.250 ;
        RECT 1083.860 648.390 1084.120 648.710 ;
        RECT 1083.920 627.970 1084.060 648.390 ;
        RECT 1083.860 627.650 1084.120 627.970 ;
        RECT 1084.780 627.650 1085.040 627.970 ;
        RECT 1084.840 573.230 1084.980 627.650 ;
        RECT 1084.780 572.910 1085.040 573.230 ;
        RECT 1084.320 572.570 1084.580 572.890 ;
        RECT 1084.380 475.990 1084.520 572.570 ;
        RECT 1084.320 475.670 1084.580 475.990 ;
        RECT 1084.320 427.730 1084.580 428.050 ;
        RECT 1084.380 352.570 1084.520 427.730 ;
        RECT 1084.320 352.250 1084.580 352.570 ;
        RECT 1083.860 351.570 1084.120 351.890 ;
        RECT 1083.920 307.090 1084.060 351.570 ;
        RECT 1083.920 306.950 1084.520 307.090 ;
        RECT 1084.380 282.870 1084.520 306.950 ;
        RECT 1084.320 282.550 1084.580 282.870 ;
        RECT 1084.780 282.550 1085.040 282.870 ;
        RECT 1084.840 276.070 1084.980 282.550 ;
        RECT 1084.780 275.750 1085.040 276.070 ;
        RECT 1084.780 227.810 1085.040 228.130 ;
        RECT 1084.840 130.290 1084.980 227.810 ;
        RECT 1084.380 130.150 1084.980 130.290 ;
        RECT 1084.380 62.550 1084.520 130.150 ;
        RECT 1084.320 62.230 1084.580 62.550 ;
        RECT 1083.860 61.890 1084.120 62.210 ;
        RECT 1083.920 43.510 1084.060 61.890 ;
        RECT 656.980 43.190 657.240 43.510 ;
        RECT 1083.860 43.190 1084.120 43.510 ;
        RECT 657.040 2.400 657.180 43.190 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 1082.930 917.520 1083.210 917.800 ;
        RECT 1083.850 917.520 1084.130 917.800 ;
        RECT 1084.310 814.840 1084.590 815.120 ;
        RECT 1083.850 814.160 1084.130 814.440 ;
      LAYER met3 ;
        RECT 1082.905 917.810 1083.235 917.825 ;
        RECT 1083.825 917.810 1084.155 917.825 ;
        RECT 1082.905 917.510 1084.155 917.810 ;
        RECT 1082.905 917.495 1083.235 917.510 ;
        RECT 1083.825 917.495 1084.155 917.510 ;
        RECT 1084.285 815.130 1084.615 815.145 ;
        RECT 1084.070 814.815 1084.615 815.130 ;
        RECT 1084.070 814.465 1084.370 814.815 ;
        RECT 1083.825 814.150 1084.370 814.465 ;
        RECT 1083.825 814.135 1084.155 814.150 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1018.050 1212.680 1018.370 1212.740 ;
        RECT 1261.390 1212.680 1261.710 1212.740 ;
        RECT 1018.050 1212.540 1261.710 1212.680 ;
        RECT 1018.050 1212.480 1018.370 1212.540 ;
        RECT 1261.390 1212.480 1261.710 1212.540 ;
        RECT 995.970 20.640 996.290 20.700 ;
        RECT 1017.590 20.640 1017.910 20.700 ;
        RECT 995.970 20.500 1017.910 20.640 ;
        RECT 995.970 20.440 996.290 20.500 ;
        RECT 1017.590 20.440 1017.910 20.500 ;
      LAYER via ;
        RECT 1018.080 1212.480 1018.340 1212.740 ;
        RECT 1261.420 1212.480 1261.680 1212.740 ;
        RECT 996.000 20.440 996.260 20.700 ;
        RECT 1017.620 20.440 1017.880 20.700 ;
      LAYER met2 ;
        RECT 1261.430 1219.680 1261.990 1228.680 ;
        RECT 1261.480 1212.770 1261.620 1219.680 ;
        RECT 1018.080 1212.450 1018.340 1212.770 ;
        RECT 1261.420 1212.450 1261.680 1212.770 ;
        RECT 1018.140 1193.130 1018.280 1212.450 ;
        RECT 1017.680 1192.990 1018.280 1193.130 ;
        RECT 1017.680 20.730 1017.820 1192.990 ;
        RECT 996.000 20.410 996.260 20.730 ;
        RECT 1017.620 20.410 1017.880 20.730 ;
        RECT 996.060 2.400 996.200 20.410 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1059.450 1214.380 1059.770 1214.440 ;
        RECT 1270.590 1214.380 1270.910 1214.440 ;
        RECT 1059.450 1214.240 1270.910 1214.380 ;
        RECT 1059.450 1214.180 1059.770 1214.240 ;
        RECT 1270.590 1214.180 1270.910 1214.240 ;
        RECT 1013.450 19.960 1013.770 20.020 ;
        RECT 1013.450 19.820 1044.040 19.960 ;
        RECT 1013.450 19.760 1013.770 19.820 ;
        RECT 1043.900 19.620 1044.040 19.820 ;
        RECT 1059.450 19.620 1059.770 19.680 ;
        RECT 1043.900 19.480 1059.770 19.620 ;
        RECT 1059.450 19.420 1059.770 19.480 ;
      LAYER via ;
        RECT 1059.480 1214.180 1059.740 1214.440 ;
        RECT 1270.620 1214.180 1270.880 1214.440 ;
        RECT 1013.480 19.760 1013.740 20.020 ;
        RECT 1059.480 19.420 1059.740 19.680 ;
      LAYER met2 ;
        RECT 1270.630 1219.680 1271.190 1228.680 ;
        RECT 1270.680 1214.470 1270.820 1219.680 ;
        RECT 1059.480 1214.150 1059.740 1214.470 ;
        RECT 1270.620 1214.150 1270.880 1214.470 ;
        RECT 1013.480 19.730 1013.740 20.050 ;
        RECT 1013.540 2.400 1013.680 19.730 ;
        RECT 1059.540 19.710 1059.680 1214.150 ;
        RECT 1059.480 19.390 1059.740 19.710 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1134.890 1208.600 1135.210 1208.660 ;
        RECT 1279.330 1208.600 1279.650 1208.660 ;
        RECT 1134.890 1208.460 1279.650 1208.600 ;
        RECT 1134.890 1208.400 1135.210 1208.460 ;
        RECT 1279.330 1208.400 1279.650 1208.460 ;
        RECT 1031.390 15.200 1031.710 15.260 ;
        RECT 1134.890 15.200 1135.210 15.260 ;
        RECT 1031.390 15.060 1135.210 15.200 ;
        RECT 1031.390 15.000 1031.710 15.060 ;
        RECT 1134.890 15.000 1135.210 15.060 ;
      LAYER via ;
        RECT 1134.920 1208.400 1135.180 1208.660 ;
        RECT 1279.360 1208.400 1279.620 1208.660 ;
        RECT 1031.420 15.000 1031.680 15.260 ;
        RECT 1134.920 15.000 1135.180 15.260 ;
      LAYER met2 ;
        RECT 1279.370 1219.680 1279.930 1228.680 ;
        RECT 1279.420 1208.690 1279.560 1219.680 ;
        RECT 1134.920 1208.370 1135.180 1208.690 ;
        RECT 1279.360 1208.370 1279.620 1208.690 ;
        RECT 1134.980 15.290 1135.120 1208.370 ;
        RECT 1031.420 14.970 1031.680 15.290 ;
        RECT 1134.920 14.970 1135.180 15.290 ;
        RECT 1031.480 2.400 1031.620 14.970 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1221.445 16.065 1221.615 18.275 ;
      LAYER mcon ;
        RECT 1221.445 18.105 1221.615 18.275 ;
      LAYER met1 ;
        RECT 1252.190 1207.580 1252.510 1207.640 ;
        RECT 1288.530 1207.580 1288.850 1207.640 ;
        RECT 1252.190 1207.440 1288.850 1207.580 ;
        RECT 1252.190 1207.380 1252.510 1207.440 ;
        RECT 1288.530 1207.380 1288.850 1207.440 ;
        RECT 1252.190 18.600 1252.510 18.660 ;
        RECT 1222.840 18.460 1252.510 18.600 ;
        RECT 1221.385 18.260 1221.675 18.305 ;
        RECT 1222.840 18.260 1222.980 18.460 ;
        RECT 1252.190 18.400 1252.510 18.460 ;
        RECT 1221.385 18.120 1222.980 18.260 ;
        RECT 1221.385 18.075 1221.675 18.120 ;
        RECT 1049.330 16.220 1049.650 16.280 ;
        RECT 1221.385 16.220 1221.675 16.265 ;
        RECT 1049.330 16.080 1221.675 16.220 ;
        RECT 1049.330 16.020 1049.650 16.080 ;
        RECT 1221.385 16.035 1221.675 16.080 ;
      LAYER via ;
        RECT 1252.220 1207.380 1252.480 1207.640 ;
        RECT 1288.560 1207.380 1288.820 1207.640 ;
        RECT 1252.220 18.400 1252.480 18.660 ;
        RECT 1049.360 16.020 1049.620 16.280 ;
      LAYER met2 ;
        RECT 1288.570 1219.680 1289.130 1228.680 ;
        RECT 1288.620 1207.670 1288.760 1219.680 ;
        RECT 1252.220 1207.350 1252.480 1207.670 ;
        RECT 1288.560 1207.350 1288.820 1207.670 ;
        RECT 1252.280 18.690 1252.420 1207.350 ;
        RECT 1252.220 18.370 1252.480 18.690 ;
        RECT 1049.360 15.990 1049.620 16.310 ;
        RECT 1049.420 2.400 1049.560 15.990 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1297.770 1219.680 1298.330 1228.680 ;
        RECT 1297.820 1210.925 1297.960 1219.680 ;
        RECT 1069.130 1210.555 1069.410 1210.925 ;
        RECT 1297.750 1210.555 1298.030 1210.925 ;
        RECT 1069.200 3.130 1069.340 1210.555 ;
        RECT 1067.360 2.990 1069.340 3.130 ;
        RECT 1067.360 2.400 1067.500 2.990 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
      LAYER via2 ;
        RECT 1069.130 1210.600 1069.410 1210.880 ;
        RECT 1297.750 1210.600 1298.030 1210.880 ;
      LAYER met3 ;
        RECT 1069.105 1210.890 1069.435 1210.905 ;
        RECT 1297.725 1210.890 1298.055 1210.905 ;
        RECT 1069.105 1210.590 1298.055 1210.890 ;
        RECT 1069.105 1210.575 1069.435 1210.590 ;
        RECT 1297.725 1210.575 1298.055 1210.590 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1100.925 15.725 1101.095 16.575 ;
        RECT 1245.365 14.025 1245.535 16.575 ;
      LAYER mcon ;
        RECT 1100.925 16.405 1101.095 16.575 ;
        RECT 1245.365 16.405 1245.535 16.575 ;
      LAYER met1 ;
        RECT 1286.690 1208.600 1287.010 1208.660 ;
        RECT 1306.930 1208.600 1307.250 1208.660 ;
        RECT 1286.690 1208.460 1307.250 1208.600 ;
        RECT 1286.690 1208.400 1287.010 1208.460 ;
        RECT 1306.930 1208.400 1307.250 1208.460 ;
        RECT 1100.865 16.560 1101.155 16.605 ;
        RECT 1245.305 16.560 1245.595 16.605 ;
        RECT 1100.865 16.420 1245.595 16.560 ;
        RECT 1100.865 16.375 1101.155 16.420 ;
        RECT 1245.305 16.375 1245.595 16.420 ;
        RECT 1085.210 15.880 1085.530 15.940 ;
        RECT 1100.865 15.880 1101.155 15.925 ;
        RECT 1085.210 15.740 1101.155 15.880 ;
        RECT 1085.210 15.680 1085.530 15.740 ;
        RECT 1100.865 15.695 1101.155 15.740 ;
        RECT 1245.305 14.180 1245.595 14.225 ;
        RECT 1286.690 14.180 1287.010 14.240 ;
        RECT 1245.305 14.040 1287.010 14.180 ;
        RECT 1245.305 13.995 1245.595 14.040 ;
        RECT 1286.690 13.980 1287.010 14.040 ;
      LAYER via ;
        RECT 1286.720 1208.400 1286.980 1208.660 ;
        RECT 1306.960 1208.400 1307.220 1208.660 ;
        RECT 1085.240 15.680 1085.500 15.940 ;
        RECT 1286.720 13.980 1286.980 14.240 ;
      LAYER met2 ;
        RECT 1306.970 1219.680 1307.530 1228.680 ;
        RECT 1307.020 1208.690 1307.160 1219.680 ;
        RECT 1286.720 1208.370 1286.980 1208.690 ;
        RECT 1306.960 1208.370 1307.220 1208.690 ;
        RECT 1085.240 15.650 1085.500 15.970 ;
        RECT 1085.300 2.400 1085.440 15.650 ;
        RECT 1286.780 14.270 1286.920 1208.370 ;
        RECT 1286.720 13.950 1286.980 14.270 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1307.390 1207.580 1307.710 1207.640 ;
        RECT 1316.130 1207.580 1316.450 1207.640 ;
        RECT 1307.390 1207.440 1316.450 1207.580 ;
        RECT 1307.390 1207.380 1307.710 1207.440 ;
        RECT 1316.130 1207.380 1316.450 1207.440 ;
        RECT 1102.690 20.300 1103.010 20.360 ;
        RECT 1307.390 20.300 1307.710 20.360 ;
        RECT 1102.690 20.160 1307.710 20.300 ;
        RECT 1102.690 20.100 1103.010 20.160 ;
        RECT 1307.390 20.100 1307.710 20.160 ;
      LAYER via ;
        RECT 1307.420 1207.380 1307.680 1207.640 ;
        RECT 1316.160 1207.380 1316.420 1207.640 ;
        RECT 1102.720 20.100 1102.980 20.360 ;
        RECT 1307.420 20.100 1307.680 20.360 ;
      LAYER met2 ;
        RECT 1316.170 1219.680 1316.730 1228.680 ;
        RECT 1316.220 1207.670 1316.360 1219.680 ;
        RECT 1307.420 1207.350 1307.680 1207.670 ;
        RECT 1316.160 1207.350 1316.420 1207.670 ;
        RECT 1307.480 20.390 1307.620 1207.350 ;
        RECT 1102.720 20.070 1102.980 20.390 ;
        RECT 1307.420 20.070 1307.680 20.390 ;
        RECT 1102.780 2.400 1102.920 20.070 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1314.290 1208.600 1314.610 1208.660 ;
        RECT 1325.330 1208.600 1325.650 1208.660 ;
        RECT 1314.290 1208.460 1325.650 1208.600 ;
        RECT 1314.290 1208.400 1314.610 1208.460 ;
        RECT 1325.330 1208.400 1325.650 1208.460 ;
        RECT 1120.630 15.880 1120.950 15.940 ;
        RECT 1314.290 15.880 1314.610 15.940 ;
        RECT 1120.630 15.740 1314.610 15.880 ;
        RECT 1120.630 15.680 1120.950 15.740 ;
        RECT 1314.290 15.680 1314.610 15.740 ;
      LAYER via ;
        RECT 1314.320 1208.400 1314.580 1208.660 ;
        RECT 1325.360 1208.400 1325.620 1208.660 ;
        RECT 1120.660 15.680 1120.920 15.940 ;
        RECT 1314.320 15.680 1314.580 15.940 ;
      LAYER met2 ;
        RECT 1325.370 1219.680 1325.930 1228.680 ;
        RECT 1325.420 1208.690 1325.560 1219.680 ;
        RECT 1314.320 1208.370 1314.580 1208.690 ;
        RECT 1325.360 1208.370 1325.620 1208.690 ;
        RECT 1314.380 15.970 1314.520 1208.370 ;
        RECT 1120.660 15.650 1120.920 15.970 ;
        RECT 1314.320 15.650 1314.580 15.970 ;
        RECT 1120.720 2.400 1120.860 15.650 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1160.725 14.365 1160.895 15.555 ;
      LAYER mcon ;
        RECT 1160.725 15.385 1160.895 15.555 ;
      LAYER met1 ;
        RECT 1160.665 15.540 1160.955 15.585 ;
        RECT 1332.230 15.540 1332.550 15.600 ;
        RECT 1160.665 15.400 1332.550 15.540 ;
        RECT 1160.665 15.355 1160.955 15.400 ;
        RECT 1332.230 15.340 1332.550 15.400 ;
        RECT 1138.570 14.520 1138.890 14.580 ;
        RECT 1160.665 14.520 1160.955 14.565 ;
        RECT 1138.570 14.380 1160.955 14.520 ;
        RECT 1138.570 14.320 1138.890 14.380 ;
        RECT 1160.665 14.335 1160.955 14.380 ;
      LAYER via ;
        RECT 1332.260 15.340 1332.520 15.600 ;
        RECT 1138.600 14.320 1138.860 14.580 ;
      LAYER met2 ;
        RECT 1334.570 1220.330 1335.130 1228.680 ;
        RECT 1332.320 1220.190 1335.130 1220.330 ;
        RECT 1332.320 15.630 1332.460 1220.190 ;
        RECT 1334.570 1219.680 1335.130 1220.190 ;
        RECT 1332.260 15.310 1332.520 15.630 ;
        RECT 1138.600 14.290 1138.860 14.610 ;
        RECT 1138.660 2.400 1138.800 14.290 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 1209.960 1159.130 1210.020 ;
        RECT 1343.730 1209.960 1344.050 1210.020 ;
        RECT 1158.810 1209.820 1344.050 1209.960 ;
        RECT 1158.810 1209.760 1159.130 1209.820 ;
        RECT 1343.730 1209.760 1344.050 1209.820 ;
        RECT 1156.510 18.260 1156.830 18.320 ;
        RECT 1158.810 18.260 1159.130 18.320 ;
        RECT 1156.510 18.120 1159.130 18.260 ;
        RECT 1156.510 18.060 1156.830 18.120 ;
        RECT 1158.810 18.060 1159.130 18.120 ;
      LAYER via ;
        RECT 1158.840 1209.760 1159.100 1210.020 ;
        RECT 1343.760 1209.760 1344.020 1210.020 ;
        RECT 1156.540 18.060 1156.800 18.320 ;
        RECT 1158.840 18.060 1159.100 18.320 ;
      LAYER met2 ;
        RECT 1343.770 1219.680 1344.330 1228.680 ;
        RECT 1343.820 1210.050 1343.960 1219.680 ;
        RECT 1158.840 1209.730 1159.100 1210.050 ;
        RECT 1343.760 1209.730 1344.020 1210.050 ;
        RECT 1158.900 18.350 1159.040 1209.730 ;
        RECT 1156.540 18.030 1156.800 18.350 ;
        RECT 1158.840 18.030 1159.100 18.350 ;
        RECT 1156.600 2.400 1156.740 18.030 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1091.265 1027.905 1091.435 1097.095 ;
        RECT 1091.265 965.685 1091.435 1007.335 ;
        RECT 1091.265 900.065 1091.435 917.235 ;
        RECT 1091.725 427.805 1091.895 475.915 ;
        RECT 1091.265 234.685 1091.435 324.275 ;
      LAYER mcon ;
        RECT 1091.265 1096.925 1091.435 1097.095 ;
        RECT 1091.265 1007.165 1091.435 1007.335 ;
        RECT 1091.265 917.065 1091.435 917.235 ;
        RECT 1091.725 475.745 1091.895 475.915 ;
        RECT 1091.265 324.105 1091.435 324.275 ;
      LAYER met1 ;
        RECT 1092.110 1124.960 1092.430 1125.020 ;
        RECT 1091.280 1124.820 1092.430 1124.960 ;
        RECT 1091.280 1124.680 1091.420 1124.820 ;
        RECT 1092.110 1124.760 1092.430 1124.820 ;
        RECT 1091.190 1124.420 1091.510 1124.680 ;
        RECT 1091.190 1103.880 1091.510 1103.940 ;
        RECT 1091.650 1103.880 1091.970 1103.940 ;
        RECT 1091.190 1103.740 1091.970 1103.880 ;
        RECT 1091.190 1103.680 1091.510 1103.740 ;
        RECT 1091.650 1103.680 1091.970 1103.740 ;
        RECT 1091.205 1097.080 1091.495 1097.125 ;
        RECT 1091.650 1097.080 1091.970 1097.140 ;
        RECT 1091.205 1096.940 1091.970 1097.080 ;
        RECT 1091.205 1096.895 1091.495 1096.940 ;
        RECT 1091.650 1096.880 1091.970 1096.940 ;
        RECT 1091.190 1028.060 1091.510 1028.120 ;
        RECT 1090.995 1027.920 1091.510 1028.060 ;
        RECT 1091.190 1027.860 1091.510 1027.920 ;
        RECT 1091.190 1007.320 1091.510 1007.380 ;
        RECT 1090.995 1007.180 1091.510 1007.320 ;
        RECT 1091.190 1007.120 1091.510 1007.180 ;
        RECT 1091.205 965.840 1091.495 965.885 ;
        RECT 1091.650 965.840 1091.970 965.900 ;
        RECT 1091.205 965.700 1091.970 965.840 ;
        RECT 1091.205 965.655 1091.495 965.700 ;
        RECT 1091.650 965.640 1091.970 965.700 ;
        RECT 1091.190 917.900 1091.510 917.960 ;
        RECT 1092.110 917.900 1092.430 917.960 ;
        RECT 1091.190 917.760 1092.430 917.900 ;
        RECT 1091.190 917.700 1091.510 917.760 ;
        RECT 1092.110 917.700 1092.430 917.760 ;
        RECT 1091.190 917.220 1091.510 917.280 ;
        RECT 1090.995 917.080 1091.510 917.220 ;
        RECT 1091.190 917.020 1091.510 917.080 ;
        RECT 1091.205 900.220 1091.495 900.265 ;
        RECT 1091.650 900.220 1091.970 900.280 ;
        RECT 1091.205 900.080 1091.970 900.220 ;
        RECT 1091.205 900.035 1091.495 900.080 ;
        RECT 1091.650 900.020 1091.970 900.080 ;
        RECT 1089.810 807.060 1090.130 807.120 ;
        RECT 1091.190 807.060 1091.510 807.120 ;
        RECT 1089.810 806.920 1091.510 807.060 ;
        RECT 1089.810 806.860 1090.130 806.920 ;
        RECT 1091.190 806.860 1091.510 806.920 ;
        RECT 1089.810 710.840 1090.130 710.900 ;
        RECT 1092.110 710.840 1092.430 710.900 ;
        RECT 1089.810 710.700 1092.430 710.840 ;
        RECT 1089.810 710.640 1090.130 710.700 ;
        RECT 1092.110 710.640 1092.430 710.700 ;
        RECT 1091.650 642.160 1091.970 642.220 ;
        RECT 1091.280 642.020 1091.970 642.160 ;
        RECT 1091.280 641.540 1091.420 642.020 ;
        RECT 1091.650 641.960 1091.970 642.020 ;
        RECT 1091.190 641.280 1091.510 641.540 ;
        RECT 1091.190 627.880 1091.510 627.940 ;
        RECT 1092.110 627.880 1092.430 627.940 ;
        RECT 1091.190 627.740 1092.430 627.880 ;
        RECT 1091.190 627.680 1091.510 627.740 ;
        RECT 1092.110 627.680 1092.430 627.740 ;
        RECT 1091.650 545.400 1091.970 545.660 ;
        RECT 1091.740 544.980 1091.880 545.400 ;
        RECT 1091.650 544.720 1091.970 544.980 ;
        RECT 1091.650 475.900 1091.970 475.960 ;
        RECT 1091.455 475.760 1091.970 475.900 ;
        RECT 1091.650 475.700 1091.970 475.760 ;
        RECT 1091.650 427.960 1091.970 428.020 ;
        RECT 1091.455 427.820 1091.970 427.960 ;
        RECT 1091.650 427.760 1091.970 427.820 ;
        RECT 1091.190 324.260 1091.510 324.320 ;
        RECT 1090.995 324.120 1091.510 324.260 ;
        RECT 1091.190 324.060 1091.510 324.120 ;
        RECT 1091.190 234.840 1091.510 234.900 ;
        RECT 1090.995 234.700 1091.510 234.840 ;
        RECT 1091.190 234.640 1091.510 234.700 ;
        RECT 1091.190 227.700 1091.510 227.760 ;
        RECT 1091.650 227.700 1091.970 227.760 ;
        RECT 1091.190 227.560 1091.970 227.700 ;
        RECT 1091.190 227.500 1091.510 227.560 ;
        RECT 1091.650 227.500 1091.970 227.560 ;
        RECT 1091.190 96.940 1091.510 97.200 ;
        RECT 1091.280 96.520 1091.420 96.940 ;
        RECT 1091.190 96.260 1091.510 96.520 ;
        RECT 674.430 43.080 674.750 43.140 ;
        RECT 1091.190 43.080 1091.510 43.140 ;
        RECT 674.430 42.940 1091.510 43.080 ;
        RECT 674.430 42.880 674.750 42.940 ;
        RECT 1091.190 42.880 1091.510 42.940 ;
      LAYER via ;
        RECT 1092.140 1124.760 1092.400 1125.020 ;
        RECT 1091.220 1124.420 1091.480 1124.680 ;
        RECT 1091.220 1103.680 1091.480 1103.940 ;
        RECT 1091.680 1103.680 1091.940 1103.940 ;
        RECT 1091.680 1096.880 1091.940 1097.140 ;
        RECT 1091.220 1027.860 1091.480 1028.120 ;
        RECT 1091.220 1007.120 1091.480 1007.380 ;
        RECT 1091.680 965.640 1091.940 965.900 ;
        RECT 1091.220 917.700 1091.480 917.960 ;
        RECT 1092.140 917.700 1092.400 917.960 ;
        RECT 1091.220 917.020 1091.480 917.280 ;
        RECT 1091.680 900.020 1091.940 900.280 ;
        RECT 1089.840 806.860 1090.100 807.120 ;
        RECT 1091.220 806.860 1091.480 807.120 ;
        RECT 1089.840 710.640 1090.100 710.900 ;
        RECT 1092.140 710.640 1092.400 710.900 ;
        RECT 1091.680 641.960 1091.940 642.220 ;
        RECT 1091.220 641.280 1091.480 641.540 ;
        RECT 1091.220 627.680 1091.480 627.940 ;
        RECT 1092.140 627.680 1092.400 627.940 ;
        RECT 1091.680 545.400 1091.940 545.660 ;
        RECT 1091.680 544.720 1091.940 544.980 ;
        RECT 1091.680 475.700 1091.940 475.960 ;
        RECT 1091.680 427.760 1091.940 428.020 ;
        RECT 1091.220 324.060 1091.480 324.320 ;
        RECT 1091.220 234.640 1091.480 234.900 ;
        RECT 1091.220 227.500 1091.480 227.760 ;
        RECT 1091.680 227.500 1091.940 227.760 ;
        RECT 1091.220 96.940 1091.480 97.200 ;
        RECT 1091.220 96.260 1091.480 96.520 ;
        RECT 674.460 42.880 674.720 43.140 ;
        RECT 1091.220 42.880 1091.480 43.140 ;
      LAYER met2 ;
        RECT 1096.290 1220.330 1096.850 1228.680 ;
        RECT 1094.960 1220.190 1096.850 1220.330 ;
        RECT 1094.960 1145.645 1095.100 1220.190 ;
        RECT 1096.290 1219.680 1096.850 1220.190 ;
        RECT 1092.130 1145.275 1092.410 1145.645 ;
        RECT 1094.890 1145.275 1095.170 1145.645 ;
        RECT 1092.200 1125.050 1092.340 1145.275 ;
        RECT 1092.140 1124.730 1092.400 1125.050 ;
        RECT 1091.220 1124.390 1091.480 1124.710 ;
        RECT 1091.280 1103.970 1091.420 1124.390 ;
        RECT 1091.220 1103.650 1091.480 1103.970 ;
        RECT 1091.680 1103.650 1091.940 1103.970 ;
        RECT 1091.740 1097.170 1091.880 1103.650 ;
        RECT 1091.680 1096.850 1091.940 1097.170 ;
        RECT 1091.220 1027.830 1091.480 1028.150 ;
        RECT 1091.280 1007.410 1091.420 1027.830 ;
        RECT 1091.220 1007.090 1091.480 1007.410 ;
        RECT 1091.680 965.610 1091.940 965.930 ;
        RECT 1091.740 959.210 1091.880 965.610 ;
        RECT 1091.740 959.070 1092.340 959.210 ;
        RECT 1092.200 917.990 1092.340 959.070 ;
        RECT 1091.220 917.670 1091.480 917.990 ;
        RECT 1092.140 917.670 1092.400 917.990 ;
        RECT 1091.280 917.310 1091.420 917.670 ;
        RECT 1091.220 916.990 1091.480 917.310 ;
        RECT 1091.680 899.990 1091.940 900.310 ;
        RECT 1091.740 815.165 1091.880 899.990 ;
        RECT 1091.670 814.795 1091.950 815.165 ;
        RECT 1091.210 814.115 1091.490 814.485 ;
        RECT 1091.280 807.150 1091.420 814.115 ;
        RECT 1089.840 806.830 1090.100 807.150 ;
        RECT 1091.220 806.830 1091.480 807.150 ;
        RECT 1089.900 759.405 1090.040 806.830 ;
        RECT 1089.830 759.035 1090.110 759.405 ;
        RECT 1089.830 758.355 1090.110 758.725 ;
        RECT 1089.900 710.930 1090.040 758.355 ;
        RECT 1089.840 710.610 1090.100 710.930 ;
        RECT 1092.140 710.610 1092.400 710.930 ;
        RECT 1092.200 689.250 1092.340 710.610 ;
        RECT 1091.740 689.110 1092.340 689.250 ;
        RECT 1091.740 642.250 1091.880 689.110 ;
        RECT 1091.680 641.930 1091.940 642.250 ;
        RECT 1091.220 641.250 1091.480 641.570 ;
        RECT 1091.280 627.970 1091.420 641.250 ;
        RECT 1091.220 627.650 1091.480 627.970 ;
        RECT 1092.140 627.650 1092.400 627.970 ;
        RECT 1092.200 596.770 1092.340 627.650 ;
        RECT 1091.740 596.630 1092.340 596.770 ;
        RECT 1091.740 545.690 1091.880 596.630 ;
        RECT 1091.680 545.370 1091.940 545.690 ;
        RECT 1091.680 544.690 1091.940 545.010 ;
        RECT 1091.740 475.990 1091.880 544.690 ;
        RECT 1091.680 475.670 1091.940 475.990 ;
        RECT 1091.680 427.730 1091.940 428.050 ;
        RECT 1091.740 355.370 1091.880 427.730 ;
        RECT 1091.280 355.230 1091.880 355.370 ;
        RECT 1091.280 324.350 1091.420 355.230 ;
        RECT 1091.220 324.030 1091.480 324.350 ;
        RECT 1091.220 234.610 1091.480 234.930 ;
        RECT 1091.280 227.790 1091.420 234.610 ;
        RECT 1091.220 227.470 1091.480 227.790 ;
        RECT 1091.680 227.470 1091.940 227.790 ;
        RECT 1091.740 186.050 1091.880 227.470 ;
        RECT 1091.280 185.910 1091.880 186.050 ;
        RECT 1091.280 97.230 1091.420 185.910 ;
        RECT 1091.220 96.910 1091.480 97.230 ;
        RECT 1091.220 96.230 1091.480 96.550 ;
        RECT 1091.280 43.170 1091.420 96.230 ;
        RECT 674.460 42.850 674.720 43.170 ;
        RECT 1091.220 42.850 1091.480 43.170 ;
        RECT 674.520 2.400 674.660 42.850 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1092.130 1145.320 1092.410 1145.600 ;
        RECT 1094.890 1145.320 1095.170 1145.600 ;
        RECT 1091.670 814.840 1091.950 815.120 ;
        RECT 1091.210 814.160 1091.490 814.440 ;
        RECT 1089.830 759.080 1090.110 759.360 ;
        RECT 1089.830 758.400 1090.110 758.680 ;
      LAYER met3 ;
        RECT 1092.105 1145.610 1092.435 1145.625 ;
        RECT 1094.865 1145.610 1095.195 1145.625 ;
        RECT 1092.105 1145.310 1095.195 1145.610 ;
        RECT 1092.105 1145.295 1092.435 1145.310 ;
        RECT 1094.865 1145.295 1095.195 1145.310 ;
        RECT 1091.645 815.130 1091.975 815.145 ;
        RECT 1091.430 814.815 1091.975 815.130 ;
        RECT 1091.430 814.465 1091.730 814.815 ;
        RECT 1091.185 814.150 1091.730 814.465 ;
        RECT 1091.185 814.135 1091.515 814.150 ;
        RECT 1089.805 759.370 1090.135 759.385 ;
        RECT 1089.805 759.070 1090.810 759.370 ;
        RECT 1089.805 759.055 1090.135 759.070 ;
        RECT 1089.805 758.690 1090.135 758.705 ;
        RECT 1090.510 758.690 1090.810 759.070 ;
        RECT 1089.805 758.390 1090.810 758.690 ;
        RECT 1089.805 758.375 1090.135 758.390 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 17.240 1174.310 17.300 ;
        RECT 1342.350 17.240 1342.670 17.300 ;
        RECT 1173.990 17.100 1342.670 17.240 ;
        RECT 1173.990 17.040 1174.310 17.100 ;
        RECT 1342.350 17.040 1342.670 17.100 ;
      LAYER via ;
        RECT 1174.020 17.040 1174.280 17.300 ;
        RECT 1342.380 17.040 1342.640 17.300 ;
      LAYER met2 ;
        RECT 1352.970 1219.680 1353.530 1228.680 ;
        RECT 1353.020 1208.205 1353.160 1219.680 ;
        RECT 1342.370 1207.835 1342.650 1208.205 ;
        RECT 1352.950 1207.835 1353.230 1208.205 ;
        RECT 1342.440 17.330 1342.580 1207.835 ;
        RECT 1174.020 17.010 1174.280 17.330 ;
        RECT 1342.380 17.010 1342.640 17.330 ;
        RECT 1174.080 2.400 1174.220 17.010 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
      LAYER via2 ;
        RECT 1342.370 1207.880 1342.650 1208.160 ;
        RECT 1352.950 1207.880 1353.230 1208.160 ;
      LAYER met3 ;
        RECT 1342.345 1208.170 1342.675 1208.185 ;
        RECT 1352.925 1208.170 1353.255 1208.185 ;
        RECT 1342.345 1207.870 1353.255 1208.170 ;
        RECT 1342.345 1207.855 1342.675 1207.870 ;
        RECT 1352.925 1207.855 1353.255 1207.870 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1193.385 1207.425 1193.555 1208.955 ;
        RECT 1192.465 862.665 1192.635 910.775 ;
        RECT 1193.385 628.065 1193.555 717.655 ;
        RECT 1192.925 572.645 1193.095 620.755 ;
        RECT 1193.385 476.085 1193.555 524.195 ;
        RECT 1193.385 379.525 1193.555 427.635 ;
        RECT 1193.385 241.485 1193.555 331.075 ;
        RECT 1192.925 186.405 1193.095 234.515 ;
        RECT 1193.385 138.465 1193.555 145.095 ;
        RECT 1192.925 48.365 1193.095 137.955 ;
      LAYER mcon ;
        RECT 1193.385 1208.785 1193.555 1208.955 ;
        RECT 1192.465 910.605 1192.635 910.775 ;
        RECT 1193.385 717.485 1193.555 717.655 ;
        RECT 1192.925 620.585 1193.095 620.755 ;
        RECT 1193.385 524.025 1193.555 524.195 ;
        RECT 1193.385 427.465 1193.555 427.635 ;
        RECT 1193.385 330.905 1193.555 331.075 ;
        RECT 1192.925 234.345 1193.095 234.515 ;
        RECT 1193.385 144.925 1193.555 145.095 ;
        RECT 1192.925 137.785 1193.095 137.955 ;
      LAYER met1 ;
        RECT 1193.325 1208.940 1193.615 1208.985 ;
        RECT 1362.130 1208.940 1362.450 1209.000 ;
        RECT 1193.325 1208.800 1362.450 1208.940 ;
        RECT 1193.325 1208.755 1193.615 1208.800 ;
        RECT 1362.130 1208.740 1362.450 1208.800 ;
        RECT 1193.310 1207.580 1193.630 1207.640 ;
        RECT 1193.115 1207.440 1193.630 1207.580 ;
        RECT 1193.310 1207.380 1193.630 1207.440 ;
        RECT 1192.390 1152.500 1192.710 1152.560 ;
        RECT 1193.310 1152.500 1193.630 1152.560 ;
        RECT 1192.390 1152.360 1193.630 1152.500 ;
        RECT 1192.390 1152.300 1192.710 1152.360 ;
        RECT 1193.310 1152.300 1193.630 1152.360 ;
        RECT 1192.390 1031.460 1192.710 1031.520 ;
        RECT 1193.310 1031.460 1193.630 1031.520 ;
        RECT 1192.390 1031.320 1193.630 1031.460 ;
        RECT 1192.390 1031.260 1192.710 1031.320 ;
        RECT 1193.310 1031.260 1193.630 1031.320 ;
        RECT 1192.390 1007.320 1192.710 1007.380 ;
        RECT 1193.310 1007.320 1193.630 1007.380 ;
        RECT 1192.390 1007.180 1193.630 1007.320 ;
        RECT 1192.390 1007.120 1192.710 1007.180 ;
        RECT 1193.310 1007.120 1193.630 1007.180 ;
        RECT 1192.390 917.900 1192.710 917.960 ;
        RECT 1193.310 917.900 1193.630 917.960 ;
        RECT 1192.390 917.760 1193.630 917.900 ;
        RECT 1192.390 917.700 1192.710 917.760 ;
        RECT 1193.310 917.700 1193.630 917.760 ;
        RECT 1192.405 910.760 1192.695 910.805 ;
        RECT 1193.310 910.760 1193.630 910.820 ;
        RECT 1192.405 910.620 1193.630 910.760 ;
        RECT 1192.405 910.575 1192.695 910.620 ;
        RECT 1193.310 910.560 1193.630 910.620 ;
        RECT 1192.390 862.820 1192.710 862.880 ;
        RECT 1192.195 862.680 1192.710 862.820 ;
        RECT 1192.390 862.620 1192.710 862.680 ;
        RECT 1192.390 821.340 1192.710 821.400 ;
        RECT 1193.310 821.340 1193.630 821.400 ;
        RECT 1192.390 821.200 1193.630 821.340 ;
        RECT 1192.390 821.140 1192.710 821.200 ;
        RECT 1193.310 821.140 1193.630 821.200 ;
        RECT 1191.930 814.200 1192.250 814.260 ;
        RECT 1193.310 814.200 1193.630 814.260 ;
        RECT 1191.930 814.060 1193.630 814.200 ;
        RECT 1191.930 814.000 1192.250 814.060 ;
        RECT 1193.310 814.000 1193.630 814.060 ;
        RECT 1192.850 724.780 1193.170 724.840 ;
        RECT 1193.310 724.780 1193.630 724.840 ;
        RECT 1192.850 724.640 1193.630 724.780 ;
        RECT 1192.850 724.580 1193.170 724.640 ;
        RECT 1193.310 724.580 1193.630 724.640 ;
        RECT 1193.310 717.640 1193.630 717.700 ;
        RECT 1193.115 717.500 1193.630 717.640 ;
        RECT 1193.310 717.440 1193.630 717.500 ;
        RECT 1193.310 628.220 1193.630 628.280 ;
        RECT 1193.115 628.080 1193.630 628.220 ;
        RECT 1193.310 628.020 1193.630 628.080 ;
        RECT 1192.865 620.740 1193.155 620.785 ;
        RECT 1193.310 620.740 1193.630 620.800 ;
        RECT 1192.865 620.600 1193.630 620.740 ;
        RECT 1192.865 620.555 1193.155 620.600 ;
        RECT 1193.310 620.540 1193.630 620.600 ;
        RECT 1192.850 572.800 1193.170 572.860 ;
        RECT 1192.655 572.660 1193.170 572.800 ;
        RECT 1192.850 572.600 1193.170 572.660 ;
        RECT 1192.850 531.660 1193.170 531.720 ;
        RECT 1193.310 531.660 1193.630 531.720 ;
        RECT 1192.850 531.520 1193.630 531.660 ;
        RECT 1192.850 531.460 1193.170 531.520 ;
        RECT 1193.310 531.460 1193.630 531.520 ;
        RECT 1193.310 524.180 1193.630 524.240 ;
        RECT 1193.115 524.040 1193.630 524.180 ;
        RECT 1193.310 523.980 1193.630 524.040 ;
        RECT 1193.310 476.240 1193.630 476.300 ;
        RECT 1193.115 476.100 1193.630 476.240 ;
        RECT 1193.310 476.040 1193.630 476.100 ;
        RECT 1193.310 427.620 1193.630 427.680 ;
        RECT 1193.115 427.480 1193.630 427.620 ;
        RECT 1193.310 427.420 1193.630 427.480 ;
        RECT 1193.310 379.680 1193.630 379.740 ;
        RECT 1193.115 379.540 1193.630 379.680 ;
        RECT 1193.310 379.480 1193.630 379.540 ;
        RECT 1193.310 331.060 1193.630 331.120 ;
        RECT 1193.115 330.920 1193.630 331.060 ;
        RECT 1193.310 330.860 1193.630 330.920 ;
        RECT 1193.310 241.640 1193.630 241.700 ;
        RECT 1193.115 241.500 1193.630 241.640 ;
        RECT 1193.310 241.440 1193.630 241.500 ;
        RECT 1192.865 234.500 1193.155 234.545 ;
        RECT 1193.310 234.500 1193.630 234.560 ;
        RECT 1192.865 234.360 1193.630 234.500 ;
        RECT 1192.865 234.315 1193.155 234.360 ;
        RECT 1193.310 234.300 1193.630 234.360 ;
        RECT 1192.865 186.560 1193.155 186.605 ;
        RECT 1193.310 186.560 1193.630 186.620 ;
        RECT 1192.865 186.420 1193.630 186.560 ;
        RECT 1192.865 186.375 1193.155 186.420 ;
        RECT 1193.310 186.360 1193.630 186.420 ;
        RECT 1193.310 145.080 1193.630 145.140 ;
        RECT 1193.115 144.940 1193.630 145.080 ;
        RECT 1193.310 144.880 1193.630 144.940 ;
        RECT 1193.310 138.620 1193.630 138.680 ;
        RECT 1193.115 138.480 1193.630 138.620 ;
        RECT 1193.310 138.420 1193.630 138.480 ;
        RECT 1192.865 137.940 1193.155 137.985 ;
        RECT 1193.310 137.940 1193.630 138.000 ;
        RECT 1192.865 137.800 1193.630 137.940 ;
        RECT 1192.865 137.755 1193.155 137.800 ;
        RECT 1193.310 137.740 1193.630 137.800 ;
        RECT 1192.850 48.520 1193.170 48.580 ;
        RECT 1192.655 48.380 1193.170 48.520 ;
        RECT 1192.850 48.320 1193.170 48.380 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1192.850 2.960 1193.170 3.020 ;
        RECT 1191.930 2.820 1193.170 2.960 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
        RECT 1192.850 2.760 1193.170 2.820 ;
      LAYER via ;
        RECT 1362.160 1208.740 1362.420 1209.000 ;
        RECT 1193.340 1207.380 1193.600 1207.640 ;
        RECT 1192.420 1152.300 1192.680 1152.560 ;
        RECT 1193.340 1152.300 1193.600 1152.560 ;
        RECT 1192.420 1031.260 1192.680 1031.520 ;
        RECT 1193.340 1031.260 1193.600 1031.520 ;
        RECT 1192.420 1007.120 1192.680 1007.380 ;
        RECT 1193.340 1007.120 1193.600 1007.380 ;
        RECT 1192.420 917.700 1192.680 917.960 ;
        RECT 1193.340 917.700 1193.600 917.960 ;
        RECT 1193.340 910.560 1193.600 910.820 ;
        RECT 1192.420 862.620 1192.680 862.880 ;
        RECT 1192.420 821.140 1192.680 821.400 ;
        RECT 1193.340 821.140 1193.600 821.400 ;
        RECT 1191.960 814.000 1192.220 814.260 ;
        RECT 1193.340 814.000 1193.600 814.260 ;
        RECT 1192.880 724.580 1193.140 724.840 ;
        RECT 1193.340 724.580 1193.600 724.840 ;
        RECT 1193.340 717.440 1193.600 717.700 ;
        RECT 1193.340 628.020 1193.600 628.280 ;
        RECT 1193.340 620.540 1193.600 620.800 ;
        RECT 1192.880 572.600 1193.140 572.860 ;
        RECT 1192.880 531.460 1193.140 531.720 ;
        RECT 1193.340 531.460 1193.600 531.720 ;
        RECT 1193.340 523.980 1193.600 524.240 ;
        RECT 1193.340 476.040 1193.600 476.300 ;
        RECT 1193.340 427.420 1193.600 427.680 ;
        RECT 1193.340 379.480 1193.600 379.740 ;
        RECT 1193.340 330.860 1193.600 331.120 ;
        RECT 1193.340 241.440 1193.600 241.700 ;
        RECT 1193.340 234.300 1193.600 234.560 ;
        RECT 1193.340 186.360 1193.600 186.620 ;
        RECT 1193.340 144.880 1193.600 145.140 ;
        RECT 1193.340 138.420 1193.600 138.680 ;
        RECT 1193.340 137.740 1193.600 138.000 ;
        RECT 1192.880 48.320 1193.140 48.580 ;
        RECT 1191.960 2.760 1192.220 3.020 ;
        RECT 1192.880 2.760 1193.140 3.020 ;
      LAYER met2 ;
        RECT 1362.170 1219.680 1362.730 1228.680 ;
        RECT 1362.220 1209.030 1362.360 1219.680 ;
        RECT 1362.160 1208.710 1362.420 1209.030 ;
        RECT 1193.340 1207.350 1193.600 1207.670 ;
        RECT 1193.400 1200.725 1193.540 1207.350 ;
        RECT 1192.410 1200.355 1192.690 1200.725 ;
        RECT 1193.330 1200.355 1193.610 1200.725 ;
        RECT 1192.480 1152.590 1192.620 1200.355 ;
        RECT 1192.420 1152.270 1192.680 1152.590 ;
        RECT 1193.340 1152.270 1193.600 1152.590 ;
        RECT 1193.400 1104.165 1193.540 1152.270 ;
        RECT 1192.410 1103.795 1192.690 1104.165 ;
        RECT 1193.330 1103.795 1193.610 1104.165 ;
        RECT 1192.480 1055.885 1192.620 1103.795 ;
        RECT 1192.410 1055.515 1192.690 1055.885 ;
        RECT 1193.330 1055.515 1193.610 1055.885 ;
        RECT 1193.400 1031.550 1193.540 1055.515 ;
        RECT 1192.420 1031.230 1192.680 1031.550 ;
        RECT 1193.340 1031.230 1193.600 1031.550 ;
        RECT 1192.480 1007.605 1192.620 1031.230 ;
        RECT 1192.410 1007.235 1192.690 1007.605 ;
        RECT 1193.330 1007.235 1193.610 1007.605 ;
        RECT 1192.420 1007.090 1192.680 1007.235 ;
        RECT 1193.340 1007.090 1193.600 1007.235 ;
        RECT 1192.480 917.990 1192.620 1007.090 ;
        RECT 1192.420 917.670 1192.680 917.990 ;
        RECT 1193.340 917.670 1193.600 917.990 ;
        RECT 1193.400 910.850 1193.540 917.670 ;
        RECT 1193.340 910.530 1193.600 910.850 ;
        RECT 1192.420 862.590 1192.680 862.910 ;
        RECT 1192.480 821.430 1192.620 862.590 ;
        RECT 1192.420 821.110 1192.680 821.430 ;
        RECT 1193.340 821.110 1193.600 821.430 ;
        RECT 1193.400 814.290 1193.540 821.110 ;
        RECT 1191.960 813.970 1192.220 814.290 ;
        RECT 1193.340 813.970 1193.600 814.290 ;
        RECT 1192.020 766.205 1192.160 813.970 ;
        RECT 1191.950 765.835 1192.230 766.205 ;
        RECT 1192.870 765.835 1193.150 766.205 ;
        RECT 1192.940 724.870 1193.080 765.835 ;
        RECT 1192.880 724.550 1193.140 724.870 ;
        RECT 1193.340 724.550 1193.600 724.870 ;
        RECT 1193.400 717.730 1193.540 724.550 ;
        RECT 1193.340 717.410 1193.600 717.730 ;
        RECT 1193.340 627.990 1193.600 628.310 ;
        RECT 1193.400 620.830 1193.540 627.990 ;
        RECT 1193.340 620.510 1193.600 620.830 ;
        RECT 1192.880 572.570 1193.140 572.890 ;
        RECT 1192.940 531.750 1193.080 572.570 ;
        RECT 1192.880 531.430 1193.140 531.750 ;
        RECT 1193.340 531.430 1193.600 531.750 ;
        RECT 1193.400 524.270 1193.540 531.430 ;
        RECT 1193.340 523.950 1193.600 524.270 ;
        RECT 1193.340 476.010 1193.600 476.330 ;
        RECT 1193.400 427.710 1193.540 476.010 ;
        RECT 1193.340 427.390 1193.600 427.710 ;
        RECT 1193.340 379.450 1193.600 379.770 ;
        RECT 1193.400 331.150 1193.540 379.450 ;
        RECT 1193.340 330.830 1193.600 331.150 ;
        RECT 1193.340 241.410 1193.600 241.730 ;
        RECT 1193.400 234.590 1193.540 241.410 ;
        RECT 1193.340 234.270 1193.600 234.590 ;
        RECT 1193.340 186.330 1193.600 186.650 ;
        RECT 1193.400 145.170 1193.540 186.330 ;
        RECT 1193.340 144.850 1193.600 145.170 ;
        RECT 1193.340 138.390 1193.600 138.710 ;
        RECT 1193.400 138.030 1193.540 138.390 ;
        RECT 1193.340 137.710 1193.600 138.030 ;
        RECT 1192.880 48.290 1193.140 48.610 ;
        RECT 1192.940 3.050 1193.080 48.290 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1192.880 2.730 1193.140 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 1192.410 1200.400 1192.690 1200.680 ;
        RECT 1193.330 1200.400 1193.610 1200.680 ;
        RECT 1192.410 1103.840 1192.690 1104.120 ;
        RECT 1193.330 1103.840 1193.610 1104.120 ;
        RECT 1192.410 1055.560 1192.690 1055.840 ;
        RECT 1193.330 1055.560 1193.610 1055.840 ;
        RECT 1192.410 1007.280 1192.690 1007.560 ;
        RECT 1193.330 1007.280 1193.610 1007.560 ;
        RECT 1191.950 765.880 1192.230 766.160 ;
        RECT 1192.870 765.880 1193.150 766.160 ;
      LAYER met3 ;
        RECT 1192.385 1200.690 1192.715 1200.705 ;
        RECT 1193.305 1200.690 1193.635 1200.705 ;
        RECT 1192.385 1200.390 1193.635 1200.690 ;
        RECT 1192.385 1200.375 1192.715 1200.390 ;
        RECT 1193.305 1200.375 1193.635 1200.390 ;
        RECT 1192.385 1104.130 1192.715 1104.145 ;
        RECT 1193.305 1104.130 1193.635 1104.145 ;
        RECT 1192.385 1103.830 1193.635 1104.130 ;
        RECT 1192.385 1103.815 1192.715 1103.830 ;
        RECT 1193.305 1103.815 1193.635 1103.830 ;
        RECT 1192.385 1055.850 1192.715 1055.865 ;
        RECT 1193.305 1055.850 1193.635 1055.865 ;
        RECT 1192.385 1055.550 1193.635 1055.850 ;
        RECT 1192.385 1055.535 1192.715 1055.550 ;
        RECT 1193.305 1055.535 1193.635 1055.550 ;
        RECT 1192.385 1007.570 1192.715 1007.585 ;
        RECT 1193.305 1007.570 1193.635 1007.585 ;
        RECT 1192.385 1007.270 1193.635 1007.570 ;
        RECT 1192.385 1007.255 1192.715 1007.270 ;
        RECT 1193.305 1007.255 1193.635 1007.270 ;
        RECT 1191.925 766.170 1192.255 766.185 ;
        RECT 1192.845 766.170 1193.175 766.185 ;
        RECT 1191.925 765.870 1193.175 766.170 ;
        RECT 1191.925 765.855 1192.255 765.870 ;
        RECT 1192.845 765.855 1193.175 765.870 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1366.805 138.125 1366.975 159.375 ;
        RECT 1318.045 17.765 1318.215 18.955 ;
        RECT 1342.425 18.105 1342.595 18.955 ;
      LAYER mcon ;
        RECT 1366.805 159.205 1366.975 159.375 ;
        RECT 1318.045 18.785 1318.215 18.955 ;
        RECT 1342.425 18.785 1342.595 18.955 ;
      LAYER met1 ;
        RECT 1366.730 159.360 1367.050 159.420 ;
        RECT 1366.535 159.220 1367.050 159.360 ;
        RECT 1366.730 159.160 1367.050 159.220 ;
        RECT 1366.730 138.280 1367.050 138.340 ;
        RECT 1366.535 138.140 1367.050 138.280 ;
        RECT 1366.730 138.080 1367.050 138.140 ;
        RECT 1317.985 18.940 1318.275 18.985 ;
        RECT 1342.365 18.940 1342.655 18.985 ;
        RECT 1317.985 18.800 1342.655 18.940 ;
        RECT 1317.985 18.755 1318.275 18.800 ;
        RECT 1342.365 18.755 1342.655 18.800 ;
        RECT 1342.365 18.260 1342.655 18.305 ;
        RECT 1366.270 18.260 1366.590 18.320 ;
        RECT 1342.365 18.120 1366.590 18.260 ;
        RECT 1342.365 18.075 1342.655 18.120 ;
        RECT 1366.270 18.060 1366.590 18.120 ;
        RECT 1209.870 17.920 1210.190 17.980 ;
        RECT 1317.985 17.920 1318.275 17.965 ;
        RECT 1209.870 17.780 1318.275 17.920 ;
        RECT 1209.870 17.720 1210.190 17.780 ;
        RECT 1317.985 17.735 1318.275 17.780 ;
      LAYER via ;
        RECT 1366.760 159.160 1367.020 159.420 ;
        RECT 1366.760 138.080 1367.020 138.340 ;
        RECT 1366.300 18.060 1366.560 18.320 ;
        RECT 1209.900 17.720 1210.160 17.980 ;
      LAYER met2 ;
        RECT 1371.370 1220.330 1371.930 1228.680 ;
        RECT 1369.580 1220.190 1371.930 1220.330 ;
        RECT 1369.580 1196.700 1369.720 1220.190 ;
        RECT 1371.370 1219.680 1371.930 1220.190 ;
        RECT 1366.360 1196.560 1369.720 1196.700 ;
        RECT 1366.360 1172.730 1366.500 1196.560 ;
        RECT 1366.360 1172.590 1366.960 1172.730 ;
        RECT 1366.820 1028.570 1366.960 1172.590 ;
        RECT 1366.360 1028.430 1366.960 1028.570 ;
        RECT 1366.360 1027.890 1366.500 1028.430 ;
        RECT 1366.360 1027.750 1366.960 1027.890 ;
        RECT 1366.820 932.010 1366.960 1027.750 ;
        RECT 1366.360 931.870 1366.960 932.010 ;
        RECT 1366.360 931.330 1366.500 931.870 ;
        RECT 1366.360 931.190 1366.960 931.330 ;
        RECT 1366.820 835.450 1366.960 931.190 ;
        RECT 1366.360 835.310 1366.960 835.450 ;
        RECT 1366.360 834.770 1366.500 835.310 ;
        RECT 1366.360 834.630 1366.960 834.770 ;
        RECT 1366.820 738.890 1366.960 834.630 ;
        RECT 1366.360 738.750 1366.960 738.890 ;
        RECT 1366.360 738.210 1366.500 738.750 ;
        RECT 1366.360 738.070 1366.960 738.210 ;
        RECT 1366.820 642.330 1366.960 738.070 ;
        RECT 1366.360 642.190 1366.960 642.330 ;
        RECT 1366.360 641.650 1366.500 642.190 ;
        RECT 1366.360 641.510 1366.960 641.650 ;
        RECT 1366.820 545.770 1366.960 641.510 ;
        RECT 1366.360 545.630 1366.960 545.770 ;
        RECT 1366.360 545.090 1366.500 545.630 ;
        RECT 1366.360 544.950 1366.960 545.090 ;
        RECT 1366.820 449.210 1366.960 544.950 ;
        RECT 1366.360 449.070 1366.960 449.210 ;
        RECT 1366.360 448.530 1366.500 449.070 ;
        RECT 1366.360 448.390 1366.960 448.530 ;
        RECT 1366.820 351.970 1366.960 448.390 ;
        RECT 1366.360 351.830 1366.960 351.970 ;
        RECT 1366.360 351.290 1366.500 351.830 ;
        RECT 1366.360 351.150 1366.960 351.290 ;
        RECT 1366.820 255.410 1366.960 351.150 ;
        RECT 1366.360 255.270 1366.960 255.410 ;
        RECT 1366.360 254.730 1366.500 255.270 ;
        RECT 1366.360 254.590 1366.960 254.730 ;
        RECT 1366.820 159.450 1366.960 254.590 ;
        RECT 1366.760 159.130 1367.020 159.450 ;
        RECT 1366.760 138.050 1367.020 138.370 ;
        RECT 1366.820 96.290 1366.960 138.050 ;
        RECT 1366.360 96.150 1366.960 96.290 ;
        RECT 1366.360 18.350 1366.500 96.150 ;
        RECT 1366.300 18.030 1366.560 18.350 ;
        RECT 1209.900 17.690 1210.160 18.010 ;
        RECT 1209.960 2.400 1210.100 17.690 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1356.685 1208.105 1356.855 1213.715 ;
      LAYER mcon ;
        RECT 1356.685 1213.545 1356.855 1213.715 ;
      LAYER met1 ;
        RECT 1228.270 1213.700 1228.590 1213.760 ;
        RECT 1356.625 1213.700 1356.915 1213.745 ;
        RECT 1228.270 1213.560 1356.915 1213.700 ;
        RECT 1228.270 1213.500 1228.590 1213.560 ;
        RECT 1356.625 1213.515 1356.915 1213.560 ;
        RECT 1356.625 1208.260 1356.915 1208.305 ;
        RECT 1356.625 1208.120 1372.480 1208.260 ;
        RECT 1356.625 1208.075 1356.915 1208.120 ;
        RECT 1372.340 1207.920 1372.480 1208.120 ;
        RECT 1380.530 1207.920 1380.850 1207.980 ;
        RECT 1372.340 1207.780 1380.850 1207.920 ;
        RECT 1380.530 1207.720 1380.850 1207.780 ;
      LAYER via ;
        RECT 1228.300 1213.500 1228.560 1213.760 ;
        RECT 1380.560 1207.720 1380.820 1207.980 ;
      LAYER met2 ;
        RECT 1380.570 1219.680 1381.130 1228.680 ;
        RECT 1228.300 1213.470 1228.560 1213.790 ;
        RECT 1228.360 1212.850 1228.500 1213.470 ;
        RECT 1227.900 1212.710 1228.500 1212.850 ;
        RECT 1227.900 2.400 1228.040 1212.710 ;
        RECT 1380.620 1208.010 1380.760 1219.680 ;
        RECT 1380.560 1207.690 1380.820 1208.010 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 1211.660 1248.830 1211.720 ;
        RECT 1389.730 1211.660 1390.050 1211.720 ;
        RECT 1248.510 1211.520 1390.050 1211.660 ;
        RECT 1248.510 1211.460 1248.830 1211.520 ;
        RECT 1389.730 1211.460 1390.050 1211.520 ;
        RECT 1245.750 18.940 1246.070 19.000 ;
        RECT 1248.510 18.940 1248.830 19.000 ;
        RECT 1245.750 18.800 1248.830 18.940 ;
        RECT 1245.750 18.740 1246.070 18.800 ;
        RECT 1248.510 18.740 1248.830 18.800 ;
      LAYER via ;
        RECT 1248.540 1211.460 1248.800 1211.720 ;
        RECT 1389.760 1211.460 1390.020 1211.720 ;
        RECT 1245.780 18.740 1246.040 19.000 ;
        RECT 1248.540 18.740 1248.800 19.000 ;
      LAYER met2 ;
        RECT 1389.770 1219.680 1390.330 1228.680 ;
        RECT 1389.820 1211.750 1389.960 1219.680 ;
        RECT 1248.540 1211.430 1248.800 1211.750 ;
        RECT 1389.760 1211.430 1390.020 1211.750 ;
        RECT 1248.600 19.030 1248.740 1211.430 ;
        RECT 1245.780 18.710 1246.040 19.030 ;
        RECT 1248.540 18.710 1248.800 19.030 ;
        RECT 1245.840 2.400 1245.980 18.710 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1394.405 1110.865 1394.575 1125.315 ;
      LAYER mcon ;
        RECT 1394.405 1125.145 1394.575 1125.315 ;
      LAYER met1 ;
        RECT 1394.345 1125.300 1394.635 1125.345 ;
        RECT 1394.790 1125.300 1395.110 1125.360 ;
        RECT 1394.345 1125.160 1395.110 1125.300 ;
        RECT 1394.345 1125.115 1394.635 1125.160 ;
        RECT 1394.790 1125.100 1395.110 1125.160 ;
        RECT 1394.330 1111.020 1394.650 1111.080 ;
        RECT 1394.135 1110.880 1394.650 1111.020 ;
        RECT 1394.330 1110.820 1394.650 1110.880 ;
        RECT 1394.330 1076.480 1394.650 1076.740 ;
        RECT 1394.420 1076.060 1394.560 1076.480 ;
        RECT 1394.330 1075.800 1394.650 1076.060 ;
        RECT 1394.330 303.320 1394.650 303.580 ;
        RECT 1394.420 303.180 1394.560 303.320 ;
        RECT 1394.790 303.180 1395.110 303.240 ;
        RECT 1394.420 303.040 1395.110 303.180 ;
        RECT 1394.790 302.980 1395.110 303.040 ;
        RECT 1263.230 18.600 1263.550 18.660 ;
        RECT 1394.330 18.600 1394.650 18.660 ;
        RECT 1263.230 18.460 1394.650 18.600 ;
        RECT 1263.230 18.400 1263.550 18.460 ;
        RECT 1394.330 18.400 1394.650 18.460 ;
      LAYER via ;
        RECT 1394.820 1125.100 1395.080 1125.360 ;
        RECT 1394.360 1110.820 1394.620 1111.080 ;
        RECT 1394.360 1076.480 1394.620 1076.740 ;
        RECT 1394.360 1075.800 1394.620 1076.060 ;
        RECT 1394.360 303.320 1394.620 303.580 ;
        RECT 1394.820 302.980 1395.080 303.240 ;
        RECT 1263.260 18.400 1263.520 18.660 ;
        RECT 1394.360 18.400 1394.620 18.660 ;
      LAYER met2 ;
        RECT 1398.970 1220.330 1399.530 1228.680 ;
        RECT 1397.180 1220.190 1399.530 1220.330 ;
        RECT 1397.180 1196.700 1397.320 1220.190 ;
        RECT 1398.970 1219.680 1399.530 1220.190 ;
        RECT 1393.960 1196.560 1397.320 1196.700 ;
        RECT 1393.960 1172.730 1394.100 1196.560 ;
        RECT 1393.960 1172.590 1395.020 1172.730 ;
        RECT 1394.880 1125.390 1395.020 1172.590 ;
        RECT 1394.820 1125.070 1395.080 1125.390 ;
        RECT 1394.360 1110.790 1394.620 1111.110 ;
        RECT 1394.420 1076.770 1394.560 1110.790 ;
        RECT 1394.360 1076.450 1394.620 1076.770 ;
        RECT 1394.360 1075.770 1394.620 1076.090 ;
        RECT 1394.420 1028.570 1394.560 1075.770 ;
        RECT 1393.960 1028.430 1394.560 1028.570 ;
        RECT 1393.960 1027.890 1394.100 1028.430 ;
        RECT 1393.960 1027.750 1394.560 1027.890 ;
        RECT 1394.420 932.010 1394.560 1027.750 ;
        RECT 1393.960 931.870 1394.560 932.010 ;
        RECT 1393.960 931.330 1394.100 931.870 ;
        RECT 1393.960 931.190 1394.560 931.330 ;
        RECT 1394.420 835.450 1394.560 931.190 ;
        RECT 1393.960 835.310 1394.560 835.450 ;
        RECT 1393.960 834.770 1394.100 835.310 ;
        RECT 1393.960 834.630 1394.560 834.770 ;
        RECT 1394.420 738.890 1394.560 834.630 ;
        RECT 1393.960 738.750 1394.560 738.890 ;
        RECT 1393.960 738.210 1394.100 738.750 ;
        RECT 1393.960 738.070 1394.560 738.210 ;
        RECT 1394.420 642.330 1394.560 738.070 ;
        RECT 1393.960 642.190 1394.560 642.330 ;
        RECT 1393.960 641.650 1394.100 642.190 ;
        RECT 1393.960 641.510 1394.560 641.650 ;
        RECT 1394.420 545.770 1394.560 641.510 ;
        RECT 1393.960 545.630 1394.560 545.770 ;
        RECT 1393.960 545.090 1394.100 545.630 ;
        RECT 1393.960 544.950 1394.560 545.090 ;
        RECT 1394.420 449.210 1394.560 544.950 ;
        RECT 1393.960 449.070 1394.560 449.210 ;
        RECT 1393.960 448.530 1394.100 449.070 ;
        RECT 1393.960 448.390 1394.560 448.530 ;
        RECT 1394.420 351.970 1394.560 448.390 ;
        RECT 1393.960 351.830 1394.560 351.970 ;
        RECT 1393.960 351.290 1394.100 351.830 ;
        RECT 1393.960 351.150 1394.560 351.290 ;
        RECT 1394.420 303.610 1394.560 351.150 ;
        RECT 1394.360 303.290 1394.620 303.610 ;
        RECT 1394.820 302.950 1395.080 303.270 ;
        RECT 1394.880 207.810 1395.020 302.950 ;
        RECT 1394.420 207.670 1395.020 207.810 ;
        RECT 1394.420 207.130 1394.560 207.670 ;
        RECT 1393.960 206.990 1394.560 207.130 ;
        RECT 1393.960 206.450 1394.100 206.990 ;
        RECT 1393.960 206.310 1394.560 206.450 ;
        RECT 1394.420 110.570 1394.560 206.310 ;
        RECT 1393.960 110.430 1394.560 110.570 ;
        RECT 1393.960 109.890 1394.100 110.430 ;
        RECT 1393.960 109.750 1394.560 109.890 ;
        RECT 1394.420 18.690 1394.560 109.750 ;
        RECT 1263.260 18.370 1263.520 18.690 ;
        RECT 1394.360 18.370 1394.620 18.690 ;
        RECT 1263.320 2.400 1263.460 18.370 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.470 1212.680 1283.790 1212.740 ;
        RECT 1407.670 1212.680 1407.990 1212.740 ;
        RECT 1283.470 1212.540 1407.990 1212.680 ;
        RECT 1283.470 1212.480 1283.790 1212.540 ;
        RECT 1407.670 1212.480 1407.990 1212.540 ;
        RECT 1281.170 2.960 1281.490 3.020 ;
        RECT 1283.010 2.960 1283.330 3.020 ;
        RECT 1281.170 2.820 1283.330 2.960 ;
        RECT 1281.170 2.760 1281.490 2.820 ;
        RECT 1283.010 2.760 1283.330 2.820 ;
      LAYER via ;
        RECT 1283.500 1212.480 1283.760 1212.740 ;
        RECT 1407.700 1212.480 1407.960 1212.740 ;
        RECT 1281.200 2.760 1281.460 3.020 ;
        RECT 1283.040 2.760 1283.300 3.020 ;
      LAYER met2 ;
        RECT 1407.710 1219.680 1408.270 1228.680 ;
        RECT 1407.760 1212.770 1407.900 1219.680 ;
        RECT 1283.500 1212.450 1283.760 1212.770 ;
        RECT 1407.700 1212.450 1407.960 1212.770 ;
        RECT 1283.560 1212.170 1283.700 1212.450 ;
        RECT 1283.100 1212.030 1283.700 1212.170 ;
        RECT 1283.100 3.050 1283.240 1212.030 ;
        RECT 1281.200 2.730 1281.460 3.050 ;
        RECT 1283.040 2.730 1283.300 3.050 ;
        RECT 1281.260 2.400 1281.400 2.730 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1403.990 1207.580 1404.310 1207.640 ;
        RECT 1416.870 1207.580 1417.190 1207.640 ;
        RECT 1403.990 1207.440 1417.190 1207.580 ;
        RECT 1403.990 1207.380 1404.310 1207.440 ;
        RECT 1416.870 1207.380 1417.190 1207.440 ;
        RECT 1299.110 16.560 1299.430 16.620 ;
        RECT 1403.990 16.560 1404.310 16.620 ;
        RECT 1299.110 16.420 1404.310 16.560 ;
        RECT 1299.110 16.360 1299.430 16.420 ;
        RECT 1403.990 16.360 1404.310 16.420 ;
      LAYER via ;
        RECT 1404.020 1207.380 1404.280 1207.640 ;
        RECT 1416.900 1207.380 1417.160 1207.640 ;
        RECT 1299.140 16.360 1299.400 16.620 ;
        RECT 1404.020 16.360 1404.280 16.620 ;
      LAYER met2 ;
        RECT 1416.910 1219.680 1417.470 1228.680 ;
        RECT 1416.960 1207.670 1417.100 1219.680 ;
        RECT 1404.020 1207.350 1404.280 1207.670 ;
        RECT 1416.900 1207.350 1417.160 1207.670 ;
        RECT 1404.080 16.650 1404.220 1207.350 ;
        RECT 1299.140 16.330 1299.400 16.650 ;
        RECT 1404.020 16.330 1404.280 16.650 ;
        RECT 1299.200 2.400 1299.340 16.330 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1422.005 786.505 1422.175 821.015 ;
        RECT 1422.005 689.605 1422.175 724.455 ;
        RECT 1422.005 593.045 1422.175 627.895 ;
        RECT 1422.005 496.485 1422.175 531.335 ;
        RECT 1422.005 386.325 1422.175 434.775 ;
        RECT 1422.465 206.805 1422.635 241.315 ;
        RECT 1422.005 144.925 1422.175 193.035 ;
      LAYER mcon ;
        RECT 1422.005 820.845 1422.175 821.015 ;
        RECT 1422.005 724.285 1422.175 724.455 ;
        RECT 1422.005 627.725 1422.175 627.895 ;
        RECT 1422.005 531.165 1422.175 531.335 ;
        RECT 1422.005 434.605 1422.175 434.775 ;
        RECT 1422.465 241.145 1422.635 241.315 ;
        RECT 1422.005 192.865 1422.175 193.035 ;
      LAYER met1 ;
        RECT 1421.470 1028.400 1421.790 1028.460 ;
        RECT 1422.390 1028.400 1422.710 1028.460 ;
        RECT 1421.470 1028.260 1422.710 1028.400 ;
        RECT 1421.470 1028.200 1421.790 1028.260 ;
        RECT 1422.390 1028.200 1422.710 1028.260 ;
        RECT 1421.470 931.840 1421.790 931.900 ;
        RECT 1422.390 931.840 1422.710 931.900 ;
        RECT 1421.470 931.700 1422.710 931.840 ;
        RECT 1421.470 931.640 1421.790 931.700 ;
        RECT 1422.390 931.640 1422.710 931.700 ;
        RECT 1422.390 869.620 1422.710 869.680 ;
        RECT 1423.310 869.620 1423.630 869.680 ;
        RECT 1422.390 869.480 1423.630 869.620 ;
        RECT 1422.390 869.420 1422.710 869.480 ;
        RECT 1423.310 869.420 1423.630 869.480 ;
        RECT 1421.470 835.280 1421.790 835.340 ;
        RECT 1422.390 835.280 1422.710 835.340 ;
        RECT 1421.470 835.140 1422.710 835.280 ;
        RECT 1421.470 835.080 1421.790 835.140 ;
        RECT 1422.390 835.080 1422.710 835.140 ;
        RECT 1421.930 821.000 1422.250 821.060 ;
        RECT 1421.735 820.860 1422.250 821.000 ;
        RECT 1421.930 820.800 1422.250 820.860 ;
        RECT 1421.930 786.660 1422.250 786.720 ;
        RECT 1421.735 786.520 1422.250 786.660 ;
        RECT 1421.930 786.460 1422.250 786.520 ;
        RECT 1421.470 738.380 1421.790 738.440 ;
        RECT 1422.390 738.380 1422.710 738.440 ;
        RECT 1421.470 738.240 1422.710 738.380 ;
        RECT 1421.470 738.180 1421.790 738.240 ;
        RECT 1422.390 738.180 1422.710 738.240 ;
        RECT 1421.930 724.440 1422.250 724.500 ;
        RECT 1421.735 724.300 1422.250 724.440 ;
        RECT 1421.930 724.240 1422.250 724.300 ;
        RECT 1421.930 689.760 1422.250 689.820 ;
        RECT 1421.735 689.620 1422.250 689.760 ;
        RECT 1421.930 689.560 1422.250 689.620 ;
        RECT 1421.470 641.820 1421.790 641.880 ;
        RECT 1422.390 641.820 1422.710 641.880 ;
        RECT 1421.470 641.680 1422.710 641.820 ;
        RECT 1421.470 641.620 1421.790 641.680 ;
        RECT 1422.390 641.620 1422.710 641.680 ;
        RECT 1421.930 627.880 1422.250 627.940 ;
        RECT 1421.735 627.740 1422.250 627.880 ;
        RECT 1421.930 627.680 1422.250 627.740 ;
        RECT 1421.930 593.200 1422.250 593.260 ;
        RECT 1421.735 593.060 1422.250 593.200 ;
        RECT 1421.930 593.000 1422.250 593.060 ;
        RECT 1421.470 545.260 1421.790 545.320 ;
        RECT 1422.390 545.260 1422.710 545.320 ;
        RECT 1421.470 545.120 1422.710 545.260 ;
        RECT 1421.470 545.060 1421.790 545.120 ;
        RECT 1422.390 545.060 1422.710 545.120 ;
        RECT 1421.930 531.320 1422.250 531.380 ;
        RECT 1421.735 531.180 1422.250 531.320 ;
        RECT 1421.930 531.120 1422.250 531.180 ;
        RECT 1421.930 496.640 1422.250 496.700 ;
        RECT 1421.735 496.500 1422.250 496.640 ;
        RECT 1421.930 496.440 1422.250 496.500 ;
        RECT 1421.470 448.700 1421.790 448.760 ;
        RECT 1422.390 448.700 1422.710 448.760 ;
        RECT 1421.470 448.560 1422.710 448.700 ;
        RECT 1421.470 448.500 1421.790 448.560 ;
        RECT 1422.390 448.500 1422.710 448.560 ;
        RECT 1421.930 434.760 1422.250 434.820 ;
        RECT 1421.735 434.620 1422.250 434.760 ;
        RECT 1421.930 434.560 1422.250 434.620 ;
        RECT 1421.945 386.480 1422.235 386.525 ;
        RECT 1422.390 386.480 1422.710 386.540 ;
        RECT 1421.945 386.340 1422.710 386.480 ;
        RECT 1421.945 386.295 1422.235 386.340 ;
        RECT 1422.390 386.280 1422.710 386.340 ;
        RECT 1421.930 331.400 1422.250 331.460 ;
        RECT 1422.390 331.400 1422.710 331.460 ;
        RECT 1421.930 331.260 1422.710 331.400 ;
        RECT 1421.930 331.200 1422.250 331.260 ;
        RECT 1422.390 331.200 1422.710 331.260 ;
        RECT 1421.930 304.000 1422.250 304.260 ;
        RECT 1422.020 303.580 1422.160 304.000 ;
        RECT 1421.930 303.320 1422.250 303.580 ;
        RECT 1421.930 255.580 1422.250 255.640 ;
        RECT 1421.560 255.440 1422.250 255.580 ;
        RECT 1421.560 255.300 1421.700 255.440 ;
        RECT 1421.930 255.380 1422.250 255.440 ;
        RECT 1421.470 255.040 1421.790 255.300 ;
        RECT 1421.470 241.300 1421.790 241.360 ;
        RECT 1422.405 241.300 1422.695 241.345 ;
        RECT 1421.470 241.160 1422.695 241.300 ;
        RECT 1421.470 241.100 1421.790 241.160 ;
        RECT 1422.405 241.115 1422.695 241.160 ;
        RECT 1422.390 206.960 1422.710 207.020 ;
        RECT 1422.195 206.820 1422.710 206.960 ;
        RECT 1422.390 206.760 1422.710 206.820 ;
        RECT 1421.945 193.020 1422.235 193.065 ;
        RECT 1422.390 193.020 1422.710 193.080 ;
        RECT 1421.945 192.880 1422.710 193.020 ;
        RECT 1421.945 192.835 1422.235 192.880 ;
        RECT 1422.390 192.820 1422.710 192.880 ;
        RECT 1421.930 145.080 1422.250 145.140 ;
        RECT 1421.735 144.940 1422.250 145.080 ;
        RECT 1421.930 144.880 1422.250 144.940 ;
        RECT 1317.050 19.620 1317.370 19.680 ;
        RECT 1422.390 19.620 1422.710 19.680 ;
        RECT 1317.050 19.480 1422.710 19.620 ;
        RECT 1317.050 19.420 1317.370 19.480 ;
        RECT 1422.390 19.420 1422.710 19.480 ;
      LAYER via ;
        RECT 1421.500 1028.200 1421.760 1028.460 ;
        RECT 1422.420 1028.200 1422.680 1028.460 ;
        RECT 1421.500 931.640 1421.760 931.900 ;
        RECT 1422.420 931.640 1422.680 931.900 ;
        RECT 1422.420 869.420 1422.680 869.680 ;
        RECT 1423.340 869.420 1423.600 869.680 ;
        RECT 1421.500 835.080 1421.760 835.340 ;
        RECT 1422.420 835.080 1422.680 835.340 ;
        RECT 1421.960 820.800 1422.220 821.060 ;
        RECT 1421.960 786.460 1422.220 786.720 ;
        RECT 1421.500 738.180 1421.760 738.440 ;
        RECT 1422.420 738.180 1422.680 738.440 ;
        RECT 1421.960 724.240 1422.220 724.500 ;
        RECT 1421.960 689.560 1422.220 689.820 ;
        RECT 1421.500 641.620 1421.760 641.880 ;
        RECT 1422.420 641.620 1422.680 641.880 ;
        RECT 1421.960 627.680 1422.220 627.940 ;
        RECT 1421.960 593.000 1422.220 593.260 ;
        RECT 1421.500 545.060 1421.760 545.320 ;
        RECT 1422.420 545.060 1422.680 545.320 ;
        RECT 1421.960 531.120 1422.220 531.380 ;
        RECT 1421.960 496.440 1422.220 496.700 ;
        RECT 1421.500 448.500 1421.760 448.760 ;
        RECT 1422.420 448.500 1422.680 448.760 ;
        RECT 1421.960 434.560 1422.220 434.820 ;
        RECT 1422.420 386.280 1422.680 386.540 ;
        RECT 1421.960 331.200 1422.220 331.460 ;
        RECT 1422.420 331.200 1422.680 331.460 ;
        RECT 1421.960 304.000 1422.220 304.260 ;
        RECT 1421.960 303.320 1422.220 303.580 ;
        RECT 1421.960 255.380 1422.220 255.640 ;
        RECT 1421.500 255.040 1421.760 255.300 ;
        RECT 1421.500 241.100 1421.760 241.360 ;
        RECT 1422.420 206.760 1422.680 207.020 ;
        RECT 1422.420 192.820 1422.680 193.080 ;
        RECT 1421.960 144.880 1422.220 145.140 ;
        RECT 1317.080 19.420 1317.340 19.680 ;
        RECT 1422.420 19.420 1422.680 19.680 ;
      LAYER met2 ;
        RECT 1426.110 1220.330 1426.670 1228.680 ;
        RECT 1424.780 1220.190 1426.670 1220.330 ;
        RECT 1424.780 1214.890 1424.920 1220.190 ;
        RECT 1426.110 1219.680 1426.670 1220.190 ;
        RECT 1423.860 1214.750 1424.920 1214.890 ;
        RECT 1423.860 1206.730 1424.000 1214.750 ;
        RECT 1421.560 1206.590 1424.000 1206.730 ;
        RECT 1421.560 1172.730 1421.700 1206.590 ;
        RECT 1421.560 1172.590 1422.160 1172.730 ;
        RECT 1422.020 1125.130 1422.160 1172.590 ;
        RECT 1422.020 1124.990 1422.620 1125.130 ;
        RECT 1422.480 1028.490 1422.620 1124.990 ;
        RECT 1421.500 1028.170 1421.760 1028.490 ;
        RECT 1422.420 1028.170 1422.680 1028.490 ;
        RECT 1421.560 1027.890 1421.700 1028.170 ;
        RECT 1421.560 1027.750 1422.160 1027.890 ;
        RECT 1422.020 980.290 1422.160 1027.750 ;
        RECT 1422.020 980.150 1422.620 980.290 ;
        RECT 1422.480 931.930 1422.620 980.150 ;
        RECT 1421.500 931.610 1421.760 931.930 ;
        RECT 1422.420 931.610 1422.680 931.930 ;
        RECT 1421.560 931.330 1421.700 931.610 ;
        RECT 1421.560 931.190 1422.160 931.330 ;
        RECT 1422.020 917.845 1422.160 931.190 ;
        RECT 1421.950 917.475 1422.230 917.845 ;
        RECT 1423.330 917.475 1423.610 917.845 ;
        RECT 1423.400 869.710 1423.540 917.475 ;
        RECT 1422.420 869.390 1422.680 869.710 ;
        RECT 1423.340 869.390 1423.600 869.710 ;
        RECT 1422.480 835.370 1422.620 869.390 ;
        RECT 1421.500 835.050 1421.760 835.370 ;
        RECT 1422.420 835.050 1422.680 835.370 ;
        RECT 1421.560 834.770 1421.700 835.050 ;
        RECT 1421.560 834.630 1422.160 834.770 ;
        RECT 1422.020 821.090 1422.160 834.630 ;
        RECT 1421.960 820.770 1422.220 821.090 ;
        RECT 1421.960 786.430 1422.220 786.750 ;
        RECT 1422.020 772.890 1422.160 786.430 ;
        RECT 1422.020 772.750 1422.620 772.890 ;
        RECT 1422.480 738.470 1422.620 772.750 ;
        RECT 1421.500 738.210 1421.760 738.470 ;
        RECT 1421.500 738.150 1422.160 738.210 ;
        RECT 1422.420 738.150 1422.680 738.470 ;
        RECT 1421.560 738.070 1422.160 738.150 ;
        RECT 1422.020 724.530 1422.160 738.070 ;
        RECT 1421.960 724.210 1422.220 724.530 ;
        RECT 1421.960 689.530 1422.220 689.850 ;
        RECT 1422.020 676.330 1422.160 689.530 ;
        RECT 1422.020 676.190 1422.620 676.330 ;
        RECT 1422.480 641.910 1422.620 676.190 ;
        RECT 1421.500 641.650 1421.760 641.910 ;
        RECT 1421.500 641.590 1422.160 641.650 ;
        RECT 1422.420 641.590 1422.680 641.910 ;
        RECT 1421.560 641.510 1422.160 641.590 ;
        RECT 1422.020 627.970 1422.160 641.510 ;
        RECT 1421.960 627.650 1422.220 627.970 ;
        RECT 1421.960 592.970 1422.220 593.290 ;
        RECT 1422.020 579.770 1422.160 592.970 ;
        RECT 1422.020 579.630 1422.620 579.770 ;
        RECT 1422.480 545.350 1422.620 579.630 ;
        RECT 1421.500 545.090 1421.760 545.350 ;
        RECT 1421.500 545.030 1422.160 545.090 ;
        RECT 1422.420 545.030 1422.680 545.350 ;
        RECT 1421.560 544.950 1422.160 545.030 ;
        RECT 1422.020 531.410 1422.160 544.950 ;
        RECT 1421.960 531.090 1422.220 531.410 ;
        RECT 1421.960 496.410 1422.220 496.730 ;
        RECT 1422.020 483.210 1422.160 496.410 ;
        RECT 1422.020 483.070 1422.620 483.210 ;
        RECT 1422.480 448.790 1422.620 483.070 ;
        RECT 1421.500 448.530 1421.760 448.790 ;
        RECT 1421.500 448.470 1422.160 448.530 ;
        RECT 1422.420 448.470 1422.680 448.790 ;
        RECT 1421.560 448.390 1422.160 448.470 ;
        RECT 1422.020 434.850 1422.160 448.390 ;
        RECT 1421.960 434.530 1422.220 434.850 ;
        RECT 1422.420 386.250 1422.680 386.570 ;
        RECT 1422.480 331.490 1422.620 386.250 ;
        RECT 1421.960 331.170 1422.220 331.490 ;
        RECT 1422.420 331.170 1422.680 331.490 ;
        RECT 1422.020 304.290 1422.160 331.170 ;
        RECT 1421.960 303.970 1422.220 304.290 ;
        RECT 1421.960 303.290 1422.220 303.610 ;
        RECT 1422.020 255.670 1422.160 303.290 ;
        RECT 1421.960 255.350 1422.220 255.670 ;
        RECT 1421.500 255.010 1421.760 255.330 ;
        RECT 1421.560 241.390 1421.700 255.010 ;
        RECT 1421.500 241.070 1421.760 241.390 ;
        RECT 1422.420 206.730 1422.680 207.050 ;
        RECT 1422.480 193.110 1422.620 206.730 ;
        RECT 1422.420 192.790 1422.680 193.110 ;
        RECT 1421.960 144.850 1422.220 145.170 ;
        RECT 1422.020 120.770 1422.160 144.850 ;
        RECT 1422.020 120.630 1422.620 120.770 ;
        RECT 1422.480 19.710 1422.620 120.630 ;
        RECT 1317.080 19.390 1317.340 19.710 ;
        RECT 1422.420 19.390 1422.680 19.710 ;
        RECT 1317.140 2.400 1317.280 19.390 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1421.950 917.520 1422.230 917.800 ;
        RECT 1423.330 917.520 1423.610 917.800 ;
      LAYER met3 ;
        RECT 1421.925 917.810 1422.255 917.825 ;
        RECT 1423.305 917.810 1423.635 917.825 ;
        RECT 1421.925 917.510 1423.635 917.810 ;
        RECT 1421.925 917.495 1422.255 917.510 ;
        RECT 1423.305 917.495 1423.635 917.510 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 1210.640 1338.530 1210.700 ;
        RECT 1435.270 1210.640 1435.590 1210.700 ;
        RECT 1338.210 1210.500 1435.590 1210.640 ;
        RECT 1338.210 1210.440 1338.530 1210.500 ;
        RECT 1435.270 1210.440 1435.590 1210.500 ;
        RECT 1334.990 15.540 1335.310 15.600 ;
        RECT 1338.210 15.540 1338.530 15.600 ;
        RECT 1334.990 15.400 1338.530 15.540 ;
        RECT 1334.990 15.340 1335.310 15.400 ;
        RECT 1338.210 15.340 1338.530 15.400 ;
      LAYER via ;
        RECT 1338.240 1210.440 1338.500 1210.700 ;
        RECT 1435.300 1210.440 1435.560 1210.700 ;
        RECT 1335.020 15.340 1335.280 15.600 ;
        RECT 1338.240 15.340 1338.500 15.600 ;
      LAYER met2 ;
        RECT 1435.310 1219.680 1435.870 1228.680 ;
        RECT 1435.360 1210.730 1435.500 1219.680 ;
        RECT 1338.240 1210.410 1338.500 1210.730 ;
        RECT 1435.300 1210.410 1435.560 1210.730 ;
        RECT 1338.300 15.630 1338.440 1210.410 ;
        RECT 1335.020 15.310 1335.280 15.630 ;
        RECT 1338.240 15.310 1338.500 15.630 ;
        RECT 1335.080 2.400 1335.220 15.310 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 42.740 692.690 42.800 ;
        RECT 1104.530 42.740 1104.850 42.800 ;
        RECT 692.370 42.600 1104.850 42.740 ;
        RECT 692.370 42.540 692.690 42.600 ;
        RECT 1104.530 42.540 1104.850 42.600 ;
      LAYER via ;
        RECT 692.400 42.540 692.660 42.800 ;
        RECT 1104.560 42.540 1104.820 42.800 ;
      LAYER met2 ;
        RECT 1105.490 1220.330 1106.050 1228.680 ;
        RECT 1104.620 1220.190 1106.050 1220.330 ;
        RECT 1104.620 42.830 1104.760 1220.190 ;
        RECT 1105.490 1219.680 1106.050 1220.190 ;
        RECT 692.400 42.510 692.660 42.830 ;
        RECT 1104.560 42.510 1104.820 42.830 ;
        RECT 692.460 2.400 692.600 42.510 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1424.690 1214.040 1425.010 1214.100 ;
        RECT 1444.470 1214.040 1444.790 1214.100 ;
        RECT 1424.690 1213.900 1444.790 1214.040 ;
        RECT 1424.690 1213.840 1425.010 1213.900 ;
        RECT 1444.470 1213.840 1444.790 1213.900 ;
        RECT 1352.470 17.240 1352.790 17.300 ;
        RECT 1352.470 17.100 1382.140 17.240 ;
        RECT 1352.470 17.040 1352.790 17.100 ;
        RECT 1382.000 16.900 1382.140 17.100 ;
        RECT 1424.690 16.900 1425.010 16.960 ;
        RECT 1382.000 16.760 1425.010 16.900 ;
        RECT 1424.690 16.700 1425.010 16.760 ;
      LAYER via ;
        RECT 1424.720 1213.840 1424.980 1214.100 ;
        RECT 1444.500 1213.840 1444.760 1214.100 ;
        RECT 1352.500 17.040 1352.760 17.300 ;
        RECT 1424.720 16.700 1424.980 16.960 ;
      LAYER met2 ;
        RECT 1444.510 1219.680 1445.070 1228.680 ;
        RECT 1444.560 1214.130 1444.700 1219.680 ;
        RECT 1424.720 1213.810 1424.980 1214.130 ;
        RECT 1444.500 1213.810 1444.760 1214.130 ;
        RECT 1352.500 17.010 1352.760 17.330 ;
        RECT 1352.560 2.400 1352.700 17.010 ;
        RECT 1424.780 16.990 1424.920 1213.810 ;
        RECT 1424.720 16.670 1424.980 16.990 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.710 1208.260 1373.030 1208.320 ;
        RECT 1453.670 1208.260 1453.990 1208.320 ;
        RECT 1372.710 1208.120 1453.990 1208.260 ;
        RECT 1372.710 1208.060 1373.030 1208.120 ;
        RECT 1453.670 1208.060 1453.990 1208.120 ;
        RECT 1370.410 20.640 1370.730 20.700 ;
        RECT 1372.710 20.640 1373.030 20.700 ;
        RECT 1370.410 20.500 1373.030 20.640 ;
        RECT 1370.410 20.440 1370.730 20.500 ;
        RECT 1372.710 20.440 1373.030 20.500 ;
      LAYER via ;
        RECT 1372.740 1208.060 1373.000 1208.320 ;
        RECT 1453.700 1208.060 1453.960 1208.320 ;
        RECT 1370.440 20.440 1370.700 20.700 ;
        RECT 1372.740 20.440 1373.000 20.700 ;
      LAYER met2 ;
        RECT 1453.710 1219.680 1454.270 1228.680 ;
        RECT 1453.760 1208.350 1453.900 1219.680 ;
        RECT 1372.740 1208.030 1373.000 1208.350 ;
        RECT 1453.700 1208.030 1453.960 1208.350 ;
        RECT 1372.800 20.730 1372.940 1208.030 ;
        RECT 1370.440 20.410 1370.700 20.730 ;
        RECT 1372.740 20.410 1373.000 20.730 ;
        RECT 1370.500 2.400 1370.640 20.410 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1431.590 1213.360 1431.910 1213.420 ;
        RECT 1462.870 1213.360 1463.190 1213.420 ;
        RECT 1431.590 1213.220 1463.190 1213.360 ;
        RECT 1431.590 1213.160 1431.910 1213.220 ;
        RECT 1462.870 1213.160 1463.190 1213.220 ;
        RECT 1388.350 17.920 1388.670 17.980 ;
        RECT 1431.590 17.920 1431.910 17.980 ;
        RECT 1388.350 17.780 1431.910 17.920 ;
        RECT 1388.350 17.720 1388.670 17.780 ;
        RECT 1431.590 17.720 1431.910 17.780 ;
      LAYER via ;
        RECT 1431.620 1213.160 1431.880 1213.420 ;
        RECT 1462.900 1213.160 1463.160 1213.420 ;
        RECT 1388.380 17.720 1388.640 17.980 ;
        RECT 1431.620 17.720 1431.880 17.980 ;
      LAYER met2 ;
        RECT 1462.910 1219.680 1463.470 1228.680 ;
        RECT 1462.960 1213.450 1463.100 1219.680 ;
        RECT 1431.620 1213.130 1431.880 1213.450 ;
        RECT 1462.900 1213.130 1463.160 1213.450 ;
        RECT 1431.680 18.010 1431.820 1213.130 ;
        RECT 1388.380 17.690 1388.640 18.010 ;
        RECT 1431.620 17.690 1431.880 18.010 ;
        RECT 1388.440 2.400 1388.580 17.690 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 1211.320 1407.530 1211.380 ;
        RECT 1472.070 1211.320 1472.390 1211.380 ;
        RECT 1407.210 1211.180 1472.390 1211.320 ;
        RECT 1407.210 1211.120 1407.530 1211.180 ;
        RECT 1472.070 1211.120 1472.390 1211.180 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1407.210 2.960 1407.530 3.020 ;
        RECT 1406.290 2.820 1407.530 2.960 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
        RECT 1407.210 2.760 1407.530 2.820 ;
      LAYER via ;
        RECT 1407.240 1211.120 1407.500 1211.380 ;
        RECT 1472.100 1211.120 1472.360 1211.380 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
        RECT 1407.240 2.760 1407.500 3.020 ;
      LAYER met2 ;
        RECT 1472.110 1219.680 1472.670 1228.680 ;
        RECT 1472.160 1211.410 1472.300 1219.680 ;
        RECT 1407.240 1211.090 1407.500 1211.410 ;
        RECT 1472.100 1211.090 1472.360 1211.410 ;
        RECT 1407.300 3.050 1407.440 1211.090 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1407.240 2.730 1407.500 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1452.290 1207.920 1452.610 1207.980 ;
        RECT 1481.270 1207.920 1481.590 1207.980 ;
        RECT 1452.290 1207.780 1481.590 1207.920 ;
        RECT 1452.290 1207.720 1452.610 1207.780 ;
        RECT 1481.270 1207.720 1481.590 1207.780 ;
        RECT 1423.770 16.560 1424.090 16.620 ;
        RECT 1452.290 16.560 1452.610 16.620 ;
        RECT 1423.770 16.420 1452.610 16.560 ;
        RECT 1423.770 16.360 1424.090 16.420 ;
        RECT 1452.290 16.360 1452.610 16.420 ;
      LAYER via ;
        RECT 1452.320 1207.720 1452.580 1207.980 ;
        RECT 1481.300 1207.720 1481.560 1207.980 ;
        RECT 1423.800 16.360 1424.060 16.620 ;
        RECT 1452.320 16.360 1452.580 16.620 ;
      LAYER met2 ;
        RECT 1481.310 1219.680 1481.870 1228.680 ;
        RECT 1481.360 1208.010 1481.500 1219.680 ;
        RECT 1452.320 1207.690 1452.580 1208.010 ;
        RECT 1481.300 1207.690 1481.560 1208.010 ;
        RECT 1452.380 16.650 1452.520 1207.690 ;
        RECT 1423.800 16.330 1424.060 16.650 ;
        RECT 1452.320 16.330 1452.580 16.650 ;
        RECT 1423.860 2.400 1424.000 16.330 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 1212.000 1442.030 1212.060 ;
        RECT 1490.470 1212.000 1490.790 1212.060 ;
        RECT 1441.710 1211.860 1490.790 1212.000 ;
        RECT 1441.710 1211.800 1442.030 1211.860 ;
        RECT 1490.470 1211.800 1490.790 1211.860 ;
      LAYER via ;
        RECT 1441.740 1211.800 1442.000 1212.060 ;
        RECT 1490.500 1211.800 1490.760 1212.060 ;
      LAYER met2 ;
        RECT 1490.510 1219.680 1491.070 1228.680 ;
        RECT 1490.560 1212.090 1490.700 1219.680 ;
        RECT 1441.740 1211.770 1442.000 1212.090 ;
        RECT 1490.500 1211.770 1490.760 1212.090 ;
        RECT 1441.800 2.400 1441.940 1211.770 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1462.410 1212.340 1462.730 1212.400 ;
        RECT 1499.670 1212.340 1499.990 1212.400 ;
        RECT 1462.410 1212.200 1499.990 1212.340 ;
        RECT 1462.410 1212.140 1462.730 1212.200 ;
        RECT 1499.670 1212.140 1499.990 1212.200 ;
        RECT 1459.650 20.640 1459.970 20.700 ;
        RECT 1462.410 20.640 1462.730 20.700 ;
        RECT 1459.650 20.500 1462.730 20.640 ;
        RECT 1459.650 20.440 1459.970 20.500 ;
        RECT 1462.410 20.440 1462.730 20.500 ;
      LAYER via ;
        RECT 1462.440 1212.140 1462.700 1212.400 ;
        RECT 1499.700 1212.140 1499.960 1212.400 ;
        RECT 1459.680 20.440 1459.940 20.700 ;
        RECT 1462.440 20.440 1462.700 20.700 ;
      LAYER met2 ;
        RECT 1499.710 1219.680 1500.270 1228.680 ;
        RECT 1499.760 1212.430 1499.900 1219.680 ;
        RECT 1462.440 1212.110 1462.700 1212.430 ;
        RECT 1499.700 1212.110 1499.960 1212.430 ;
        RECT 1462.500 20.730 1462.640 1212.110 ;
        RECT 1459.680 20.410 1459.940 20.730 ;
        RECT 1462.440 20.410 1462.700 20.730 ;
        RECT 1459.740 2.400 1459.880 20.410 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1493.690 1208.260 1494.010 1208.320 ;
        RECT 1508.870 1208.260 1509.190 1208.320 ;
        RECT 1493.690 1208.120 1509.190 1208.260 ;
        RECT 1493.690 1208.060 1494.010 1208.120 ;
        RECT 1508.870 1208.060 1509.190 1208.120 ;
        RECT 1477.590 20.640 1477.910 20.700 ;
        RECT 1493.690 20.640 1494.010 20.700 ;
        RECT 1477.590 20.500 1494.010 20.640 ;
        RECT 1477.590 20.440 1477.910 20.500 ;
        RECT 1493.690 20.440 1494.010 20.500 ;
      LAYER via ;
        RECT 1493.720 1208.060 1493.980 1208.320 ;
        RECT 1508.900 1208.060 1509.160 1208.320 ;
        RECT 1477.620 20.440 1477.880 20.700 ;
        RECT 1493.720 20.440 1493.980 20.700 ;
      LAYER met2 ;
        RECT 1508.910 1219.680 1509.470 1228.680 ;
        RECT 1508.960 1208.350 1509.100 1219.680 ;
        RECT 1493.720 1208.030 1493.980 1208.350 ;
        RECT 1508.900 1208.030 1509.160 1208.350 ;
        RECT 1493.780 20.730 1493.920 1208.030 ;
        RECT 1477.620 20.410 1477.880 20.730 ;
        RECT 1493.720 20.410 1493.980 20.730 ;
        RECT 1477.680 2.400 1477.820 20.410 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1507.490 1207.920 1507.810 1207.980 ;
        RECT 1518.070 1207.920 1518.390 1207.980 ;
        RECT 1507.490 1207.780 1518.390 1207.920 ;
        RECT 1507.490 1207.720 1507.810 1207.780 ;
        RECT 1518.070 1207.720 1518.390 1207.780 ;
        RECT 1495.530 15.880 1495.850 15.940 ;
        RECT 1507.490 15.880 1507.810 15.940 ;
        RECT 1495.530 15.740 1507.810 15.880 ;
        RECT 1495.530 15.680 1495.850 15.740 ;
        RECT 1507.490 15.680 1507.810 15.740 ;
      LAYER via ;
        RECT 1507.520 1207.720 1507.780 1207.980 ;
        RECT 1518.100 1207.720 1518.360 1207.980 ;
        RECT 1495.560 15.680 1495.820 15.940 ;
        RECT 1507.520 15.680 1507.780 15.940 ;
      LAYER met2 ;
        RECT 1518.110 1219.680 1518.670 1228.680 ;
        RECT 1518.160 1208.010 1518.300 1219.680 ;
        RECT 1507.520 1207.690 1507.780 1208.010 ;
        RECT 1518.100 1207.690 1518.360 1208.010 ;
        RECT 1507.580 15.970 1507.720 1207.690 ;
        RECT 1495.560 15.650 1495.820 15.970 ;
        RECT 1507.520 15.650 1507.780 15.970 ;
        RECT 1495.620 2.400 1495.760 15.650 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1521.290 1207.920 1521.610 1207.980 ;
        RECT 1526.810 1207.920 1527.130 1207.980 ;
        RECT 1521.290 1207.780 1527.130 1207.920 ;
        RECT 1521.290 1207.720 1521.610 1207.780 ;
        RECT 1526.810 1207.720 1527.130 1207.780 ;
        RECT 1513.010 20.300 1513.330 20.360 ;
        RECT 1521.290 20.300 1521.610 20.360 ;
        RECT 1513.010 20.160 1521.610 20.300 ;
        RECT 1513.010 20.100 1513.330 20.160 ;
        RECT 1521.290 20.100 1521.610 20.160 ;
      LAYER via ;
        RECT 1521.320 1207.720 1521.580 1207.980 ;
        RECT 1526.840 1207.720 1527.100 1207.980 ;
        RECT 1513.040 20.100 1513.300 20.360 ;
        RECT 1521.320 20.100 1521.580 20.360 ;
      LAYER met2 ;
        RECT 1526.850 1219.680 1527.410 1228.680 ;
        RECT 1526.900 1208.010 1527.040 1219.680 ;
        RECT 1521.320 1207.690 1521.580 1208.010 ;
        RECT 1526.840 1207.690 1527.100 1208.010 ;
        RECT 1521.380 20.390 1521.520 1207.690 ;
        RECT 1513.040 20.070 1513.300 20.390 ;
        RECT 1521.320 20.070 1521.580 20.390 ;
        RECT 1513.100 2.400 1513.240 20.070 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1112.425 144.925 1112.595 210.375 ;
      LAYER mcon ;
        RECT 1112.425 210.205 1112.595 210.375 ;
      LAYER met1 ;
        RECT 1112.350 1183.440 1112.670 1183.500 ;
        RECT 1113.270 1183.440 1113.590 1183.500 ;
        RECT 1112.350 1183.300 1113.590 1183.440 ;
        RECT 1112.350 1183.240 1112.670 1183.300 ;
        RECT 1113.270 1183.240 1113.590 1183.300 ;
        RECT 1112.810 1077.020 1113.130 1077.080 ;
        RECT 1112.440 1076.880 1113.130 1077.020 ;
        RECT 1112.440 1076.400 1112.580 1076.880 ;
        RECT 1112.810 1076.820 1113.130 1076.880 ;
        RECT 1112.350 1076.140 1112.670 1076.400 ;
        RECT 1112.350 1014.460 1112.670 1014.520 ;
        RECT 1112.810 1014.460 1113.130 1014.520 ;
        RECT 1112.350 1014.320 1113.130 1014.460 ;
        RECT 1112.350 1014.260 1112.670 1014.320 ;
        RECT 1112.810 1014.260 1113.130 1014.320 ;
        RECT 1112.810 1007.320 1113.130 1007.380 ;
        RECT 1113.270 1007.320 1113.590 1007.380 ;
        RECT 1112.810 1007.180 1113.590 1007.320 ;
        RECT 1112.810 1007.120 1113.130 1007.180 ;
        RECT 1113.270 1007.120 1113.590 1007.180 ;
        RECT 1112.350 869.620 1112.670 869.680 ;
        RECT 1113.270 869.620 1113.590 869.680 ;
        RECT 1112.350 869.480 1113.590 869.620 ;
        RECT 1112.350 869.420 1112.670 869.480 ;
        RECT 1113.270 869.420 1113.590 869.480 ;
        RECT 1112.350 772.720 1112.670 772.780 ;
        RECT 1113.270 772.720 1113.590 772.780 ;
        RECT 1112.350 772.580 1113.590 772.720 ;
        RECT 1112.350 772.520 1112.670 772.580 ;
        RECT 1113.270 772.520 1113.590 772.580 ;
        RECT 1112.810 593.680 1113.130 593.940 ;
        RECT 1112.900 593.260 1113.040 593.680 ;
        RECT 1112.810 593.000 1113.130 593.260 ;
        RECT 1112.350 531.320 1112.670 531.380 ;
        RECT 1112.810 531.320 1113.130 531.380 ;
        RECT 1112.350 531.180 1113.130 531.320 ;
        RECT 1112.350 531.120 1112.670 531.180 ;
        RECT 1112.810 531.120 1113.130 531.180 ;
        RECT 1112.350 523.980 1112.670 524.240 ;
        RECT 1112.440 523.840 1112.580 523.980 ;
        RECT 1112.810 523.840 1113.130 523.900 ;
        RECT 1112.440 523.700 1113.130 523.840 ;
        RECT 1112.810 523.640 1113.130 523.700 ;
        RECT 1112.350 434.760 1112.670 434.820 ;
        RECT 1112.810 434.760 1113.130 434.820 ;
        RECT 1112.350 434.620 1113.130 434.760 ;
        RECT 1112.350 434.560 1112.670 434.620 ;
        RECT 1112.810 434.560 1113.130 434.620 ;
        RECT 1112.350 338.200 1112.670 338.260 ;
        RECT 1112.810 338.200 1113.130 338.260 ;
        RECT 1112.350 338.060 1113.130 338.200 ;
        RECT 1112.350 338.000 1112.670 338.060 ;
        RECT 1112.810 338.000 1113.130 338.060 ;
        RECT 1112.350 210.360 1112.670 210.420 ;
        RECT 1112.155 210.220 1112.670 210.360 ;
        RECT 1112.350 210.160 1112.670 210.220 ;
        RECT 1112.365 145.080 1112.655 145.125 ;
        RECT 1113.270 145.080 1113.590 145.140 ;
        RECT 1112.365 144.940 1113.590 145.080 ;
        RECT 1112.365 144.895 1112.655 144.940 ;
        RECT 1113.270 144.880 1113.590 144.940 ;
        RECT 710.310 42.400 710.630 42.460 ;
        RECT 1111.890 42.400 1112.210 42.460 ;
        RECT 710.310 42.260 1112.210 42.400 ;
        RECT 710.310 42.200 710.630 42.260 ;
        RECT 1111.890 42.200 1112.210 42.260 ;
      LAYER via ;
        RECT 1112.380 1183.240 1112.640 1183.500 ;
        RECT 1113.300 1183.240 1113.560 1183.500 ;
        RECT 1112.840 1076.820 1113.100 1077.080 ;
        RECT 1112.380 1076.140 1112.640 1076.400 ;
        RECT 1112.380 1014.260 1112.640 1014.520 ;
        RECT 1112.840 1014.260 1113.100 1014.520 ;
        RECT 1112.840 1007.120 1113.100 1007.380 ;
        RECT 1113.300 1007.120 1113.560 1007.380 ;
        RECT 1112.380 869.420 1112.640 869.680 ;
        RECT 1113.300 869.420 1113.560 869.680 ;
        RECT 1112.380 772.520 1112.640 772.780 ;
        RECT 1113.300 772.520 1113.560 772.780 ;
        RECT 1112.840 593.680 1113.100 593.940 ;
        RECT 1112.840 593.000 1113.100 593.260 ;
        RECT 1112.380 531.120 1112.640 531.380 ;
        RECT 1112.840 531.120 1113.100 531.380 ;
        RECT 1112.380 523.980 1112.640 524.240 ;
        RECT 1112.840 523.640 1113.100 523.900 ;
        RECT 1112.380 434.560 1112.640 434.820 ;
        RECT 1112.840 434.560 1113.100 434.820 ;
        RECT 1112.380 338.000 1112.640 338.260 ;
        RECT 1112.840 338.000 1113.100 338.260 ;
        RECT 1112.380 210.160 1112.640 210.420 ;
        RECT 1113.300 144.880 1113.560 145.140 ;
        RECT 710.340 42.200 710.600 42.460 ;
        RECT 1111.920 42.200 1112.180 42.460 ;
      LAYER met2 ;
        RECT 1114.690 1220.330 1115.250 1228.680 ;
        RECT 1113.360 1220.190 1115.250 1220.330 ;
        RECT 1113.360 1183.530 1113.500 1220.190 ;
        RECT 1114.690 1219.680 1115.250 1220.190 ;
        RECT 1112.380 1183.210 1112.640 1183.530 ;
        RECT 1113.300 1183.210 1113.560 1183.530 ;
        RECT 1112.440 1159.130 1112.580 1183.210 ;
        RECT 1112.440 1158.990 1113.040 1159.130 ;
        RECT 1112.900 1077.110 1113.040 1158.990 ;
        RECT 1112.840 1076.790 1113.100 1077.110 ;
        RECT 1112.380 1076.110 1112.640 1076.430 ;
        RECT 1112.440 1014.550 1112.580 1076.110 ;
        RECT 1112.380 1014.230 1112.640 1014.550 ;
        RECT 1112.840 1014.230 1113.100 1014.550 ;
        RECT 1112.900 1007.410 1113.040 1014.230 ;
        RECT 1112.840 1007.090 1113.100 1007.410 ;
        RECT 1113.300 1007.090 1113.560 1007.410 ;
        RECT 1113.360 869.710 1113.500 1007.090 ;
        RECT 1112.380 869.390 1112.640 869.710 ;
        RECT 1113.300 869.390 1113.560 869.710 ;
        RECT 1112.440 847.010 1112.580 869.390 ;
        RECT 1112.440 846.870 1113.040 847.010 ;
        RECT 1112.900 796.010 1113.040 846.870 ;
        RECT 1112.440 795.870 1113.040 796.010 ;
        RECT 1112.440 772.810 1112.580 795.870 ;
        RECT 1112.380 772.490 1112.640 772.810 ;
        RECT 1113.300 772.490 1113.560 772.810 ;
        RECT 1113.360 676.445 1113.500 772.490 ;
        RECT 1112.370 676.075 1112.650 676.445 ;
        RECT 1113.290 676.075 1113.570 676.445 ;
        RECT 1112.440 628.050 1112.580 676.075 ;
        RECT 1112.440 627.910 1113.040 628.050 ;
        RECT 1112.900 593.970 1113.040 627.910 ;
        RECT 1112.840 593.650 1113.100 593.970 ;
        RECT 1112.840 592.970 1113.100 593.290 ;
        RECT 1112.900 531.410 1113.040 592.970 ;
        RECT 1112.380 531.090 1112.640 531.410 ;
        RECT 1112.840 531.090 1113.100 531.410 ;
        RECT 1112.440 524.270 1112.580 531.090 ;
        RECT 1112.380 523.950 1112.640 524.270 ;
        RECT 1112.840 523.610 1113.100 523.930 ;
        RECT 1112.900 434.850 1113.040 523.610 ;
        RECT 1112.380 434.530 1112.640 434.850 ;
        RECT 1112.840 434.530 1113.100 434.850 ;
        RECT 1112.440 413.850 1112.580 434.530 ;
        RECT 1112.440 413.710 1113.040 413.850 ;
        RECT 1112.900 338.290 1113.040 413.710 ;
        RECT 1112.380 337.970 1112.640 338.290 ;
        RECT 1112.840 337.970 1113.100 338.290 ;
        RECT 1112.440 289.410 1112.580 337.970 ;
        RECT 1111.980 289.270 1112.580 289.410 ;
        RECT 1111.980 241.810 1112.120 289.270 ;
        RECT 1111.980 241.670 1112.580 241.810 ;
        RECT 1112.440 210.450 1112.580 241.670 ;
        RECT 1112.380 210.130 1112.640 210.450 ;
        RECT 1113.300 144.850 1113.560 145.170 ;
        RECT 1113.360 72.490 1113.500 144.850 ;
        RECT 1111.980 72.350 1113.500 72.490 ;
        RECT 1111.980 42.490 1112.120 72.350 ;
        RECT 710.340 42.170 710.600 42.490 ;
        RECT 1111.920 42.170 1112.180 42.490 ;
        RECT 710.400 2.400 710.540 42.170 ;
        RECT 710.190 -4.800 710.750 2.400 ;
      LAYER via2 ;
        RECT 1112.370 676.120 1112.650 676.400 ;
        RECT 1113.290 676.120 1113.570 676.400 ;
      LAYER met3 ;
        RECT 1112.345 676.410 1112.675 676.425 ;
        RECT 1113.265 676.410 1113.595 676.425 ;
        RECT 1112.345 676.110 1113.595 676.410 ;
        RECT 1112.345 676.095 1112.675 676.110 ;
        RECT 1113.265 676.095 1113.595 676.110 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1536.010 1207.580 1536.330 1207.640 ;
        RECT 1531.500 1207.440 1536.330 1207.580 ;
        RECT 1531.500 1207.300 1531.640 1207.440 ;
        RECT 1536.010 1207.380 1536.330 1207.440 ;
        RECT 1531.410 1207.040 1531.730 1207.300 ;
      LAYER via ;
        RECT 1536.040 1207.380 1536.300 1207.640 ;
        RECT 1531.440 1207.040 1531.700 1207.300 ;
      LAYER met2 ;
        RECT 1536.050 1219.680 1536.610 1228.680 ;
        RECT 1536.100 1207.670 1536.240 1219.680 ;
        RECT 1536.040 1207.350 1536.300 1207.670 ;
        RECT 1531.440 1207.010 1531.700 1207.330 ;
        RECT 1531.500 20.130 1531.640 1207.010 ;
        RECT 1531.040 19.990 1531.640 20.130 ;
        RECT 1531.040 2.400 1531.180 19.990 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1547.050 48.520 1547.370 48.580 ;
        RECT 1548.890 48.520 1549.210 48.580 ;
        RECT 1547.050 48.380 1549.210 48.520 ;
        RECT 1547.050 48.320 1547.370 48.380 ;
        RECT 1548.890 48.320 1549.210 48.380 ;
      LAYER via ;
        RECT 1547.080 48.320 1547.340 48.580 ;
        RECT 1548.920 48.320 1549.180 48.580 ;
      LAYER met2 ;
        RECT 1545.250 1219.680 1545.810 1228.680 ;
        RECT 1545.300 1207.920 1545.440 1219.680 ;
        RECT 1545.300 1207.780 1546.820 1207.920 ;
        RECT 1546.680 72.490 1546.820 1207.780 ;
        RECT 1546.680 72.350 1547.280 72.490 ;
        RECT 1547.140 48.610 1547.280 72.350 ;
        RECT 1547.080 48.290 1547.340 48.610 ;
        RECT 1548.920 48.290 1549.180 48.610 ;
        RECT 1548.980 2.400 1549.120 48.290 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1554.410 1207.580 1554.730 1207.640 ;
        RECT 1562.690 1207.580 1563.010 1207.640 ;
        RECT 1554.410 1207.440 1563.010 1207.580 ;
        RECT 1554.410 1207.380 1554.730 1207.440 ;
        RECT 1562.690 1207.380 1563.010 1207.440 ;
        RECT 1562.690 17.580 1563.010 17.640 ;
        RECT 1566.830 17.580 1567.150 17.640 ;
        RECT 1562.690 17.440 1567.150 17.580 ;
        RECT 1562.690 17.380 1563.010 17.440 ;
        RECT 1566.830 17.380 1567.150 17.440 ;
      LAYER via ;
        RECT 1554.440 1207.380 1554.700 1207.640 ;
        RECT 1562.720 1207.380 1562.980 1207.640 ;
        RECT 1562.720 17.380 1562.980 17.640 ;
        RECT 1566.860 17.380 1567.120 17.640 ;
      LAYER met2 ;
        RECT 1554.450 1219.680 1555.010 1228.680 ;
        RECT 1554.500 1207.670 1554.640 1219.680 ;
        RECT 1554.440 1207.350 1554.700 1207.670 ;
        RECT 1562.720 1207.350 1562.980 1207.670 ;
        RECT 1562.780 17.670 1562.920 1207.350 ;
        RECT 1562.720 17.350 1562.980 17.670 ;
        RECT 1566.860 17.350 1567.120 17.670 ;
        RECT 1566.920 2.400 1567.060 17.350 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1563.610 1214.380 1563.930 1214.440 ;
        RECT 1580.170 1214.380 1580.490 1214.440 ;
        RECT 1563.610 1214.240 1580.490 1214.380 ;
        RECT 1563.610 1214.180 1563.930 1214.240 ;
        RECT 1580.170 1214.180 1580.490 1214.240 ;
      LAYER via ;
        RECT 1563.640 1214.180 1563.900 1214.440 ;
        RECT 1580.200 1214.180 1580.460 1214.440 ;
      LAYER met2 ;
        RECT 1563.650 1219.680 1564.210 1228.680 ;
        RECT 1563.700 1214.470 1563.840 1219.680 ;
        RECT 1563.640 1214.150 1563.900 1214.470 ;
        RECT 1580.200 1214.150 1580.460 1214.470 ;
        RECT 1580.260 16.730 1580.400 1214.150 ;
        RECT 1580.260 16.590 1585.000 16.730 ;
        RECT 1584.860 2.400 1585.000 16.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.810 1213.700 1573.130 1213.760 ;
        RECT 1583.850 1213.700 1584.170 1213.760 ;
        RECT 1572.810 1213.560 1584.170 1213.700 ;
        RECT 1572.810 1213.500 1573.130 1213.560 ;
        RECT 1583.850 1213.500 1584.170 1213.560 ;
        RECT 1583.850 18.260 1584.170 18.320 ;
        RECT 1602.250 18.260 1602.570 18.320 ;
        RECT 1583.850 18.120 1602.570 18.260 ;
        RECT 1583.850 18.060 1584.170 18.120 ;
        RECT 1602.250 18.060 1602.570 18.120 ;
      LAYER via ;
        RECT 1572.840 1213.500 1573.100 1213.760 ;
        RECT 1583.880 1213.500 1584.140 1213.760 ;
        RECT 1583.880 18.060 1584.140 18.320 ;
        RECT 1602.280 18.060 1602.540 18.320 ;
      LAYER met2 ;
        RECT 1572.850 1219.680 1573.410 1228.680 ;
        RECT 1572.900 1213.790 1573.040 1219.680 ;
        RECT 1572.840 1213.470 1573.100 1213.790 ;
        RECT 1583.880 1213.470 1584.140 1213.790 ;
        RECT 1583.940 18.350 1584.080 1213.470 ;
        RECT 1583.880 18.030 1584.140 18.350 ;
        RECT 1602.280 18.030 1602.540 18.350 ;
        RECT 1602.340 2.400 1602.480 18.030 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1582.010 1207.920 1582.330 1207.980 ;
        RECT 1604.090 1207.920 1604.410 1207.980 ;
        RECT 1582.010 1207.780 1604.410 1207.920 ;
        RECT 1582.010 1207.720 1582.330 1207.780 ;
        RECT 1604.090 1207.720 1604.410 1207.780 ;
        RECT 1604.090 16.220 1604.410 16.280 ;
        RECT 1620.190 16.220 1620.510 16.280 ;
        RECT 1604.090 16.080 1620.510 16.220 ;
        RECT 1604.090 16.020 1604.410 16.080 ;
        RECT 1620.190 16.020 1620.510 16.080 ;
      LAYER via ;
        RECT 1582.040 1207.720 1582.300 1207.980 ;
        RECT 1604.120 1207.720 1604.380 1207.980 ;
        RECT 1604.120 16.020 1604.380 16.280 ;
        RECT 1620.220 16.020 1620.480 16.280 ;
      LAYER met2 ;
        RECT 1582.050 1219.680 1582.610 1228.680 ;
        RECT 1582.100 1208.010 1582.240 1219.680 ;
        RECT 1582.040 1207.690 1582.300 1208.010 ;
        RECT 1604.120 1207.690 1604.380 1208.010 ;
        RECT 1604.180 16.310 1604.320 1207.690 ;
        RECT 1604.120 15.990 1604.380 16.310 ;
        RECT 1620.220 15.990 1620.480 16.310 ;
        RECT 1620.280 2.400 1620.420 15.990 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1591.210 1210.980 1591.530 1211.040 ;
        RECT 1636.290 1210.980 1636.610 1211.040 ;
        RECT 1591.210 1210.840 1636.610 1210.980 ;
        RECT 1591.210 1210.780 1591.530 1210.840 ;
        RECT 1636.290 1210.780 1636.610 1210.840 ;
      LAYER via ;
        RECT 1591.240 1210.780 1591.500 1211.040 ;
        RECT 1636.320 1210.780 1636.580 1211.040 ;
      LAYER met2 ;
        RECT 1591.250 1219.680 1591.810 1228.680 ;
        RECT 1591.300 1211.070 1591.440 1219.680 ;
        RECT 1591.240 1210.750 1591.500 1211.070 ;
        RECT 1636.320 1210.750 1636.580 1211.070 ;
        RECT 1636.380 3.130 1636.520 1210.750 ;
        RECT 1636.380 2.990 1638.360 3.130 ;
        RECT 1638.220 2.400 1638.360 2.990 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.410 18.940 1600.730 19.000 ;
        RECT 1656.070 18.940 1656.390 19.000 ;
        RECT 1600.410 18.800 1656.390 18.940 ;
        RECT 1600.410 18.740 1600.730 18.800 ;
        RECT 1656.070 18.740 1656.390 18.800 ;
      LAYER via ;
        RECT 1600.440 18.740 1600.700 19.000 ;
        RECT 1656.100 18.740 1656.360 19.000 ;
      LAYER met2 ;
        RECT 1600.450 1219.680 1601.010 1228.680 ;
        RECT 1600.500 19.030 1600.640 1219.680 ;
        RECT 1600.440 18.710 1600.700 19.030 ;
        RECT 1656.100 18.710 1656.360 19.030 ;
        RECT 1656.160 2.400 1656.300 18.710 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1609.610 1207.580 1609.930 1207.640 ;
        RECT 1614.210 1207.580 1614.530 1207.640 ;
        RECT 1609.610 1207.440 1614.530 1207.580 ;
        RECT 1609.610 1207.380 1609.930 1207.440 ;
        RECT 1614.210 1207.380 1614.530 1207.440 ;
        RECT 1614.670 16.900 1614.990 16.960 ;
        RECT 1673.550 16.900 1673.870 16.960 ;
        RECT 1614.670 16.760 1673.870 16.900 ;
        RECT 1614.670 16.700 1614.990 16.760 ;
        RECT 1673.550 16.700 1673.870 16.760 ;
      LAYER via ;
        RECT 1609.640 1207.380 1609.900 1207.640 ;
        RECT 1614.240 1207.380 1614.500 1207.640 ;
        RECT 1614.700 16.700 1614.960 16.960 ;
        RECT 1673.580 16.700 1673.840 16.960 ;
      LAYER met2 ;
        RECT 1609.650 1219.680 1610.210 1228.680 ;
        RECT 1609.700 1207.670 1609.840 1219.680 ;
        RECT 1609.640 1207.350 1609.900 1207.670 ;
        RECT 1614.240 1207.350 1614.500 1207.670 ;
        RECT 1614.300 18.090 1614.440 1207.350 ;
        RECT 1614.300 17.950 1614.900 18.090 ;
        RECT 1614.760 16.990 1614.900 17.950 ;
        RECT 1614.700 16.670 1614.960 16.990 ;
        RECT 1673.580 16.670 1673.840 16.990 ;
        RECT 1673.640 2.400 1673.780 16.670 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1621.110 17.920 1621.430 17.980 ;
        RECT 1691.490 17.920 1691.810 17.980 ;
        RECT 1621.110 17.780 1691.810 17.920 ;
        RECT 1621.110 17.720 1621.430 17.780 ;
        RECT 1691.490 17.720 1691.810 17.780 ;
      LAYER via ;
        RECT 1621.140 17.720 1621.400 17.980 ;
        RECT 1691.520 17.720 1691.780 17.980 ;
      LAYER met2 ;
        RECT 1618.850 1220.330 1619.410 1228.680 ;
        RECT 1618.850 1220.190 1621.340 1220.330 ;
        RECT 1618.850 1219.680 1619.410 1220.190 ;
        RECT 1621.200 18.010 1621.340 1220.190 ;
        RECT 1621.140 17.690 1621.400 18.010 ;
        RECT 1691.520 17.690 1691.780 18.010 ;
        RECT 1691.580 2.400 1691.720 17.690 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1119.325 1104.065 1119.495 1111.035 ;
        RECT 1118.865 476.085 1119.035 524.195 ;
        RECT 1118.865 372.725 1119.035 427.635 ;
        RECT 1118.405 276.165 1118.575 324.275 ;
        RECT 1118.865 144.925 1119.035 210.375 ;
        RECT 1118.405 48.365 1118.575 137.955 ;
      LAYER mcon ;
        RECT 1119.325 1110.865 1119.495 1111.035 ;
        RECT 1118.865 524.025 1119.035 524.195 ;
        RECT 1118.865 427.465 1119.035 427.635 ;
        RECT 1118.405 324.105 1118.575 324.275 ;
        RECT 1118.865 210.205 1119.035 210.375 ;
        RECT 1118.405 137.785 1118.575 137.955 ;
      LAYER met1 ;
        RECT 1118.790 1183.440 1119.110 1183.500 ;
        RECT 1122.010 1183.440 1122.330 1183.500 ;
        RECT 1118.790 1183.300 1122.330 1183.440 ;
        RECT 1118.790 1183.240 1119.110 1183.300 ;
        RECT 1122.010 1183.240 1122.330 1183.300 ;
        RECT 1119.250 1111.020 1119.570 1111.080 ;
        RECT 1119.055 1110.880 1119.570 1111.020 ;
        RECT 1119.250 1110.820 1119.570 1110.880 ;
        RECT 1119.250 1104.220 1119.570 1104.280 ;
        RECT 1119.055 1104.080 1119.570 1104.220 ;
        RECT 1119.250 1104.020 1119.570 1104.080 ;
        RECT 1119.250 1014.460 1119.570 1014.520 ;
        RECT 1119.710 1014.460 1120.030 1014.520 ;
        RECT 1119.250 1014.320 1120.030 1014.460 ;
        RECT 1119.250 1014.260 1119.570 1014.320 ;
        RECT 1119.710 1014.260 1120.030 1014.320 ;
        RECT 1119.250 980.460 1119.570 980.520 ;
        RECT 1118.880 980.320 1119.570 980.460 ;
        RECT 1118.880 979.840 1119.020 980.320 ;
        RECT 1119.250 980.260 1119.570 980.320 ;
        RECT 1118.790 979.580 1119.110 979.840 ;
        RECT 1118.790 959.040 1119.110 959.100 ;
        RECT 1120.170 959.040 1120.490 959.100 ;
        RECT 1118.790 958.900 1120.490 959.040 ;
        RECT 1118.790 958.840 1119.110 958.900 ;
        RECT 1120.170 958.840 1120.490 958.900 ;
        RECT 1118.790 772.720 1119.110 772.780 ;
        RECT 1119.710 772.720 1120.030 772.780 ;
        RECT 1118.790 772.580 1120.030 772.720 ;
        RECT 1118.790 772.520 1119.110 772.580 ;
        RECT 1119.710 772.520 1120.030 772.580 ;
        RECT 1119.250 593.680 1119.570 593.940 ;
        RECT 1119.340 593.260 1119.480 593.680 ;
        RECT 1119.250 593.000 1119.570 593.260 ;
        RECT 1118.790 531.320 1119.110 531.380 ;
        RECT 1119.250 531.320 1119.570 531.380 ;
        RECT 1118.790 531.180 1119.570 531.320 ;
        RECT 1118.790 531.120 1119.110 531.180 ;
        RECT 1119.250 531.120 1119.570 531.180 ;
        RECT 1118.790 524.180 1119.110 524.240 ;
        RECT 1118.595 524.040 1119.110 524.180 ;
        RECT 1118.790 523.980 1119.110 524.040 ;
        RECT 1118.805 476.240 1119.095 476.285 ;
        RECT 1120.170 476.240 1120.490 476.300 ;
        RECT 1118.805 476.100 1120.490 476.240 ;
        RECT 1118.805 476.055 1119.095 476.100 ;
        RECT 1120.170 476.040 1120.490 476.100 ;
        RECT 1118.790 434.760 1119.110 434.820 ;
        RECT 1119.250 434.760 1119.570 434.820 ;
        RECT 1118.790 434.620 1119.570 434.760 ;
        RECT 1118.790 434.560 1119.110 434.620 ;
        RECT 1119.250 434.560 1119.570 434.620 ;
        RECT 1118.790 427.620 1119.110 427.680 ;
        RECT 1118.595 427.480 1119.110 427.620 ;
        RECT 1118.790 427.420 1119.110 427.480 ;
        RECT 1118.790 372.880 1119.110 372.940 ;
        RECT 1118.595 372.740 1119.110 372.880 ;
        RECT 1118.790 372.680 1119.110 372.740 ;
        RECT 1118.345 324.260 1118.635 324.305 ;
        RECT 1118.790 324.260 1119.110 324.320 ;
        RECT 1118.345 324.120 1119.110 324.260 ;
        RECT 1118.345 324.075 1118.635 324.120 ;
        RECT 1118.790 324.060 1119.110 324.120 ;
        RECT 1118.330 276.320 1118.650 276.380 ;
        RECT 1118.135 276.180 1118.650 276.320 ;
        RECT 1118.330 276.120 1118.650 276.180 ;
        RECT 1118.790 210.360 1119.110 210.420 ;
        RECT 1118.595 210.220 1119.110 210.360 ;
        RECT 1118.790 210.160 1119.110 210.220 ;
        RECT 1118.790 145.080 1119.110 145.140 ;
        RECT 1118.595 144.940 1119.110 145.080 ;
        RECT 1118.790 144.880 1119.110 144.940 ;
        RECT 1118.345 137.940 1118.635 137.985 ;
        RECT 1118.790 137.940 1119.110 138.000 ;
        RECT 1118.345 137.800 1119.110 137.940 ;
        RECT 1118.345 137.755 1118.635 137.800 ;
        RECT 1118.790 137.740 1119.110 137.800 ;
        RECT 1118.330 48.520 1118.650 48.580 ;
        RECT 1118.135 48.380 1118.650 48.520 ;
        RECT 1118.330 48.320 1118.650 48.380 ;
        RECT 728.250 42.060 728.570 42.120 ;
        RECT 1118.330 42.060 1118.650 42.120 ;
        RECT 728.250 41.920 1118.650 42.060 ;
        RECT 728.250 41.860 728.570 41.920 ;
        RECT 1118.330 41.860 1118.650 41.920 ;
      LAYER via ;
        RECT 1118.820 1183.240 1119.080 1183.500 ;
        RECT 1122.040 1183.240 1122.300 1183.500 ;
        RECT 1119.280 1110.820 1119.540 1111.080 ;
        RECT 1119.280 1104.020 1119.540 1104.280 ;
        RECT 1119.280 1014.260 1119.540 1014.520 ;
        RECT 1119.740 1014.260 1120.000 1014.520 ;
        RECT 1119.280 980.260 1119.540 980.520 ;
        RECT 1118.820 979.580 1119.080 979.840 ;
        RECT 1118.820 958.840 1119.080 959.100 ;
        RECT 1120.200 958.840 1120.460 959.100 ;
        RECT 1118.820 772.520 1119.080 772.780 ;
        RECT 1119.740 772.520 1120.000 772.780 ;
        RECT 1119.280 593.680 1119.540 593.940 ;
        RECT 1119.280 593.000 1119.540 593.260 ;
        RECT 1118.820 531.120 1119.080 531.380 ;
        RECT 1119.280 531.120 1119.540 531.380 ;
        RECT 1118.820 523.980 1119.080 524.240 ;
        RECT 1120.200 476.040 1120.460 476.300 ;
        RECT 1118.820 434.560 1119.080 434.820 ;
        RECT 1119.280 434.560 1119.540 434.820 ;
        RECT 1118.820 427.420 1119.080 427.680 ;
        RECT 1118.820 372.680 1119.080 372.940 ;
        RECT 1118.820 324.060 1119.080 324.320 ;
        RECT 1118.360 276.120 1118.620 276.380 ;
        RECT 1118.820 210.160 1119.080 210.420 ;
        RECT 1118.820 144.880 1119.080 145.140 ;
        RECT 1118.820 137.740 1119.080 138.000 ;
        RECT 1118.360 48.320 1118.620 48.580 ;
        RECT 728.280 41.860 728.540 42.120 ;
        RECT 1118.360 41.860 1118.620 42.120 ;
      LAYER met2 ;
        RECT 1123.890 1220.330 1124.450 1228.680 ;
        RECT 1122.100 1220.190 1124.450 1220.330 ;
        RECT 1122.100 1183.530 1122.240 1220.190 ;
        RECT 1123.890 1219.680 1124.450 1220.190 ;
        RECT 1118.820 1183.210 1119.080 1183.530 ;
        RECT 1122.040 1183.210 1122.300 1183.530 ;
        RECT 1118.880 1159.245 1119.020 1183.210 ;
        RECT 1118.810 1158.875 1119.090 1159.245 ;
        RECT 1119.730 1158.875 1120.010 1159.245 ;
        RECT 1119.800 1152.330 1119.940 1158.875 ;
        RECT 1119.340 1152.190 1119.940 1152.330 ;
        RECT 1119.340 1111.110 1119.480 1152.190 ;
        RECT 1119.280 1110.790 1119.540 1111.110 ;
        RECT 1119.340 1104.310 1119.480 1104.465 ;
        RECT 1119.280 1104.050 1119.540 1104.310 ;
        RECT 1118.880 1103.990 1119.540 1104.050 ;
        RECT 1118.880 1103.910 1119.480 1103.990 ;
        RECT 1118.880 1055.885 1119.020 1103.910 ;
        RECT 1118.810 1055.515 1119.090 1055.885 ;
        RECT 1119.730 1055.515 1120.010 1055.885 ;
        RECT 1119.800 1014.550 1119.940 1055.515 ;
        RECT 1119.280 1014.230 1119.540 1014.550 ;
        RECT 1119.740 1014.230 1120.000 1014.550 ;
        RECT 1119.340 980.550 1119.480 1014.230 ;
        RECT 1119.280 980.230 1119.540 980.550 ;
        RECT 1118.820 979.550 1119.080 979.870 ;
        RECT 1118.880 959.130 1119.020 979.550 ;
        RECT 1118.820 958.810 1119.080 959.130 ;
        RECT 1120.200 958.810 1120.460 959.130 ;
        RECT 1120.260 911.045 1120.400 958.810 ;
        RECT 1119.270 910.675 1119.550 911.045 ;
        RECT 1120.190 910.675 1120.470 911.045 ;
        RECT 1119.340 784.450 1119.480 910.675 ;
        RECT 1118.880 784.310 1119.480 784.450 ;
        RECT 1118.880 772.810 1119.020 784.310 ;
        RECT 1118.820 772.490 1119.080 772.810 ;
        RECT 1119.740 772.490 1120.000 772.810 ;
        RECT 1119.800 676.445 1119.940 772.490 ;
        RECT 1118.810 676.075 1119.090 676.445 ;
        RECT 1119.730 676.075 1120.010 676.445 ;
        RECT 1118.880 628.050 1119.020 676.075 ;
        RECT 1118.880 627.910 1119.480 628.050 ;
        RECT 1119.340 593.970 1119.480 627.910 ;
        RECT 1119.280 593.650 1119.540 593.970 ;
        RECT 1119.280 592.970 1119.540 593.290 ;
        RECT 1119.340 531.410 1119.480 592.970 ;
        RECT 1118.820 531.090 1119.080 531.410 ;
        RECT 1119.280 531.090 1119.540 531.410 ;
        RECT 1118.880 524.270 1119.020 531.090 ;
        RECT 1118.820 523.950 1119.080 524.270 ;
        RECT 1120.200 476.010 1120.460 476.330 ;
        RECT 1120.260 435.725 1120.400 476.010 ;
        RECT 1120.190 435.355 1120.470 435.725 ;
        RECT 1118.820 434.530 1119.080 434.850 ;
        RECT 1119.270 434.675 1119.550 435.045 ;
        RECT 1119.280 434.530 1119.540 434.675 ;
        RECT 1118.880 427.710 1119.020 434.530 ;
        RECT 1118.820 427.390 1119.080 427.710 ;
        RECT 1118.820 372.650 1119.080 372.970 ;
        RECT 1118.880 324.350 1119.020 372.650 ;
        RECT 1118.820 324.030 1119.080 324.350 ;
        RECT 1118.360 276.090 1118.620 276.410 ;
        RECT 1118.420 241.810 1118.560 276.090 ;
        RECT 1118.420 241.670 1119.020 241.810 ;
        RECT 1118.880 210.450 1119.020 241.670 ;
        RECT 1118.820 210.130 1119.080 210.450 ;
        RECT 1118.820 144.850 1119.080 145.170 ;
        RECT 1118.880 138.030 1119.020 144.850 ;
        RECT 1118.820 137.710 1119.080 138.030 ;
        RECT 1118.360 48.290 1118.620 48.610 ;
        RECT 1118.420 42.150 1118.560 48.290 ;
        RECT 728.280 41.830 728.540 42.150 ;
        RECT 1118.360 41.830 1118.620 42.150 ;
        RECT 728.340 2.400 728.480 41.830 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 1118.810 1158.920 1119.090 1159.200 ;
        RECT 1119.730 1158.920 1120.010 1159.200 ;
        RECT 1118.810 1055.560 1119.090 1055.840 ;
        RECT 1119.730 1055.560 1120.010 1055.840 ;
        RECT 1119.270 910.720 1119.550 911.000 ;
        RECT 1120.190 910.720 1120.470 911.000 ;
        RECT 1118.810 676.120 1119.090 676.400 ;
        RECT 1119.730 676.120 1120.010 676.400 ;
        RECT 1120.190 435.400 1120.470 435.680 ;
        RECT 1119.270 434.720 1119.550 435.000 ;
      LAYER met3 ;
        RECT 1118.785 1159.210 1119.115 1159.225 ;
        RECT 1119.705 1159.210 1120.035 1159.225 ;
        RECT 1118.785 1158.910 1120.035 1159.210 ;
        RECT 1118.785 1158.895 1119.115 1158.910 ;
        RECT 1119.705 1158.895 1120.035 1158.910 ;
        RECT 1118.785 1055.850 1119.115 1055.865 ;
        RECT 1119.705 1055.850 1120.035 1055.865 ;
        RECT 1118.785 1055.550 1120.035 1055.850 ;
        RECT 1118.785 1055.535 1119.115 1055.550 ;
        RECT 1119.705 1055.535 1120.035 1055.550 ;
        RECT 1119.245 911.010 1119.575 911.025 ;
        RECT 1120.165 911.010 1120.495 911.025 ;
        RECT 1119.245 910.710 1120.495 911.010 ;
        RECT 1119.245 910.695 1119.575 910.710 ;
        RECT 1120.165 910.695 1120.495 910.710 ;
        RECT 1118.785 676.410 1119.115 676.425 ;
        RECT 1119.705 676.410 1120.035 676.425 ;
        RECT 1118.785 676.110 1120.035 676.410 ;
        RECT 1118.785 676.095 1119.115 676.110 ;
        RECT 1119.705 676.095 1120.035 676.110 ;
        RECT 1120.165 435.690 1120.495 435.705 ;
        RECT 1119.030 435.390 1120.495 435.690 ;
        RECT 1119.030 435.025 1119.330 435.390 ;
        RECT 1120.165 435.375 1120.495 435.390 ;
        RECT 1119.030 434.710 1119.575 435.025 ;
        RECT 1119.245 434.695 1119.575 434.710 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.010 1213.020 1628.330 1213.080 ;
        RECT 1693.790 1213.020 1694.110 1213.080 ;
        RECT 1628.010 1212.880 1694.110 1213.020 ;
        RECT 1628.010 1212.820 1628.330 1212.880 ;
        RECT 1693.790 1212.820 1694.110 1212.880 ;
        RECT 1693.790 15.200 1694.110 15.260 ;
        RECT 1709.430 15.200 1709.750 15.260 ;
        RECT 1693.790 15.060 1709.750 15.200 ;
        RECT 1693.790 15.000 1694.110 15.060 ;
        RECT 1709.430 15.000 1709.750 15.060 ;
      LAYER via ;
        RECT 1628.040 1212.820 1628.300 1213.080 ;
        RECT 1693.820 1212.820 1694.080 1213.080 ;
        RECT 1693.820 15.000 1694.080 15.260 ;
        RECT 1709.460 15.000 1709.720 15.260 ;
      LAYER met2 ;
        RECT 1628.050 1219.680 1628.610 1228.680 ;
        RECT 1628.100 1213.110 1628.240 1219.680 ;
        RECT 1628.040 1212.790 1628.300 1213.110 ;
        RECT 1693.820 1212.790 1694.080 1213.110 ;
        RECT 1693.880 15.290 1694.020 1212.790 ;
        RECT 1693.820 14.970 1694.080 15.290 ;
        RECT 1709.460 14.970 1709.720 15.290 ;
        RECT 1709.520 2.400 1709.660 14.970 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1637.210 1207.580 1637.530 1207.640 ;
        RECT 1641.810 1207.580 1642.130 1207.640 ;
        RECT 1637.210 1207.440 1642.130 1207.580 ;
        RECT 1637.210 1207.380 1637.530 1207.440 ;
        RECT 1641.810 1207.380 1642.130 1207.440 ;
        RECT 1641.810 19.960 1642.130 20.020 ;
        RECT 1727.370 19.960 1727.690 20.020 ;
        RECT 1641.810 19.820 1727.690 19.960 ;
        RECT 1641.810 19.760 1642.130 19.820 ;
        RECT 1727.370 19.760 1727.690 19.820 ;
      LAYER via ;
        RECT 1637.240 1207.380 1637.500 1207.640 ;
        RECT 1641.840 1207.380 1642.100 1207.640 ;
        RECT 1641.840 19.760 1642.100 20.020 ;
        RECT 1727.400 19.760 1727.660 20.020 ;
      LAYER met2 ;
        RECT 1637.250 1219.680 1637.810 1228.680 ;
        RECT 1637.300 1207.670 1637.440 1219.680 ;
        RECT 1637.240 1207.350 1637.500 1207.670 ;
        RECT 1641.840 1207.350 1642.100 1207.670 ;
        RECT 1641.900 20.050 1642.040 1207.350 ;
        RECT 1641.840 19.730 1642.100 20.050 ;
        RECT 1727.400 19.730 1727.660 20.050 ;
        RECT 1727.460 2.400 1727.600 19.730 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1713.645 16.745 1713.815 20.315 ;
      LAYER mcon ;
        RECT 1713.645 20.145 1713.815 20.315 ;
      LAYER met1 ;
        RECT 1645.950 1207.920 1646.270 1207.980 ;
        RECT 1666.190 1207.920 1666.510 1207.980 ;
        RECT 1645.950 1207.780 1666.510 1207.920 ;
        RECT 1645.950 1207.720 1646.270 1207.780 ;
        RECT 1666.190 1207.720 1666.510 1207.780 ;
        RECT 1666.190 20.300 1666.510 20.360 ;
        RECT 1713.585 20.300 1713.875 20.345 ;
        RECT 1666.190 20.160 1713.875 20.300 ;
        RECT 1666.190 20.100 1666.510 20.160 ;
        RECT 1713.585 20.115 1713.875 20.160 ;
        RECT 1713.585 16.900 1713.875 16.945 ;
        RECT 1745.310 16.900 1745.630 16.960 ;
        RECT 1713.585 16.760 1745.630 16.900 ;
        RECT 1713.585 16.715 1713.875 16.760 ;
        RECT 1745.310 16.700 1745.630 16.760 ;
      LAYER via ;
        RECT 1645.980 1207.720 1646.240 1207.980 ;
        RECT 1666.220 1207.720 1666.480 1207.980 ;
        RECT 1666.220 20.100 1666.480 20.360 ;
        RECT 1745.340 16.700 1745.600 16.960 ;
      LAYER met2 ;
        RECT 1645.990 1219.680 1646.550 1228.680 ;
        RECT 1646.040 1208.010 1646.180 1219.680 ;
        RECT 1645.980 1207.690 1646.240 1208.010 ;
        RECT 1666.220 1207.690 1666.480 1208.010 ;
        RECT 1666.280 20.390 1666.420 1207.690 ;
        RECT 1666.220 20.070 1666.480 20.390 ;
        RECT 1745.340 16.670 1745.600 16.990 ;
        RECT 1745.400 2.400 1745.540 16.670 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 19.280 1655.930 19.340 ;
        RECT 1762.790 19.280 1763.110 19.340 ;
        RECT 1655.610 19.140 1763.110 19.280 ;
        RECT 1655.610 19.080 1655.930 19.140 ;
        RECT 1762.790 19.080 1763.110 19.140 ;
      LAYER via ;
        RECT 1655.640 19.080 1655.900 19.340 ;
        RECT 1762.820 19.080 1763.080 19.340 ;
      LAYER met2 ;
        RECT 1655.190 1220.330 1655.750 1228.680 ;
        RECT 1655.190 1219.680 1655.840 1220.330 ;
        RECT 1655.700 19.370 1655.840 1219.680 ;
        RECT 1655.640 19.050 1655.900 19.370 ;
        RECT 1762.820 19.050 1763.080 19.370 ;
        RECT 1762.880 2.400 1763.020 19.050 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1664.350 1207.580 1664.670 1207.640 ;
        RECT 1669.410 1207.580 1669.730 1207.640 ;
        RECT 1664.350 1207.440 1669.730 1207.580 ;
        RECT 1664.350 1207.380 1664.670 1207.440 ;
        RECT 1669.410 1207.380 1669.730 1207.440 ;
        RECT 1669.410 18.940 1669.730 19.000 ;
        RECT 1780.730 18.940 1781.050 19.000 ;
        RECT 1669.410 18.800 1781.050 18.940 ;
        RECT 1669.410 18.740 1669.730 18.800 ;
        RECT 1780.730 18.740 1781.050 18.800 ;
      LAYER via ;
        RECT 1664.380 1207.380 1664.640 1207.640 ;
        RECT 1669.440 1207.380 1669.700 1207.640 ;
        RECT 1669.440 18.740 1669.700 19.000 ;
        RECT 1780.760 18.740 1781.020 19.000 ;
      LAYER met2 ;
        RECT 1664.390 1219.680 1664.950 1228.680 ;
        RECT 1664.440 1207.670 1664.580 1219.680 ;
        RECT 1664.380 1207.350 1664.640 1207.670 ;
        RECT 1669.440 1207.350 1669.700 1207.670 ;
        RECT 1669.500 19.030 1669.640 1207.350 ;
        RECT 1669.440 18.710 1669.700 19.030 ;
        RECT 1780.760 18.710 1781.020 19.030 ;
        RECT 1780.820 2.400 1780.960 18.710 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1676.310 18.600 1676.630 18.660 ;
        RECT 1798.670 18.600 1798.990 18.660 ;
        RECT 1676.310 18.460 1798.990 18.600 ;
        RECT 1676.310 18.400 1676.630 18.460 ;
        RECT 1798.670 18.400 1798.990 18.460 ;
      LAYER via ;
        RECT 1676.340 18.400 1676.600 18.660 ;
        RECT 1798.700 18.400 1798.960 18.660 ;
      LAYER met2 ;
        RECT 1673.590 1220.330 1674.150 1228.680 ;
        RECT 1673.590 1220.190 1676.540 1220.330 ;
        RECT 1673.590 1219.680 1674.150 1220.190 ;
        RECT 1676.400 18.690 1676.540 1220.190 ;
        RECT 1676.340 18.370 1676.600 18.690 ;
        RECT 1798.700 18.370 1798.960 18.690 ;
        RECT 1798.760 2.400 1798.900 18.370 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1728.825 18.105 1728.995 20.315 ;
      LAYER mcon ;
        RECT 1728.825 20.145 1728.995 20.315 ;
      LAYER met1 ;
        RECT 1682.750 1207.920 1683.070 1207.980 ;
        RECT 1694.250 1207.920 1694.570 1207.980 ;
        RECT 1682.750 1207.780 1694.570 1207.920 ;
        RECT 1682.750 1207.720 1683.070 1207.780 ;
        RECT 1694.250 1207.720 1694.570 1207.780 ;
        RECT 1694.250 20.640 1694.570 20.700 ;
        RECT 1694.250 20.500 1714.260 20.640 ;
        RECT 1694.250 20.440 1694.570 20.500 ;
        RECT 1714.120 20.300 1714.260 20.500 ;
        RECT 1728.765 20.300 1729.055 20.345 ;
        RECT 1714.120 20.160 1729.055 20.300 ;
        RECT 1728.765 20.115 1729.055 20.160 ;
        RECT 1728.765 18.260 1729.055 18.305 ;
        RECT 1816.610 18.260 1816.930 18.320 ;
        RECT 1728.765 18.120 1816.930 18.260 ;
        RECT 1728.765 18.075 1729.055 18.120 ;
        RECT 1816.610 18.060 1816.930 18.120 ;
      LAYER via ;
        RECT 1682.780 1207.720 1683.040 1207.980 ;
        RECT 1694.280 1207.720 1694.540 1207.980 ;
        RECT 1694.280 20.440 1694.540 20.700 ;
        RECT 1816.640 18.060 1816.900 18.320 ;
      LAYER met2 ;
        RECT 1682.790 1219.680 1683.350 1228.680 ;
        RECT 1682.840 1208.010 1682.980 1219.680 ;
        RECT 1682.780 1207.690 1683.040 1208.010 ;
        RECT 1694.280 1207.690 1694.540 1208.010 ;
        RECT 1694.340 20.730 1694.480 1207.690 ;
        RECT 1694.280 20.410 1694.540 20.730 ;
        RECT 1816.640 18.030 1816.900 18.350 ;
        RECT 1816.700 2.400 1816.840 18.030 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1691.950 1207.580 1692.270 1207.640 ;
        RECT 1697.010 1207.580 1697.330 1207.640 ;
        RECT 1691.950 1207.440 1697.330 1207.580 ;
        RECT 1691.950 1207.380 1692.270 1207.440 ;
        RECT 1697.010 1207.380 1697.330 1207.440 ;
        RECT 1697.010 18.260 1697.330 18.320 ;
        RECT 1697.010 18.120 1728.520 18.260 ;
        RECT 1697.010 18.060 1697.330 18.120 ;
        RECT 1728.380 17.920 1728.520 18.120 ;
        RECT 1834.550 17.920 1834.870 17.980 ;
        RECT 1728.380 17.780 1834.870 17.920 ;
        RECT 1834.550 17.720 1834.870 17.780 ;
      LAYER via ;
        RECT 1691.980 1207.380 1692.240 1207.640 ;
        RECT 1697.040 1207.380 1697.300 1207.640 ;
        RECT 1697.040 18.060 1697.300 18.320 ;
        RECT 1834.580 17.720 1834.840 17.980 ;
      LAYER met2 ;
        RECT 1691.990 1219.680 1692.550 1228.680 ;
        RECT 1692.040 1207.670 1692.180 1219.680 ;
        RECT 1691.980 1207.350 1692.240 1207.670 ;
        RECT 1697.040 1207.350 1697.300 1207.670 ;
        RECT 1697.100 18.350 1697.240 1207.350 ;
        RECT 1697.040 18.030 1697.300 18.350 ;
        RECT 1834.580 17.690 1834.840 18.010 ;
        RECT 1834.640 2.400 1834.780 17.690 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1727.905 15.385 1728.075 17.935 ;
        RECT 1752.285 15.385 1752.455 17.595 ;
      LAYER mcon ;
        RECT 1727.905 17.765 1728.075 17.935 ;
        RECT 1752.285 17.425 1752.455 17.595 ;
      LAYER met1 ;
        RECT 1703.910 17.920 1704.230 17.980 ;
        RECT 1727.845 17.920 1728.135 17.965 ;
        RECT 1703.910 17.780 1728.135 17.920 ;
        RECT 1703.910 17.720 1704.230 17.780 ;
        RECT 1727.845 17.735 1728.135 17.780 ;
        RECT 1752.225 17.580 1752.515 17.625 ;
        RECT 1852.030 17.580 1852.350 17.640 ;
        RECT 1752.225 17.440 1852.350 17.580 ;
        RECT 1752.225 17.395 1752.515 17.440 ;
        RECT 1852.030 17.380 1852.350 17.440 ;
        RECT 1727.845 15.540 1728.135 15.585 ;
        RECT 1752.225 15.540 1752.515 15.585 ;
        RECT 1727.845 15.400 1752.515 15.540 ;
        RECT 1727.845 15.355 1728.135 15.400 ;
        RECT 1752.225 15.355 1752.515 15.400 ;
      LAYER via ;
        RECT 1703.940 17.720 1704.200 17.980 ;
        RECT 1852.060 17.380 1852.320 17.640 ;
      LAYER met2 ;
        RECT 1701.190 1220.330 1701.750 1228.680 ;
        RECT 1701.190 1220.190 1704.140 1220.330 ;
        RECT 1701.190 1219.680 1701.750 1220.190 ;
        RECT 1704.000 18.010 1704.140 1220.190 ;
        RECT 1703.940 17.690 1704.200 18.010 ;
        RECT 1852.060 17.350 1852.320 17.670 ;
        RECT 1852.120 2.400 1852.260 17.350 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1836.005 1213.545 1836.635 1213.715 ;
        RECT 1836.465 1213.205 1836.635 1213.545 ;
        RECT 1871.425 766.105 1871.595 814.215 ;
        RECT 1871.425 669.545 1871.595 717.655 ;
        RECT 1871.425 572.645 1871.595 620.755 ;
        RECT 1871.425 476.085 1871.595 524.195 ;
        RECT 1871.425 379.525 1871.595 427.635 ;
        RECT 1871.425 282.965 1871.595 331.075 ;
        RECT 1871.425 186.405 1871.595 234.515 ;
        RECT 1871.425 89.845 1871.595 137.955 ;
        RECT 1870.965 48.365 1871.135 62.815 ;
        RECT 1870.045 2.805 1870.215 13.515 ;
      LAYER mcon ;
        RECT 1871.425 814.045 1871.595 814.215 ;
        RECT 1871.425 717.485 1871.595 717.655 ;
        RECT 1871.425 620.585 1871.595 620.755 ;
        RECT 1871.425 524.025 1871.595 524.195 ;
        RECT 1871.425 427.465 1871.595 427.635 ;
        RECT 1871.425 330.905 1871.595 331.075 ;
        RECT 1871.425 234.345 1871.595 234.515 ;
        RECT 1871.425 137.785 1871.595 137.955 ;
        RECT 1870.965 62.645 1871.135 62.815 ;
        RECT 1870.045 13.345 1870.215 13.515 ;
      LAYER met1 ;
        RECT 1835.945 1213.700 1836.235 1213.745 ;
        RECT 1752.300 1213.560 1836.235 1213.700 ;
        RECT 1710.350 1213.360 1710.670 1213.420 ;
        RECT 1752.300 1213.360 1752.440 1213.560 ;
        RECT 1835.945 1213.515 1836.235 1213.560 ;
        RECT 1710.350 1213.220 1752.440 1213.360 ;
        RECT 1836.405 1213.360 1836.695 1213.405 ;
        RECT 1838.230 1213.360 1838.550 1213.420 ;
        RECT 1836.405 1213.220 1838.550 1213.360 ;
        RECT 1710.350 1213.160 1710.670 1213.220 ;
        RECT 1836.405 1213.175 1836.695 1213.220 ;
        RECT 1838.230 1213.160 1838.550 1213.220 ;
        RECT 1871.350 1152.500 1871.670 1152.560 ;
        RECT 1872.270 1152.500 1872.590 1152.560 ;
        RECT 1871.350 1152.360 1872.590 1152.500 ;
        RECT 1871.350 1152.300 1871.670 1152.360 ;
        RECT 1872.270 1152.300 1872.590 1152.360 ;
        RECT 1871.350 1007.320 1871.670 1007.380 ;
        RECT 1872.270 1007.320 1872.590 1007.380 ;
        RECT 1871.350 1007.180 1872.590 1007.320 ;
        RECT 1871.350 1007.120 1871.670 1007.180 ;
        RECT 1872.270 1007.120 1872.590 1007.180 ;
        RECT 1871.350 910.760 1871.670 910.820 ;
        RECT 1872.270 910.760 1872.590 910.820 ;
        RECT 1871.350 910.620 1872.590 910.760 ;
        RECT 1871.350 910.560 1871.670 910.620 ;
        RECT 1872.270 910.560 1872.590 910.620 ;
        RECT 1871.350 814.200 1871.670 814.260 ;
        RECT 1871.155 814.060 1871.670 814.200 ;
        RECT 1871.350 814.000 1871.670 814.060 ;
        RECT 1871.350 766.260 1871.670 766.320 ;
        RECT 1871.155 766.120 1871.670 766.260 ;
        RECT 1871.350 766.060 1871.670 766.120 ;
        RECT 1871.350 717.640 1871.670 717.700 ;
        RECT 1871.155 717.500 1871.670 717.640 ;
        RECT 1871.350 717.440 1871.670 717.500 ;
        RECT 1871.350 669.700 1871.670 669.760 ;
        RECT 1871.155 669.560 1871.670 669.700 ;
        RECT 1871.350 669.500 1871.670 669.560 ;
        RECT 1871.350 620.740 1871.670 620.800 ;
        RECT 1871.155 620.600 1871.670 620.740 ;
        RECT 1871.350 620.540 1871.670 620.600 ;
        RECT 1871.350 572.800 1871.670 572.860 ;
        RECT 1871.155 572.660 1871.670 572.800 ;
        RECT 1871.350 572.600 1871.670 572.660 ;
        RECT 1871.350 524.180 1871.670 524.240 ;
        RECT 1871.155 524.040 1871.670 524.180 ;
        RECT 1871.350 523.980 1871.670 524.040 ;
        RECT 1871.350 476.240 1871.670 476.300 ;
        RECT 1871.155 476.100 1871.670 476.240 ;
        RECT 1871.350 476.040 1871.670 476.100 ;
        RECT 1871.350 427.620 1871.670 427.680 ;
        RECT 1871.155 427.480 1871.670 427.620 ;
        RECT 1871.350 427.420 1871.670 427.480 ;
        RECT 1871.350 379.680 1871.670 379.740 ;
        RECT 1871.155 379.540 1871.670 379.680 ;
        RECT 1871.350 379.480 1871.670 379.540 ;
        RECT 1871.350 331.060 1871.670 331.120 ;
        RECT 1871.155 330.920 1871.670 331.060 ;
        RECT 1871.350 330.860 1871.670 330.920 ;
        RECT 1871.350 283.120 1871.670 283.180 ;
        RECT 1871.155 282.980 1871.670 283.120 ;
        RECT 1871.350 282.920 1871.670 282.980 ;
        RECT 1871.350 234.500 1871.670 234.560 ;
        RECT 1871.155 234.360 1871.670 234.500 ;
        RECT 1871.350 234.300 1871.670 234.360 ;
        RECT 1871.350 186.560 1871.670 186.620 ;
        RECT 1871.155 186.420 1871.670 186.560 ;
        RECT 1871.350 186.360 1871.670 186.420 ;
        RECT 1871.350 137.940 1871.670 138.000 ;
        RECT 1871.155 137.800 1871.670 137.940 ;
        RECT 1871.350 137.740 1871.670 137.800 ;
        RECT 1871.350 90.000 1871.670 90.060 ;
        RECT 1871.155 89.860 1871.670 90.000 ;
        RECT 1871.350 89.800 1871.670 89.860 ;
        RECT 1870.905 62.800 1871.195 62.845 ;
        RECT 1871.350 62.800 1871.670 62.860 ;
        RECT 1870.905 62.660 1871.670 62.800 ;
        RECT 1870.905 62.615 1871.195 62.660 ;
        RECT 1871.350 62.600 1871.670 62.660 ;
        RECT 1870.890 48.520 1871.210 48.580 ;
        RECT 1870.695 48.380 1871.210 48.520 ;
        RECT 1870.890 48.320 1871.210 48.380 ;
        RECT 1869.985 13.500 1870.275 13.545 ;
        RECT 1871.350 13.500 1871.670 13.560 ;
        RECT 1869.985 13.360 1871.670 13.500 ;
        RECT 1869.985 13.315 1870.275 13.360 ;
        RECT 1871.350 13.300 1871.670 13.360 ;
        RECT 1869.970 2.960 1870.290 3.020 ;
        RECT 1869.775 2.820 1870.290 2.960 ;
        RECT 1869.970 2.760 1870.290 2.820 ;
      LAYER via ;
        RECT 1710.380 1213.160 1710.640 1213.420 ;
        RECT 1838.260 1213.160 1838.520 1213.420 ;
        RECT 1871.380 1152.300 1871.640 1152.560 ;
        RECT 1872.300 1152.300 1872.560 1152.560 ;
        RECT 1871.380 1007.120 1871.640 1007.380 ;
        RECT 1872.300 1007.120 1872.560 1007.380 ;
        RECT 1871.380 910.560 1871.640 910.820 ;
        RECT 1872.300 910.560 1872.560 910.820 ;
        RECT 1871.380 814.000 1871.640 814.260 ;
        RECT 1871.380 766.060 1871.640 766.320 ;
        RECT 1871.380 717.440 1871.640 717.700 ;
        RECT 1871.380 669.500 1871.640 669.760 ;
        RECT 1871.380 620.540 1871.640 620.800 ;
        RECT 1871.380 572.600 1871.640 572.860 ;
        RECT 1871.380 523.980 1871.640 524.240 ;
        RECT 1871.380 476.040 1871.640 476.300 ;
        RECT 1871.380 427.420 1871.640 427.680 ;
        RECT 1871.380 379.480 1871.640 379.740 ;
        RECT 1871.380 330.860 1871.640 331.120 ;
        RECT 1871.380 282.920 1871.640 283.180 ;
        RECT 1871.380 234.300 1871.640 234.560 ;
        RECT 1871.380 186.360 1871.640 186.620 ;
        RECT 1871.380 137.740 1871.640 138.000 ;
        RECT 1871.380 89.800 1871.640 90.060 ;
        RECT 1871.380 62.600 1871.640 62.860 ;
        RECT 1870.920 48.320 1871.180 48.580 ;
        RECT 1871.380 13.300 1871.640 13.560 ;
        RECT 1870.000 2.760 1870.260 3.020 ;
      LAYER met2 ;
        RECT 1710.390 1219.680 1710.950 1228.680 ;
        RECT 1710.440 1213.450 1710.580 1219.680 ;
        RECT 1710.380 1213.130 1710.640 1213.450 ;
        RECT 1838.260 1213.130 1838.520 1213.450 ;
        RECT 1838.320 1208.885 1838.460 1213.130 ;
        RECT 1838.250 1208.515 1838.530 1208.885 ;
        RECT 1871.370 1207.325 1871.650 1207.695 ;
        RECT 1871.440 1200.725 1871.580 1207.325 ;
        RECT 1871.370 1200.355 1871.650 1200.725 ;
        RECT 1872.290 1200.355 1872.570 1200.725 ;
        RECT 1872.360 1152.590 1872.500 1200.355 ;
        RECT 1871.380 1152.270 1871.640 1152.590 ;
        RECT 1872.300 1152.270 1872.560 1152.590 ;
        RECT 1871.440 1104.165 1871.580 1152.270 ;
        RECT 1871.370 1103.795 1871.650 1104.165 ;
        RECT 1872.290 1103.795 1872.570 1104.165 ;
        RECT 1872.360 1055.885 1872.500 1103.795 ;
        RECT 1871.370 1055.515 1871.650 1055.885 ;
        RECT 1872.290 1055.515 1872.570 1055.885 ;
        RECT 1871.440 1007.410 1871.580 1055.515 ;
        RECT 1871.380 1007.090 1871.640 1007.410 ;
        RECT 1872.300 1007.090 1872.560 1007.410 ;
        RECT 1872.360 959.325 1872.500 1007.090 ;
        RECT 1871.370 958.955 1871.650 959.325 ;
        RECT 1872.290 958.955 1872.570 959.325 ;
        RECT 1871.440 910.850 1871.580 958.955 ;
        RECT 1871.380 910.530 1871.640 910.850 ;
        RECT 1872.300 910.530 1872.560 910.850 ;
        RECT 1872.360 862.765 1872.500 910.530 ;
        RECT 1871.370 862.395 1871.650 862.765 ;
        RECT 1872.290 862.395 1872.570 862.765 ;
        RECT 1871.440 814.290 1871.580 862.395 ;
        RECT 1871.380 813.970 1871.640 814.290 ;
        RECT 1871.380 766.030 1871.640 766.350 ;
        RECT 1871.440 717.730 1871.580 766.030 ;
        RECT 1871.380 717.410 1871.640 717.730 ;
        RECT 1871.380 669.470 1871.640 669.790 ;
        RECT 1871.440 620.830 1871.580 669.470 ;
        RECT 1871.380 620.510 1871.640 620.830 ;
        RECT 1871.380 572.570 1871.640 572.890 ;
        RECT 1871.440 524.270 1871.580 572.570 ;
        RECT 1871.380 523.950 1871.640 524.270 ;
        RECT 1871.380 476.010 1871.640 476.330 ;
        RECT 1871.440 427.710 1871.580 476.010 ;
        RECT 1871.380 427.390 1871.640 427.710 ;
        RECT 1871.380 379.450 1871.640 379.770 ;
        RECT 1871.440 331.150 1871.580 379.450 ;
        RECT 1871.380 330.830 1871.640 331.150 ;
        RECT 1871.380 282.890 1871.640 283.210 ;
        RECT 1871.440 234.590 1871.580 282.890 ;
        RECT 1871.380 234.270 1871.640 234.590 ;
        RECT 1871.380 186.330 1871.640 186.650 ;
        RECT 1871.440 138.030 1871.580 186.330 ;
        RECT 1871.380 137.710 1871.640 138.030 ;
        RECT 1871.380 89.770 1871.640 90.090 ;
        RECT 1871.440 62.890 1871.580 89.770 ;
        RECT 1871.380 62.570 1871.640 62.890 ;
        RECT 1870.920 48.290 1871.180 48.610 ;
        RECT 1870.980 48.010 1871.120 48.290 ;
        RECT 1870.980 47.870 1871.580 48.010 ;
        RECT 1871.440 13.590 1871.580 47.870 ;
        RECT 1871.380 13.270 1871.640 13.590 ;
        RECT 1870.000 2.730 1870.260 3.050 ;
        RECT 1870.060 2.400 1870.200 2.730 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
      LAYER via2 ;
        RECT 1838.250 1208.560 1838.530 1208.840 ;
        RECT 1871.370 1207.370 1871.650 1207.650 ;
        RECT 1871.370 1200.400 1871.650 1200.680 ;
        RECT 1872.290 1200.400 1872.570 1200.680 ;
        RECT 1871.370 1103.840 1871.650 1104.120 ;
        RECT 1872.290 1103.840 1872.570 1104.120 ;
        RECT 1871.370 1055.560 1871.650 1055.840 ;
        RECT 1872.290 1055.560 1872.570 1055.840 ;
        RECT 1871.370 959.000 1871.650 959.280 ;
        RECT 1872.290 959.000 1872.570 959.280 ;
        RECT 1871.370 862.440 1871.650 862.720 ;
        RECT 1872.290 862.440 1872.570 862.720 ;
      LAYER met3 ;
        RECT 1838.225 1208.850 1838.555 1208.865 ;
        RECT 1838.225 1208.550 1870.970 1208.850 ;
        RECT 1838.225 1208.535 1838.555 1208.550 ;
        RECT 1870.670 1207.660 1870.970 1208.550 ;
        RECT 1871.345 1207.660 1871.675 1207.675 ;
        RECT 1870.670 1207.360 1871.675 1207.660 ;
        RECT 1871.345 1207.345 1871.675 1207.360 ;
        RECT 1871.345 1200.690 1871.675 1200.705 ;
        RECT 1872.265 1200.690 1872.595 1200.705 ;
        RECT 1871.345 1200.390 1872.595 1200.690 ;
        RECT 1871.345 1200.375 1871.675 1200.390 ;
        RECT 1872.265 1200.375 1872.595 1200.390 ;
        RECT 1871.345 1104.130 1871.675 1104.145 ;
        RECT 1872.265 1104.130 1872.595 1104.145 ;
        RECT 1871.345 1103.830 1872.595 1104.130 ;
        RECT 1871.345 1103.815 1871.675 1103.830 ;
        RECT 1872.265 1103.815 1872.595 1103.830 ;
        RECT 1871.345 1055.850 1871.675 1055.865 ;
        RECT 1872.265 1055.850 1872.595 1055.865 ;
        RECT 1871.345 1055.550 1872.595 1055.850 ;
        RECT 1871.345 1055.535 1871.675 1055.550 ;
        RECT 1872.265 1055.535 1872.595 1055.550 ;
        RECT 1871.345 959.290 1871.675 959.305 ;
        RECT 1872.265 959.290 1872.595 959.305 ;
        RECT 1871.345 958.990 1872.595 959.290 ;
        RECT 1871.345 958.975 1871.675 958.990 ;
        RECT 1872.265 958.975 1872.595 958.990 ;
        RECT 1871.345 862.730 1871.675 862.745 ;
        RECT 1872.265 862.730 1872.595 862.745 ;
        RECT 1871.345 862.430 1872.595 862.730 ;
        RECT 1871.345 862.415 1871.675 862.430 ;
        RECT 1872.265 862.415 1872.595 862.430 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 746.190 24.380 746.510 24.440 ;
        RECT 1131.670 24.380 1131.990 24.440 ;
        RECT 746.190 24.240 1131.990 24.380 ;
        RECT 746.190 24.180 746.510 24.240 ;
        RECT 1131.670 24.180 1131.990 24.240 ;
      LAYER via ;
        RECT 746.220 24.180 746.480 24.440 ;
        RECT 1131.700 24.180 1131.960 24.440 ;
      LAYER met2 ;
        RECT 1133.090 1220.330 1133.650 1228.680 ;
        RECT 1131.760 1220.190 1133.650 1220.330 ;
        RECT 1131.760 24.470 1131.900 1220.190 ;
        RECT 1133.090 1219.680 1133.650 1220.190 ;
        RECT 746.220 24.150 746.480 24.470 ;
        RECT 1131.700 24.150 1131.960 24.470 ;
        RECT 746.280 2.400 746.420 24.150 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1719.550 1210.640 1719.870 1210.700 ;
        RECT 1719.550 1210.500 1871.120 1210.640 ;
        RECT 1719.550 1210.440 1719.870 1210.500 ;
        RECT 1870.980 1210.300 1871.120 1210.500 ;
        RECT 1880.090 1210.300 1880.410 1210.360 ;
        RECT 1870.980 1210.160 1880.410 1210.300 ;
        RECT 1880.090 1210.100 1880.410 1210.160 ;
        RECT 1880.090 20.640 1880.410 20.700 ;
        RECT 1887.910 20.640 1888.230 20.700 ;
        RECT 1880.090 20.500 1888.230 20.640 ;
        RECT 1880.090 20.440 1880.410 20.500 ;
        RECT 1887.910 20.440 1888.230 20.500 ;
      LAYER via ;
        RECT 1719.580 1210.440 1719.840 1210.700 ;
        RECT 1880.120 1210.100 1880.380 1210.360 ;
        RECT 1880.120 20.440 1880.380 20.700 ;
        RECT 1887.940 20.440 1888.200 20.700 ;
      LAYER met2 ;
        RECT 1719.590 1219.680 1720.150 1228.680 ;
        RECT 1719.640 1210.730 1719.780 1219.680 ;
        RECT 1719.580 1210.410 1719.840 1210.730 ;
        RECT 1880.120 1210.070 1880.380 1210.390 ;
        RECT 1880.180 20.730 1880.320 1210.070 ;
        RECT 1880.120 20.410 1880.380 20.730 ;
        RECT 1887.940 20.410 1888.200 20.730 ;
        RECT 1888.000 2.400 1888.140 20.410 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1731.125 786.505 1731.295 821.015 ;
        RECT 1731.125 689.605 1731.295 724.455 ;
        RECT 1731.125 593.045 1731.295 627.895 ;
        RECT 1731.125 496.485 1731.295 531.335 ;
        RECT 1731.125 386.325 1731.295 434.775 ;
        RECT 1731.125 110.245 1731.295 137.955 ;
      LAYER mcon ;
        RECT 1731.125 820.845 1731.295 821.015 ;
        RECT 1731.125 724.285 1731.295 724.455 ;
        RECT 1731.125 627.725 1731.295 627.895 ;
        RECT 1731.125 531.165 1731.295 531.335 ;
        RECT 1731.125 434.605 1731.295 434.775 ;
        RECT 1731.125 137.785 1731.295 137.955 ;
      LAYER met1 ;
        RECT 1730.590 1124.960 1730.910 1125.020 ;
        RECT 1731.510 1124.960 1731.830 1125.020 ;
        RECT 1730.590 1124.820 1731.830 1124.960 ;
        RECT 1730.590 1124.760 1730.910 1124.820 ;
        RECT 1731.510 1124.760 1731.830 1124.820 ;
        RECT 1730.590 1028.400 1730.910 1028.460 ;
        RECT 1731.510 1028.400 1731.830 1028.460 ;
        RECT 1730.590 1028.260 1731.830 1028.400 ;
        RECT 1730.590 1028.200 1730.910 1028.260 ;
        RECT 1731.510 1028.200 1731.830 1028.260 ;
        RECT 1730.590 931.840 1730.910 931.900 ;
        RECT 1731.510 931.840 1731.830 931.900 ;
        RECT 1730.590 931.700 1731.830 931.840 ;
        RECT 1730.590 931.640 1730.910 931.700 ;
        RECT 1731.510 931.640 1731.830 931.700 ;
        RECT 1730.130 869.620 1730.450 869.680 ;
        RECT 1731.510 869.620 1731.830 869.680 ;
        RECT 1730.130 869.480 1731.830 869.620 ;
        RECT 1730.130 869.420 1730.450 869.480 ;
        RECT 1731.510 869.420 1731.830 869.480 ;
        RECT 1730.590 835.280 1730.910 835.340 ;
        RECT 1731.510 835.280 1731.830 835.340 ;
        RECT 1730.590 835.140 1731.830 835.280 ;
        RECT 1730.590 835.080 1730.910 835.140 ;
        RECT 1731.510 835.080 1731.830 835.140 ;
        RECT 1731.050 821.000 1731.370 821.060 ;
        RECT 1730.855 820.860 1731.370 821.000 ;
        RECT 1731.050 820.800 1731.370 820.860 ;
        RECT 1731.050 786.660 1731.370 786.720 ;
        RECT 1730.855 786.520 1731.370 786.660 ;
        RECT 1731.050 786.460 1731.370 786.520 ;
        RECT 1730.590 738.380 1730.910 738.440 ;
        RECT 1731.510 738.380 1731.830 738.440 ;
        RECT 1730.590 738.240 1731.830 738.380 ;
        RECT 1730.590 738.180 1730.910 738.240 ;
        RECT 1731.510 738.180 1731.830 738.240 ;
        RECT 1731.050 724.440 1731.370 724.500 ;
        RECT 1730.855 724.300 1731.370 724.440 ;
        RECT 1731.050 724.240 1731.370 724.300 ;
        RECT 1731.050 689.760 1731.370 689.820 ;
        RECT 1730.855 689.620 1731.370 689.760 ;
        RECT 1731.050 689.560 1731.370 689.620 ;
        RECT 1730.590 641.820 1730.910 641.880 ;
        RECT 1731.510 641.820 1731.830 641.880 ;
        RECT 1730.590 641.680 1731.830 641.820 ;
        RECT 1730.590 641.620 1730.910 641.680 ;
        RECT 1731.510 641.620 1731.830 641.680 ;
        RECT 1731.050 627.880 1731.370 627.940 ;
        RECT 1730.855 627.740 1731.370 627.880 ;
        RECT 1731.050 627.680 1731.370 627.740 ;
        RECT 1731.050 593.200 1731.370 593.260 ;
        RECT 1730.855 593.060 1731.370 593.200 ;
        RECT 1731.050 593.000 1731.370 593.060 ;
        RECT 1730.590 545.260 1730.910 545.320 ;
        RECT 1731.510 545.260 1731.830 545.320 ;
        RECT 1730.590 545.120 1731.830 545.260 ;
        RECT 1730.590 545.060 1730.910 545.120 ;
        RECT 1731.510 545.060 1731.830 545.120 ;
        RECT 1731.050 531.320 1731.370 531.380 ;
        RECT 1730.855 531.180 1731.370 531.320 ;
        RECT 1731.050 531.120 1731.370 531.180 ;
        RECT 1731.050 496.640 1731.370 496.700 ;
        RECT 1730.855 496.500 1731.370 496.640 ;
        RECT 1731.050 496.440 1731.370 496.500 ;
        RECT 1730.590 448.700 1730.910 448.760 ;
        RECT 1731.510 448.700 1731.830 448.760 ;
        RECT 1730.590 448.560 1731.830 448.700 ;
        RECT 1730.590 448.500 1730.910 448.560 ;
        RECT 1731.510 448.500 1731.830 448.560 ;
        RECT 1731.050 434.760 1731.370 434.820 ;
        RECT 1730.855 434.620 1731.370 434.760 ;
        RECT 1731.050 434.560 1731.370 434.620 ;
        RECT 1731.065 386.480 1731.355 386.525 ;
        RECT 1731.510 386.480 1731.830 386.540 ;
        RECT 1731.065 386.340 1731.830 386.480 ;
        RECT 1731.065 386.295 1731.355 386.340 ;
        RECT 1731.510 386.280 1731.830 386.340 ;
        RECT 1730.590 352.140 1730.910 352.200 ;
        RECT 1730.590 352.000 1731.280 352.140 ;
        RECT 1730.590 351.940 1730.910 352.000 ;
        RECT 1731.140 351.860 1731.280 352.000 ;
        RECT 1731.050 351.600 1731.370 351.860 ;
        RECT 1731.050 241.640 1731.370 241.700 ;
        RECT 1731.510 241.640 1731.830 241.700 ;
        RECT 1731.050 241.500 1731.830 241.640 ;
        RECT 1731.050 241.440 1731.370 241.500 ;
        RECT 1731.510 241.440 1731.830 241.500 ;
        RECT 1730.590 158.820 1730.910 159.080 ;
        RECT 1730.680 158.340 1730.820 158.820 ;
        RECT 1731.050 158.340 1731.370 158.400 ;
        RECT 1730.680 158.200 1731.370 158.340 ;
        RECT 1731.050 158.140 1731.370 158.200 ;
        RECT 1731.050 137.940 1731.370 138.000 ;
        RECT 1730.855 137.800 1731.370 137.940 ;
        RECT 1731.050 137.740 1731.370 137.800 ;
        RECT 1731.050 110.400 1731.370 110.460 ;
        RECT 1730.855 110.260 1731.370 110.400 ;
        RECT 1731.050 110.200 1731.370 110.260 ;
        RECT 1731.050 20.980 1731.370 21.040 ;
        RECT 1905.850 20.980 1906.170 21.040 ;
        RECT 1731.050 20.840 1906.170 20.980 ;
        RECT 1731.050 20.780 1731.370 20.840 ;
        RECT 1905.850 20.780 1906.170 20.840 ;
      LAYER via ;
        RECT 1730.620 1124.760 1730.880 1125.020 ;
        RECT 1731.540 1124.760 1731.800 1125.020 ;
        RECT 1730.620 1028.200 1730.880 1028.460 ;
        RECT 1731.540 1028.200 1731.800 1028.460 ;
        RECT 1730.620 931.640 1730.880 931.900 ;
        RECT 1731.540 931.640 1731.800 931.900 ;
        RECT 1730.160 869.420 1730.420 869.680 ;
        RECT 1731.540 869.420 1731.800 869.680 ;
        RECT 1730.620 835.080 1730.880 835.340 ;
        RECT 1731.540 835.080 1731.800 835.340 ;
        RECT 1731.080 820.800 1731.340 821.060 ;
        RECT 1731.080 786.460 1731.340 786.720 ;
        RECT 1730.620 738.180 1730.880 738.440 ;
        RECT 1731.540 738.180 1731.800 738.440 ;
        RECT 1731.080 724.240 1731.340 724.500 ;
        RECT 1731.080 689.560 1731.340 689.820 ;
        RECT 1730.620 641.620 1730.880 641.880 ;
        RECT 1731.540 641.620 1731.800 641.880 ;
        RECT 1731.080 627.680 1731.340 627.940 ;
        RECT 1731.080 593.000 1731.340 593.260 ;
        RECT 1730.620 545.060 1730.880 545.320 ;
        RECT 1731.540 545.060 1731.800 545.320 ;
        RECT 1731.080 531.120 1731.340 531.380 ;
        RECT 1731.080 496.440 1731.340 496.700 ;
        RECT 1730.620 448.500 1730.880 448.760 ;
        RECT 1731.540 448.500 1731.800 448.760 ;
        RECT 1731.080 434.560 1731.340 434.820 ;
        RECT 1731.540 386.280 1731.800 386.540 ;
        RECT 1730.620 351.940 1730.880 352.200 ;
        RECT 1731.080 351.600 1731.340 351.860 ;
        RECT 1731.080 241.440 1731.340 241.700 ;
        RECT 1731.540 241.440 1731.800 241.700 ;
        RECT 1730.620 158.820 1730.880 159.080 ;
        RECT 1731.080 158.140 1731.340 158.400 ;
        RECT 1731.080 137.740 1731.340 138.000 ;
        RECT 1731.080 110.200 1731.340 110.460 ;
        RECT 1731.080 20.780 1731.340 21.040 ;
        RECT 1905.880 20.780 1906.140 21.040 ;
      LAYER met2 ;
        RECT 1728.790 1221.010 1729.350 1228.680 ;
        RECT 1728.790 1220.870 1731.280 1221.010 ;
        RECT 1728.790 1219.680 1729.350 1220.870 ;
        RECT 1731.140 1196.530 1731.280 1220.870 ;
        RECT 1731.140 1196.390 1731.740 1196.530 ;
        RECT 1731.600 1125.050 1731.740 1196.390 ;
        RECT 1730.620 1124.730 1730.880 1125.050 ;
        RECT 1731.540 1124.730 1731.800 1125.050 ;
        RECT 1730.680 1124.450 1730.820 1124.730 ;
        RECT 1730.680 1124.310 1731.280 1124.450 ;
        RECT 1731.140 1076.850 1731.280 1124.310 ;
        RECT 1731.140 1076.710 1731.740 1076.850 ;
        RECT 1731.600 1028.490 1731.740 1076.710 ;
        RECT 1730.620 1028.170 1730.880 1028.490 ;
        RECT 1731.540 1028.170 1731.800 1028.490 ;
        RECT 1730.680 1027.890 1730.820 1028.170 ;
        RECT 1730.680 1027.750 1731.280 1027.890 ;
        RECT 1731.140 980.290 1731.280 1027.750 ;
        RECT 1731.140 980.150 1731.740 980.290 ;
        RECT 1731.600 931.930 1731.740 980.150 ;
        RECT 1730.620 931.610 1730.880 931.930 ;
        RECT 1731.540 931.610 1731.800 931.930 ;
        RECT 1730.680 931.330 1730.820 931.610 ;
        RECT 1730.680 931.190 1731.280 931.330 ;
        RECT 1731.140 917.845 1731.280 931.190 ;
        RECT 1730.150 917.475 1730.430 917.845 ;
        RECT 1731.070 917.475 1731.350 917.845 ;
        RECT 1730.220 869.710 1730.360 917.475 ;
        RECT 1730.160 869.390 1730.420 869.710 ;
        RECT 1731.540 869.390 1731.800 869.710 ;
        RECT 1731.600 835.370 1731.740 869.390 ;
        RECT 1730.620 835.050 1730.880 835.370 ;
        RECT 1731.540 835.050 1731.800 835.370 ;
        RECT 1730.680 834.770 1730.820 835.050 ;
        RECT 1730.680 834.630 1731.280 834.770 ;
        RECT 1731.140 821.090 1731.280 834.630 ;
        RECT 1731.080 820.770 1731.340 821.090 ;
        RECT 1731.080 786.430 1731.340 786.750 ;
        RECT 1731.140 772.890 1731.280 786.430 ;
        RECT 1731.140 772.750 1731.740 772.890 ;
        RECT 1731.600 738.470 1731.740 772.750 ;
        RECT 1730.620 738.210 1730.880 738.470 ;
        RECT 1730.620 738.150 1731.280 738.210 ;
        RECT 1731.540 738.150 1731.800 738.470 ;
        RECT 1730.680 738.070 1731.280 738.150 ;
        RECT 1731.140 724.530 1731.280 738.070 ;
        RECT 1731.080 724.210 1731.340 724.530 ;
        RECT 1731.080 689.530 1731.340 689.850 ;
        RECT 1731.140 676.330 1731.280 689.530 ;
        RECT 1731.140 676.190 1731.740 676.330 ;
        RECT 1731.600 641.910 1731.740 676.190 ;
        RECT 1730.620 641.650 1730.880 641.910 ;
        RECT 1730.620 641.590 1731.280 641.650 ;
        RECT 1731.540 641.590 1731.800 641.910 ;
        RECT 1730.680 641.510 1731.280 641.590 ;
        RECT 1731.140 627.970 1731.280 641.510 ;
        RECT 1731.080 627.650 1731.340 627.970 ;
        RECT 1731.080 592.970 1731.340 593.290 ;
        RECT 1731.140 579.770 1731.280 592.970 ;
        RECT 1731.140 579.630 1731.740 579.770 ;
        RECT 1731.600 545.350 1731.740 579.630 ;
        RECT 1730.620 545.090 1730.880 545.350 ;
        RECT 1730.620 545.030 1731.280 545.090 ;
        RECT 1731.540 545.030 1731.800 545.350 ;
        RECT 1730.680 544.950 1731.280 545.030 ;
        RECT 1731.140 531.410 1731.280 544.950 ;
        RECT 1731.080 531.090 1731.340 531.410 ;
        RECT 1731.080 496.410 1731.340 496.730 ;
        RECT 1731.140 483.210 1731.280 496.410 ;
        RECT 1731.140 483.070 1731.740 483.210 ;
        RECT 1731.600 448.790 1731.740 483.070 ;
        RECT 1730.620 448.530 1730.880 448.790 ;
        RECT 1730.620 448.470 1731.280 448.530 ;
        RECT 1731.540 448.470 1731.800 448.790 ;
        RECT 1730.680 448.390 1731.280 448.470 ;
        RECT 1731.140 434.850 1731.280 448.390 ;
        RECT 1731.080 434.530 1731.340 434.850 ;
        RECT 1731.540 386.250 1731.800 386.570 ;
        RECT 1731.600 386.085 1731.740 386.250 ;
        RECT 1730.610 385.715 1730.890 386.085 ;
        RECT 1731.530 385.715 1731.810 386.085 ;
        RECT 1730.680 352.230 1730.820 385.715 ;
        RECT 1730.620 351.910 1730.880 352.230 ;
        RECT 1731.080 351.570 1731.340 351.890 ;
        RECT 1731.140 303.690 1731.280 351.570 ;
        RECT 1731.140 303.550 1731.740 303.690 ;
        RECT 1731.600 241.730 1731.740 303.550 ;
        RECT 1731.080 241.410 1731.340 241.730 ;
        RECT 1731.540 241.410 1731.800 241.730 ;
        RECT 1731.140 241.130 1731.280 241.410 ;
        RECT 1730.680 240.990 1731.280 241.130 ;
        RECT 1730.680 207.130 1730.820 240.990 ;
        RECT 1730.680 206.990 1731.280 207.130 ;
        RECT 1731.140 193.530 1731.280 206.990 ;
        RECT 1730.680 193.390 1731.280 193.530 ;
        RECT 1730.680 159.110 1730.820 193.390 ;
        RECT 1730.620 158.790 1730.880 159.110 ;
        RECT 1731.080 158.110 1731.340 158.430 ;
        RECT 1731.140 138.030 1731.280 158.110 ;
        RECT 1731.080 137.710 1731.340 138.030 ;
        RECT 1731.080 110.170 1731.340 110.490 ;
        RECT 1731.140 21.070 1731.280 110.170 ;
        RECT 1731.080 20.750 1731.340 21.070 ;
        RECT 1905.880 20.750 1906.140 21.070 ;
        RECT 1905.940 2.400 1906.080 20.750 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
      LAYER via2 ;
        RECT 1730.150 917.520 1730.430 917.800 ;
        RECT 1731.070 917.520 1731.350 917.800 ;
        RECT 1730.610 385.760 1730.890 386.040 ;
        RECT 1731.530 385.760 1731.810 386.040 ;
      LAYER met3 ;
        RECT 1730.125 917.810 1730.455 917.825 ;
        RECT 1731.045 917.810 1731.375 917.825 ;
        RECT 1730.125 917.510 1731.375 917.810 ;
        RECT 1730.125 917.495 1730.455 917.510 ;
        RECT 1731.045 917.495 1731.375 917.510 ;
        RECT 1730.585 386.050 1730.915 386.065 ;
        RECT 1731.505 386.050 1731.835 386.065 ;
        RECT 1730.585 385.750 1731.835 386.050 ;
        RECT 1730.585 385.735 1730.915 385.750 ;
        RECT 1731.505 385.735 1731.835 385.750 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1738.410 21.320 1738.730 21.380 ;
        RECT 1923.330 21.320 1923.650 21.380 ;
        RECT 1738.410 21.180 1923.650 21.320 ;
        RECT 1738.410 21.120 1738.730 21.180 ;
        RECT 1923.330 21.120 1923.650 21.180 ;
      LAYER via ;
        RECT 1738.440 21.120 1738.700 21.380 ;
        RECT 1923.360 21.120 1923.620 21.380 ;
      LAYER met2 ;
        RECT 1737.990 1220.330 1738.550 1228.680 ;
        RECT 1737.990 1219.680 1738.640 1220.330 ;
        RECT 1738.500 21.410 1738.640 1219.680 ;
        RECT 1738.440 21.090 1738.700 21.410 ;
        RECT 1923.360 21.090 1923.620 21.410 ;
        RECT 1923.420 2.400 1923.560 21.090 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1747.150 1208.600 1747.470 1208.660 ;
        RECT 1752.210 1208.600 1752.530 1208.660 ;
        RECT 1747.150 1208.460 1752.530 1208.600 ;
        RECT 1747.150 1208.400 1747.470 1208.460 ;
        RECT 1752.210 1208.400 1752.530 1208.460 ;
        RECT 1752.210 21.660 1752.530 21.720 ;
        RECT 1941.270 21.660 1941.590 21.720 ;
        RECT 1752.210 21.520 1941.590 21.660 ;
        RECT 1752.210 21.460 1752.530 21.520 ;
        RECT 1941.270 21.460 1941.590 21.520 ;
      LAYER via ;
        RECT 1747.180 1208.400 1747.440 1208.660 ;
        RECT 1752.240 1208.400 1752.500 1208.660 ;
        RECT 1752.240 21.460 1752.500 21.720 ;
        RECT 1941.300 21.460 1941.560 21.720 ;
      LAYER met2 ;
        RECT 1747.190 1219.680 1747.750 1228.680 ;
        RECT 1747.240 1208.690 1747.380 1219.680 ;
        RECT 1747.180 1208.370 1747.440 1208.690 ;
        RECT 1752.240 1208.370 1752.500 1208.690 ;
        RECT 1752.300 21.750 1752.440 1208.370 ;
        RECT 1752.240 21.430 1752.500 21.750 ;
        RECT 1941.300 21.430 1941.560 21.750 ;
        RECT 1941.360 2.400 1941.500 21.430 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1759.110 22.340 1759.430 22.400 ;
        RECT 1959.210 22.340 1959.530 22.400 ;
        RECT 1759.110 22.200 1959.530 22.340 ;
        RECT 1759.110 22.140 1759.430 22.200 ;
        RECT 1959.210 22.140 1959.530 22.200 ;
      LAYER via ;
        RECT 1759.140 22.140 1759.400 22.400 ;
        RECT 1959.240 22.140 1959.500 22.400 ;
      LAYER met2 ;
        RECT 1756.390 1220.330 1756.950 1228.680 ;
        RECT 1756.390 1220.190 1758.880 1220.330 ;
        RECT 1756.390 1219.680 1756.950 1220.190 ;
        RECT 1758.740 1196.530 1758.880 1220.190 ;
        RECT 1758.740 1196.390 1759.340 1196.530 ;
        RECT 1759.200 22.430 1759.340 1196.390 ;
        RECT 1759.140 22.110 1759.400 22.430 ;
        RECT 1959.240 22.110 1959.500 22.430 ;
        RECT 1959.300 2.400 1959.440 22.110 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1765.550 32.200 1765.870 32.260 ;
        RECT 1976.690 32.200 1977.010 32.260 ;
        RECT 1765.550 32.060 1977.010 32.200 ;
        RECT 1765.550 32.000 1765.870 32.060 ;
        RECT 1976.690 32.000 1977.010 32.060 ;
      LAYER via ;
        RECT 1765.580 32.000 1765.840 32.260 ;
        RECT 1976.720 32.000 1976.980 32.260 ;
      LAYER met2 ;
        RECT 1765.130 1220.330 1765.690 1228.680 ;
        RECT 1765.130 1219.680 1765.780 1220.330 ;
        RECT 1765.640 32.290 1765.780 1219.680 ;
        RECT 1765.580 31.970 1765.840 32.290 ;
        RECT 1976.720 31.970 1976.980 32.290 ;
        RECT 1976.780 20.130 1976.920 31.970 ;
        RECT 1976.780 19.990 1977.380 20.130 ;
        RECT 1977.240 2.400 1977.380 19.990 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1774.290 1207.580 1774.610 1207.640 ;
        RECT 1779.350 1207.580 1779.670 1207.640 ;
        RECT 1774.290 1207.440 1779.670 1207.580 ;
        RECT 1774.290 1207.380 1774.610 1207.440 ;
        RECT 1779.350 1207.380 1779.670 1207.440 ;
        RECT 1779.350 31.860 1779.670 31.920 ;
        RECT 1995.090 31.860 1995.410 31.920 ;
        RECT 1779.350 31.720 1995.410 31.860 ;
        RECT 1779.350 31.660 1779.670 31.720 ;
        RECT 1995.090 31.660 1995.410 31.720 ;
      LAYER via ;
        RECT 1774.320 1207.380 1774.580 1207.640 ;
        RECT 1779.380 1207.380 1779.640 1207.640 ;
        RECT 1779.380 31.660 1779.640 31.920 ;
        RECT 1995.120 31.660 1995.380 31.920 ;
      LAYER met2 ;
        RECT 1774.330 1219.680 1774.890 1228.680 ;
        RECT 1774.380 1207.670 1774.520 1219.680 ;
        RECT 1774.320 1207.350 1774.580 1207.670 ;
        RECT 1779.380 1207.350 1779.640 1207.670 ;
        RECT 1779.440 31.950 1779.580 1207.350 ;
        RECT 1779.380 31.630 1779.640 31.950 ;
        RECT 1995.120 31.630 1995.380 31.950 ;
        RECT 1995.180 2.400 1995.320 31.630 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1941.805 20.825 1941.975 21.675 ;
      LAYER mcon ;
        RECT 1941.805 21.505 1941.975 21.675 ;
      LAYER met1 ;
        RECT 1922.410 1208.940 1922.730 1209.000 ;
        RECT 1898.120 1208.800 1922.730 1208.940 ;
        RECT 1898.120 1208.600 1898.260 1208.800 ;
        RECT 1922.410 1208.740 1922.730 1208.800 ;
        RECT 1801.520 1208.460 1898.260 1208.600 ;
        RECT 1785.330 1207.920 1785.650 1207.980 ;
        RECT 1801.520 1207.920 1801.660 1208.460 ;
        RECT 1785.330 1207.780 1801.660 1207.920 ;
        RECT 1785.330 1207.720 1785.650 1207.780 ;
        RECT 1922.410 620.540 1922.730 620.800 ;
        RECT 1922.500 620.120 1922.640 620.540 ;
        RECT 1922.410 619.860 1922.730 620.120 ;
        RECT 1941.745 21.660 1942.035 21.705 ;
        RECT 1941.745 21.520 1970.020 21.660 ;
        RECT 1941.745 21.475 1942.035 21.520 ;
        RECT 1969.880 21.320 1970.020 21.520 ;
        RECT 2012.570 21.320 2012.890 21.380 ;
        RECT 1969.880 21.180 2012.890 21.320 ;
        RECT 2012.570 21.120 2012.890 21.180 ;
        RECT 1924.250 20.980 1924.570 21.040 ;
        RECT 1941.745 20.980 1942.035 21.025 ;
        RECT 1924.250 20.840 1942.035 20.980 ;
        RECT 1924.250 20.780 1924.570 20.840 ;
        RECT 1941.745 20.795 1942.035 20.840 ;
      LAYER via ;
        RECT 1922.440 1208.740 1922.700 1209.000 ;
        RECT 1785.360 1207.720 1785.620 1207.980 ;
        RECT 1922.440 620.540 1922.700 620.800 ;
        RECT 1922.440 619.860 1922.700 620.120 ;
        RECT 2012.600 21.120 2012.860 21.380 ;
        RECT 1924.280 20.780 1924.540 21.040 ;
      LAYER met2 ;
        RECT 1783.530 1220.330 1784.090 1228.680 ;
        RECT 1783.530 1220.190 1785.560 1220.330 ;
        RECT 1783.530 1219.680 1784.090 1220.190 ;
        RECT 1785.420 1208.010 1785.560 1220.190 ;
        RECT 1922.440 1208.710 1922.700 1209.030 ;
        RECT 1785.360 1207.690 1785.620 1208.010 ;
        RECT 1922.500 620.830 1922.640 1208.710 ;
        RECT 1922.440 620.510 1922.700 620.830 ;
        RECT 1922.440 619.830 1922.700 620.150 ;
        RECT 1922.500 41.890 1922.640 619.830 ;
        RECT 1922.500 41.750 1924.480 41.890 ;
        RECT 1924.340 21.070 1924.480 41.750 ;
        RECT 2012.600 21.090 2012.860 21.410 ;
        RECT 1924.280 20.750 1924.540 21.070 ;
        RECT 2012.660 2.400 2012.800 21.090 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1793.150 31.520 1793.470 31.580 ;
        RECT 2030.510 31.520 2030.830 31.580 ;
        RECT 1793.150 31.380 2030.830 31.520 ;
        RECT 1793.150 31.320 1793.470 31.380 ;
        RECT 2030.510 31.320 2030.830 31.380 ;
      LAYER via ;
        RECT 1793.180 31.320 1793.440 31.580 ;
        RECT 2030.540 31.320 2030.800 31.580 ;
      LAYER met2 ;
        RECT 1792.730 1220.330 1793.290 1228.680 ;
        RECT 1792.730 1219.680 1793.380 1220.330 ;
        RECT 1793.240 31.610 1793.380 1219.680 ;
        RECT 1793.180 31.290 1793.440 31.610 ;
        RECT 2030.540 31.290 2030.800 31.610 ;
        RECT 2030.600 2.400 2030.740 31.290 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1898.105 1208.955 1898.275 1210.995 ;
        RECT 1897.645 1208.785 1898.275 1208.955 ;
        RECT 1969.405 21.165 1969.575 22.015 ;
      LAYER mcon ;
        RECT 1898.105 1210.825 1898.275 1210.995 ;
        RECT 1969.405 21.845 1969.575 22.015 ;
      LAYER met1 ;
        RECT 1898.045 1210.980 1898.335 1211.025 ;
        RECT 1943.110 1210.980 1943.430 1211.040 ;
        RECT 1898.045 1210.840 1943.430 1210.980 ;
        RECT 1898.045 1210.795 1898.335 1210.840 ;
        RECT 1943.110 1210.780 1943.430 1210.840 ;
        RECT 1845.590 1208.940 1845.910 1209.000 ;
        RECT 1897.585 1208.940 1897.875 1208.985 ;
        RECT 1845.590 1208.800 1897.875 1208.940 ;
        RECT 1845.590 1208.740 1845.910 1208.800 ;
        RECT 1897.585 1208.755 1897.875 1208.800 ;
        RECT 1801.890 1208.260 1802.210 1208.320 ;
        RECT 1845.590 1208.260 1845.910 1208.320 ;
        RECT 1801.890 1208.120 1845.910 1208.260 ;
        RECT 1801.890 1208.060 1802.210 1208.120 ;
        RECT 1845.590 1208.060 1845.910 1208.120 ;
        RECT 1969.345 22.000 1969.635 22.045 ;
        RECT 1969.345 21.860 1970.480 22.000 ;
        RECT 1969.345 21.815 1969.635 21.860 ;
        RECT 1970.340 21.660 1970.480 21.860 ;
        RECT 2048.450 21.660 2048.770 21.720 ;
        RECT 1970.340 21.520 2048.770 21.660 ;
        RECT 2048.450 21.460 2048.770 21.520 ;
        RECT 1943.110 21.320 1943.430 21.380 ;
        RECT 1969.345 21.320 1969.635 21.365 ;
        RECT 1943.110 21.180 1969.635 21.320 ;
        RECT 1943.110 21.120 1943.430 21.180 ;
        RECT 1969.345 21.135 1969.635 21.180 ;
      LAYER via ;
        RECT 1943.140 1210.780 1943.400 1211.040 ;
        RECT 1845.620 1208.740 1845.880 1209.000 ;
        RECT 1801.920 1208.060 1802.180 1208.320 ;
        RECT 1845.620 1208.060 1845.880 1208.320 ;
        RECT 2048.480 21.460 2048.740 21.720 ;
        RECT 1943.140 21.120 1943.400 21.380 ;
      LAYER met2 ;
        RECT 1801.930 1219.680 1802.490 1228.680 ;
        RECT 1801.980 1208.350 1802.120 1219.680 ;
        RECT 1943.140 1210.750 1943.400 1211.070 ;
        RECT 1845.620 1208.710 1845.880 1209.030 ;
        RECT 1845.680 1208.350 1845.820 1208.710 ;
        RECT 1801.920 1208.030 1802.180 1208.350 ;
        RECT 1845.620 1208.030 1845.880 1208.350 ;
        RECT 1943.200 21.410 1943.340 1210.750 ;
        RECT 2048.480 21.430 2048.740 21.750 ;
        RECT 1943.140 21.090 1943.400 21.410 ;
        RECT 2048.540 2.400 2048.680 21.430 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 917.845 23.545 918.015 27.455 ;
        RECT 941.765 21.845 941.935 23.715 ;
      LAYER mcon ;
        RECT 917.845 27.285 918.015 27.455 ;
        RECT 941.765 23.545 941.935 23.715 ;
      LAYER met1 ;
        RECT 1003.790 1209.960 1004.110 1210.020 ;
        RECT 1142.250 1209.960 1142.570 1210.020 ;
        RECT 1003.790 1209.820 1142.570 1209.960 ;
        RECT 1003.790 1209.760 1004.110 1209.820 ;
        RECT 1142.250 1209.760 1142.570 1209.820 ;
        RECT 917.310 27.440 917.630 27.500 ;
        RECT 917.785 27.440 918.075 27.485 ;
        RECT 917.310 27.300 918.075 27.440 ;
        RECT 917.310 27.240 917.630 27.300 ;
        RECT 917.785 27.255 918.075 27.300 ;
        RECT 763.670 26.760 763.990 26.820 ;
        RECT 763.670 26.620 810.820 26.760 ;
        RECT 763.670 26.560 763.990 26.620 ;
        RECT 810.680 26.420 810.820 26.620 ;
        RECT 893.390 26.420 893.710 26.480 ;
        RECT 810.680 26.280 893.710 26.420 ;
        RECT 893.390 26.220 893.710 26.280 ;
        RECT 917.785 23.700 918.075 23.745 ;
        RECT 941.705 23.700 941.995 23.745 ;
        RECT 917.785 23.560 941.995 23.700 ;
        RECT 917.785 23.515 918.075 23.560 ;
        RECT 941.705 23.515 941.995 23.560 ;
        RECT 941.705 22.000 941.995 22.045 ;
        RECT 941.705 21.860 946.060 22.000 ;
        RECT 941.705 21.815 941.995 21.860 ;
        RECT 945.920 21.660 946.060 21.860 ;
        RECT 1003.790 21.660 1004.110 21.720 ;
        RECT 945.920 21.520 1004.110 21.660 ;
        RECT 1003.790 21.460 1004.110 21.520 ;
      LAYER via ;
        RECT 1003.820 1209.760 1004.080 1210.020 ;
        RECT 1142.280 1209.760 1142.540 1210.020 ;
        RECT 917.340 27.240 917.600 27.500 ;
        RECT 763.700 26.560 763.960 26.820 ;
        RECT 893.420 26.220 893.680 26.480 ;
        RECT 1003.820 21.460 1004.080 21.720 ;
      LAYER met2 ;
        RECT 1142.290 1219.680 1142.850 1228.680 ;
        RECT 1142.340 1210.050 1142.480 1219.680 ;
        RECT 1003.820 1209.730 1004.080 1210.050 ;
        RECT 1142.280 1209.730 1142.540 1210.050 ;
        RECT 917.340 27.210 917.600 27.530 ;
        RECT 917.400 27.045 917.540 27.210 ;
        RECT 763.700 26.530 763.960 26.850 ;
        RECT 893.410 26.675 893.690 27.045 ;
        RECT 917.330 26.675 917.610 27.045 ;
        RECT 763.760 2.400 763.900 26.530 ;
        RECT 893.480 26.510 893.620 26.675 ;
        RECT 893.420 26.190 893.680 26.510 ;
        RECT 1003.880 21.750 1004.020 1209.730 ;
        RECT 1003.820 21.430 1004.080 21.750 ;
        RECT 763.550 -4.800 764.110 2.400 ;
      LAYER via2 ;
        RECT 893.410 26.720 893.690 27.000 ;
        RECT 917.330 26.720 917.610 27.000 ;
      LAYER met3 ;
        RECT 893.385 27.010 893.715 27.025 ;
        RECT 917.305 27.010 917.635 27.025 ;
        RECT 893.385 26.710 917.635 27.010 ;
        RECT 893.385 26.695 893.715 26.710 ;
        RECT 917.305 26.695 917.635 26.710 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1813.390 31.180 1813.710 31.240 ;
        RECT 2066.390 31.180 2066.710 31.240 ;
        RECT 1813.390 31.040 2066.710 31.180 ;
        RECT 1813.390 30.980 1813.710 31.040 ;
        RECT 2066.390 30.980 2066.710 31.040 ;
      LAYER via ;
        RECT 1813.420 30.980 1813.680 31.240 ;
        RECT 2066.420 30.980 2066.680 31.240 ;
      LAYER met2 ;
        RECT 1811.130 1220.330 1811.690 1228.680 ;
        RECT 1811.130 1220.190 1813.620 1220.330 ;
        RECT 1811.130 1219.680 1811.690 1220.190 ;
        RECT 1813.480 31.270 1813.620 1220.190 ;
        RECT 1813.420 30.950 1813.680 31.270 ;
        RECT 2066.420 30.950 2066.680 31.270 ;
        RECT 2066.480 2.400 2066.620 30.950 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1820.750 30.840 1821.070 30.900 ;
        RECT 2084.330 30.840 2084.650 30.900 ;
        RECT 1820.750 30.700 2084.650 30.840 ;
        RECT 1820.750 30.640 1821.070 30.700 ;
        RECT 2084.330 30.640 2084.650 30.700 ;
      LAYER via ;
        RECT 1820.780 30.640 1821.040 30.900 ;
        RECT 2084.360 30.640 2084.620 30.900 ;
      LAYER met2 ;
        RECT 1820.330 1220.330 1820.890 1228.680 ;
        RECT 1820.330 1219.680 1820.980 1220.330 ;
        RECT 1820.840 30.930 1820.980 1219.680 ;
        RECT 1820.780 30.610 1821.040 30.930 ;
        RECT 2084.360 30.610 2084.620 30.930 ;
        RECT 2084.420 2.400 2084.560 30.610 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1829.490 1207.580 1829.810 1207.640 ;
        RECT 1835.010 1207.580 1835.330 1207.640 ;
        RECT 1829.490 1207.440 1835.330 1207.580 ;
        RECT 1829.490 1207.380 1829.810 1207.440 ;
        RECT 1835.010 1207.380 1835.330 1207.440 ;
        RECT 1835.010 18.940 1835.330 19.000 ;
        RECT 2101.810 18.940 2102.130 19.000 ;
        RECT 1835.010 18.800 2102.130 18.940 ;
        RECT 1835.010 18.740 1835.330 18.800 ;
        RECT 2101.810 18.740 2102.130 18.800 ;
      LAYER via ;
        RECT 1829.520 1207.380 1829.780 1207.640 ;
        RECT 1835.040 1207.380 1835.300 1207.640 ;
        RECT 1835.040 18.740 1835.300 19.000 ;
        RECT 2101.840 18.740 2102.100 19.000 ;
      LAYER met2 ;
        RECT 1829.530 1219.680 1830.090 1228.680 ;
        RECT 1829.580 1207.670 1829.720 1219.680 ;
        RECT 1829.520 1207.350 1829.780 1207.670 ;
        RECT 1835.040 1207.350 1835.300 1207.670 ;
        RECT 1835.100 19.030 1835.240 1207.350 ;
        RECT 1835.040 18.710 1835.300 19.030 ;
        RECT 2101.840 18.710 2102.100 19.030 ;
        RECT 2101.900 2.400 2102.040 18.710 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1849.805 1207.425 1849.975 1214.735 ;
      LAYER mcon ;
        RECT 1849.805 1214.565 1849.975 1214.735 ;
      LAYER met1 ;
        RECT 1838.690 1214.720 1839.010 1214.780 ;
        RECT 1849.745 1214.720 1850.035 1214.765 ;
        RECT 1838.690 1214.580 1850.035 1214.720 ;
        RECT 1838.690 1214.520 1839.010 1214.580 ;
        RECT 1849.745 1214.535 1850.035 1214.580 ;
        RECT 1956.450 1208.600 1956.770 1208.660 ;
        RECT 1905.020 1208.460 1956.770 1208.600 ;
        RECT 1905.020 1207.920 1905.160 1208.460 ;
        RECT 1956.450 1208.400 1956.770 1208.460 ;
        RECT 1899.500 1207.780 1905.160 1207.920 ;
        RECT 1849.745 1207.580 1850.035 1207.625 ;
        RECT 1899.500 1207.580 1899.640 1207.780 ;
        RECT 1849.745 1207.440 1850.420 1207.580 ;
        RECT 1849.745 1207.395 1850.035 1207.440 ;
        RECT 1850.280 1207.240 1850.420 1207.440 ;
        RECT 1856.260 1207.440 1862.840 1207.580 ;
        RECT 1856.260 1207.240 1856.400 1207.440 ;
        RECT 1850.280 1207.100 1856.400 1207.240 ;
        RECT 1862.700 1207.240 1862.840 1207.440 ;
        RECT 1876.960 1207.440 1899.640 1207.580 ;
        RECT 1876.960 1207.240 1877.100 1207.440 ;
        RECT 1862.700 1207.100 1877.100 1207.240 ;
        RECT 1973.470 22.340 1973.790 22.400 ;
        RECT 2119.750 22.340 2120.070 22.400 ;
        RECT 1973.470 22.200 2120.070 22.340 ;
        RECT 1973.470 22.140 1973.790 22.200 ;
        RECT 2119.750 22.140 2120.070 22.200 ;
      LAYER via ;
        RECT 1838.720 1214.520 1838.980 1214.780 ;
        RECT 1956.480 1208.400 1956.740 1208.660 ;
        RECT 1973.500 22.140 1973.760 22.400 ;
        RECT 2119.780 22.140 2120.040 22.400 ;
      LAYER met2 ;
        RECT 1838.730 1219.680 1839.290 1228.680 ;
        RECT 1838.780 1214.810 1838.920 1219.680 ;
        RECT 1838.720 1214.490 1838.980 1214.810 ;
        RECT 1956.480 1208.370 1956.740 1208.690 ;
        RECT 1956.540 22.965 1956.680 1208.370 ;
        RECT 1956.470 22.595 1956.750 22.965 ;
        RECT 1973.490 22.595 1973.770 22.965 ;
        RECT 1973.560 22.430 1973.700 22.595 ;
        RECT 1973.500 22.110 1973.760 22.430 ;
        RECT 2119.780 22.110 2120.040 22.430 ;
        RECT 2119.840 2.400 2119.980 22.110 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
      LAYER via2 ;
        RECT 1956.470 22.640 1956.750 22.920 ;
        RECT 1973.490 22.640 1973.770 22.920 ;
      LAYER met3 ;
        RECT 1956.445 22.930 1956.775 22.945 ;
        RECT 1973.465 22.930 1973.795 22.945 ;
        RECT 1956.445 22.630 1973.795 22.930 ;
        RECT 1956.445 22.615 1956.775 22.630 ;
        RECT 1973.465 22.615 1973.795 22.630 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1848.350 38.320 1848.670 38.380 ;
        RECT 2137.690 38.320 2138.010 38.380 ;
        RECT 1848.350 38.180 2138.010 38.320 ;
        RECT 1848.350 38.120 1848.670 38.180 ;
        RECT 2137.690 38.120 2138.010 38.180 ;
      LAYER via ;
        RECT 1848.380 38.120 1848.640 38.380 ;
        RECT 2137.720 38.120 2137.980 38.380 ;
      LAYER met2 ;
        RECT 1847.930 1220.330 1848.490 1228.680 ;
        RECT 1847.930 1219.680 1848.580 1220.330 ;
        RECT 1848.440 38.410 1848.580 1219.680 ;
        RECT 1848.380 38.090 1848.640 38.410 ;
        RECT 2137.720 38.090 2137.980 38.410 ;
        RECT 2137.780 2.400 2137.920 38.090 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2139.145 21.845 2139.315 24.055 ;
      LAYER mcon ;
        RECT 2139.145 23.885 2139.315 24.055 ;
      LAYER met1 ;
        RECT 1956.910 1209.620 1957.230 1209.680 ;
        RECT 1921.580 1209.480 1957.230 1209.620 ;
        RECT 1857.090 1209.280 1857.410 1209.340 ;
        RECT 1921.580 1209.280 1921.720 1209.480 ;
        RECT 1956.910 1209.420 1957.230 1209.480 ;
        RECT 1857.090 1209.140 1921.720 1209.280 ;
        RECT 1857.090 1209.080 1857.410 1209.140 ;
        RECT 2139.085 24.040 2139.375 24.085 ;
        RECT 2155.630 24.040 2155.950 24.100 ;
        RECT 2139.085 23.900 2155.950 24.040 ;
        RECT 2139.085 23.855 2139.375 23.900 ;
        RECT 2155.630 23.840 2155.950 23.900 ;
        RECT 1959.760 22.200 1973.240 22.340 ;
        RECT 1956.910 22.000 1957.230 22.060 ;
        RECT 1959.760 22.000 1959.900 22.200 ;
        RECT 1956.910 21.860 1959.900 22.000 ;
        RECT 1973.100 22.000 1973.240 22.200 ;
        RECT 2139.085 22.000 2139.375 22.045 ;
        RECT 1973.100 21.860 2139.375 22.000 ;
        RECT 1956.910 21.800 1957.230 21.860 ;
        RECT 2139.085 21.815 2139.375 21.860 ;
      LAYER via ;
        RECT 1857.120 1209.080 1857.380 1209.340 ;
        RECT 1956.940 1209.420 1957.200 1209.680 ;
        RECT 2155.660 23.840 2155.920 24.100 ;
        RECT 1956.940 21.800 1957.200 22.060 ;
      LAYER met2 ;
        RECT 1857.130 1219.680 1857.690 1228.680 ;
        RECT 1857.180 1209.370 1857.320 1219.680 ;
        RECT 1956.940 1209.390 1957.200 1209.710 ;
        RECT 1857.120 1209.050 1857.380 1209.370 ;
        RECT 1957.000 22.090 1957.140 1209.390 ;
        RECT 2155.660 23.810 2155.920 24.130 ;
        RECT 1956.940 21.770 1957.200 22.090 ;
        RECT 2155.720 2.400 2155.860 23.810 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2172.650 37.980 2172.970 38.040 ;
        RECT 1882.940 37.840 2172.970 37.980 ;
        RECT 1868.590 37.300 1868.910 37.360 ;
        RECT 1882.940 37.300 1883.080 37.840 ;
        RECT 2172.650 37.780 2172.970 37.840 ;
        RECT 1868.590 37.160 1883.080 37.300 ;
        RECT 1868.590 37.100 1868.910 37.160 ;
      LAYER via ;
        RECT 1868.620 37.100 1868.880 37.360 ;
        RECT 2172.680 37.780 2172.940 38.040 ;
      LAYER met2 ;
        RECT 1866.330 1220.330 1866.890 1228.680 ;
        RECT 1866.330 1220.190 1868.820 1220.330 ;
        RECT 1866.330 1219.680 1866.890 1220.190 ;
        RECT 1868.680 37.390 1868.820 1220.190 ;
        RECT 2172.680 37.750 2172.940 38.070 ;
        RECT 1868.620 37.070 1868.880 37.390 ;
        RECT 2172.740 8.570 2172.880 37.750 ;
        RECT 2172.740 8.430 2173.340 8.570 ;
        RECT 2173.200 2.400 2173.340 8.430 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1970.325 96.645 1970.495 144.755 ;
        RECT 2163.065 24.225 2164.155 24.395 ;
        RECT 2163.065 23.885 2163.235 24.225 ;
        RECT 2018.165 21.165 2018.335 23.035 ;
        RECT 2062.325 21.165 2062.495 23.035 ;
      LAYER mcon ;
        RECT 1970.325 144.585 1970.495 144.755 ;
        RECT 2163.985 24.225 2164.155 24.395 ;
        RECT 2018.165 22.865 2018.335 23.035 ;
        RECT 2062.325 22.865 2062.495 23.035 ;
      LAYER met1 ;
        RECT 1875.490 1209.960 1875.810 1210.020 ;
        RECT 1970.250 1209.960 1970.570 1210.020 ;
        RECT 1875.490 1209.820 1970.570 1209.960 ;
        RECT 1875.490 1209.760 1875.810 1209.820 ;
        RECT 1970.250 1209.760 1970.570 1209.820 ;
        RECT 1968.870 1159.300 1969.190 1159.360 ;
        RECT 1969.790 1159.300 1970.110 1159.360 ;
        RECT 1968.870 1159.160 1970.110 1159.300 ;
        RECT 1968.870 1159.100 1969.190 1159.160 ;
        RECT 1969.790 1159.100 1970.110 1159.160 ;
        RECT 1969.790 158.680 1970.110 158.740 ;
        RECT 1970.710 158.680 1971.030 158.740 ;
        RECT 1969.790 158.540 1971.030 158.680 ;
        RECT 1969.790 158.480 1970.110 158.540 ;
        RECT 1970.710 158.480 1971.030 158.540 ;
        RECT 1970.265 144.740 1970.555 144.785 ;
        RECT 1970.710 144.740 1971.030 144.800 ;
        RECT 1970.265 144.600 1971.030 144.740 ;
        RECT 1970.265 144.555 1970.555 144.600 ;
        RECT 1970.710 144.540 1971.030 144.600 ;
        RECT 1970.250 96.800 1970.570 96.860 ;
        RECT 1970.055 96.660 1970.570 96.800 ;
        RECT 1970.250 96.600 1970.570 96.660 ;
        RECT 2163.925 24.380 2164.215 24.425 ;
        RECT 2191.050 24.380 2191.370 24.440 ;
        RECT 2163.925 24.240 2191.370 24.380 ;
        RECT 2163.925 24.195 2164.215 24.240 ;
        RECT 2191.050 24.180 2191.370 24.240 ;
        RECT 2163.005 23.855 2163.295 24.085 ;
        RECT 2163.080 23.700 2163.220 23.855 ;
        RECT 2114.780 23.560 2163.220 23.700 ;
        RECT 1972.090 23.020 1972.410 23.080 ;
        RECT 2018.105 23.020 2018.395 23.065 ;
        RECT 1972.090 22.880 2018.395 23.020 ;
        RECT 1972.090 22.820 1972.410 22.880 ;
        RECT 2018.105 22.835 2018.395 22.880 ;
        RECT 2062.265 23.020 2062.555 23.065 ;
        RECT 2114.780 23.020 2114.920 23.560 ;
        RECT 2062.265 22.880 2114.920 23.020 ;
        RECT 2062.265 22.835 2062.555 22.880 ;
        RECT 2018.105 21.320 2018.395 21.365 ;
        RECT 2062.265 21.320 2062.555 21.365 ;
        RECT 2018.105 21.180 2062.555 21.320 ;
        RECT 2018.105 21.135 2018.395 21.180 ;
        RECT 2062.265 21.135 2062.555 21.180 ;
      LAYER via ;
        RECT 1875.520 1209.760 1875.780 1210.020 ;
        RECT 1970.280 1209.760 1970.540 1210.020 ;
        RECT 1968.900 1159.100 1969.160 1159.360 ;
        RECT 1969.820 1159.100 1970.080 1159.360 ;
        RECT 1969.820 158.480 1970.080 158.740 ;
        RECT 1970.740 158.480 1971.000 158.740 ;
        RECT 1970.740 144.540 1971.000 144.800 ;
        RECT 1970.280 96.600 1970.540 96.860 ;
        RECT 2191.080 24.180 2191.340 24.440 ;
        RECT 1972.120 22.820 1972.380 23.080 ;
      LAYER met2 ;
        RECT 1875.530 1219.680 1876.090 1228.680 ;
        RECT 1875.580 1210.050 1875.720 1219.680 ;
        RECT 1875.520 1209.730 1875.780 1210.050 ;
        RECT 1970.280 1209.730 1970.540 1210.050 ;
        RECT 1970.340 1207.525 1970.480 1209.730 ;
        RECT 1968.890 1207.155 1969.170 1207.525 ;
        RECT 1970.270 1207.155 1970.550 1207.525 ;
        RECT 1968.960 1159.390 1969.100 1207.155 ;
        RECT 1968.900 1159.070 1969.160 1159.390 ;
        RECT 1969.820 1159.070 1970.080 1159.390 ;
        RECT 1969.880 158.770 1970.020 1159.070 ;
        RECT 1969.820 158.450 1970.080 158.770 ;
        RECT 1970.740 158.450 1971.000 158.770 ;
        RECT 1970.800 144.830 1970.940 158.450 ;
        RECT 1970.740 144.510 1971.000 144.830 ;
        RECT 1970.280 96.570 1970.540 96.890 ;
        RECT 1970.340 62.290 1970.480 96.570 ;
        RECT 1970.340 62.150 1972.320 62.290 ;
        RECT 1972.180 23.110 1972.320 62.150 ;
        RECT 2191.080 24.150 2191.340 24.470 ;
        RECT 1972.120 22.790 1972.380 23.110 ;
        RECT 2191.140 2.400 2191.280 24.150 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
      LAYER via2 ;
        RECT 1968.890 1207.200 1969.170 1207.480 ;
        RECT 1970.270 1207.200 1970.550 1207.480 ;
      LAYER met3 ;
        RECT 1968.865 1207.490 1969.195 1207.505 ;
        RECT 1970.245 1207.490 1970.575 1207.505 ;
        RECT 1968.865 1207.190 1970.575 1207.490 ;
        RECT 1968.865 1207.175 1969.195 1207.190 ;
        RECT 1970.245 1207.175 1970.575 1207.190 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1897.645 1213.545 1897.815 1214.395 ;
        RECT 2113.845 23.885 2114.935 24.055 ;
        RECT 2113.845 23.205 2114.015 23.885 ;
        RECT 2114.765 23.715 2114.935 23.885 ;
        RECT 2116.145 23.715 2116.315 25.075 ;
        RECT 2114.765 23.545 2116.315 23.715 ;
      LAYER mcon ;
        RECT 1897.645 1214.225 1897.815 1214.395 ;
        RECT 2116.145 24.905 2116.315 25.075 ;
      LAYER met1 ;
        RECT 1897.585 1214.380 1897.875 1214.425 ;
        RECT 1990.490 1214.380 1990.810 1214.440 ;
        RECT 1897.585 1214.240 1990.810 1214.380 ;
        RECT 1897.585 1214.195 1897.875 1214.240 ;
        RECT 1990.490 1214.180 1990.810 1214.240 ;
        RECT 1897.585 1213.515 1897.875 1213.745 ;
        RECT 1884.690 1213.360 1885.010 1213.420 ;
        RECT 1897.660 1213.360 1897.800 1213.515 ;
        RECT 1884.690 1213.220 1897.800 1213.360 ;
        RECT 1884.690 1213.160 1885.010 1213.220 ;
        RECT 2116.085 25.060 2116.375 25.105 ;
        RECT 2116.085 24.920 2162.760 25.060 ;
        RECT 2116.085 24.875 2116.375 24.920 ;
        RECT 2162.620 24.380 2162.760 24.920 ;
        RECT 2162.620 24.240 2163.680 24.380 ;
        RECT 2163.540 24.040 2163.680 24.240 ;
        RECT 2208.990 24.040 2209.310 24.100 ;
        RECT 2163.540 23.900 2209.310 24.040 ;
        RECT 2208.990 23.840 2209.310 23.900 ;
        RECT 1990.490 23.360 1990.810 23.420 ;
        RECT 1994.170 23.360 1994.490 23.420 ;
        RECT 2113.785 23.360 2114.075 23.405 ;
        RECT 1990.490 23.220 1994.490 23.360 ;
        RECT 1990.490 23.160 1990.810 23.220 ;
        RECT 1994.170 23.160 1994.490 23.220 ;
        RECT 2061.880 23.220 2114.075 23.360 ;
        RECT 2018.550 23.020 2018.870 23.080 ;
        RECT 2061.880 23.020 2062.020 23.220 ;
        RECT 2113.785 23.175 2114.075 23.220 ;
        RECT 2018.550 22.880 2062.020 23.020 ;
        RECT 2018.550 22.820 2018.870 22.880 ;
        RECT 2007.050 22.680 2007.370 22.740 ;
        RECT 2017.170 22.680 2017.490 22.740 ;
        RECT 2007.050 22.540 2017.490 22.680 ;
        RECT 2007.050 22.480 2007.370 22.540 ;
        RECT 2017.170 22.480 2017.490 22.540 ;
      LAYER via ;
        RECT 1990.520 1214.180 1990.780 1214.440 ;
        RECT 1884.720 1213.160 1884.980 1213.420 ;
        RECT 2209.020 23.840 2209.280 24.100 ;
        RECT 1990.520 23.160 1990.780 23.420 ;
        RECT 1994.200 23.160 1994.460 23.420 ;
        RECT 2018.580 22.820 2018.840 23.080 ;
        RECT 2007.080 22.480 2007.340 22.740 ;
        RECT 2017.200 22.480 2017.460 22.740 ;
      LAYER met2 ;
        RECT 1884.730 1219.680 1885.290 1228.680 ;
        RECT 1884.780 1213.450 1884.920 1219.680 ;
        RECT 1990.520 1214.150 1990.780 1214.470 ;
        RECT 1884.720 1213.130 1884.980 1213.450 ;
        RECT 1990.580 23.450 1990.720 1214.150 ;
        RECT 2209.020 23.810 2209.280 24.130 ;
        RECT 1990.520 23.130 1990.780 23.450 ;
        RECT 1994.200 23.130 1994.460 23.450 ;
        RECT 1994.260 22.965 1994.400 23.130 ;
        RECT 1994.190 22.595 1994.470 22.965 ;
        RECT 2007.070 22.595 2007.350 22.965 ;
        RECT 2018.580 22.850 2018.840 23.110 ;
        RECT 2017.260 22.790 2018.840 22.850 ;
        RECT 2017.260 22.770 2018.780 22.790 ;
        RECT 2017.200 22.710 2018.780 22.770 ;
        RECT 2007.080 22.450 2007.340 22.595 ;
        RECT 2017.200 22.450 2017.460 22.710 ;
        RECT 2209.080 2.400 2209.220 23.810 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
      LAYER via2 ;
        RECT 1994.190 22.640 1994.470 22.920 ;
        RECT 2007.070 22.640 2007.350 22.920 ;
      LAYER met3 ;
        RECT 1994.165 22.930 1994.495 22.945 ;
        RECT 2007.045 22.930 2007.375 22.945 ;
        RECT 1994.165 22.630 2007.375 22.930 ;
        RECT 1994.165 22.615 1994.495 22.630 ;
        RECT 2007.045 22.615 2007.375 22.630 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1895.345 786.505 1895.515 814.215 ;
        RECT 1895.805 662.405 1895.975 710.515 ;
        RECT 1895.805 614.125 1895.975 661.895 ;
        RECT 1895.805 446.845 1895.975 500.395 ;
        RECT 1895.805 283.305 1895.975 331.075 ;
        RECT 1895.805 234.685 1895.975 282.795 ;
        RECT 1896.265 110.245 1896.435 137.615 ;
      LAYER mcon ;
        RECT 1895.345 814.045 1895.515 814.215 ;
        RECT 1895.805 710.345 1895.975 710.515 ;
        RECT 1895.805 661.725 1895.975 661.895 ;
        RECT 1895.805 500.225 1895.975 500.395 ;
        RECT 1895.805 330.905 1895.975 331.075 ;
        RECT 1895.805 282.625 1895.975 282.795 ;
        RECT 1896.265 137.445 1896.435 137.615 ;
      LAYER met1 ;
        RECT 1895.270 1104.220 1895.590 1104.280 ;
        RECT 1896.190 1104.220 1896.510 1104.280 ;
        RECT 1895.270 1104.080 1896.510 1104.220 ;
        RECT 1895.270 1104.020 1895.590 1104.080 ;
        RECT 1896.190 1104.020 1896.510 1104.080 ;
        RECT 1895.730 1103.880 1896.050 1103.940 ;
        RECT 1896.650 1103.880 1896.970 1103.940 ;
        RECT 1895.730 1103.740 1896.970 1103.880 ;
        RECT 1895.730 1103.680 1896.050 1103.740 ;
        RECT 1896.650 1103.680 1896.970 1103.740 ;
        RECT 1895.730 1055.600 1896.050 1055.660 ;
        RECT 1896.190 1055.600 1896.510 1055.660 ;
        RECT 1895.730 1055.460 1896.510 1055.600 ;
        RECT 1895.730 1055.400 1896.050 1055.460 ;
        RECT 1896.190 1055.400 1896.510 1055.460 ;
        RECT 1894.350 918.240 1894.670 918.300 ;
        RECT 1895.270 918.240 1895.590 918.300 ;
        RECT 1894.350 918.100 1895.590 918.240 ;
        RECT 1894.350 918.040 1894.670 918.100 ;
        RECT 1895.270 918.040 1895.590 918.100 ;
        RECT 1895.270 910.760 1895.590 910.820 ;
        RECT 1896.650 910.760 1896.970 910.820 ;
        RECT 1895.270 910.620 1896.970 910.760 ;
        RECT 1895.270 910.560 1895.590 910.620 ;
        RECT 1896.650 910.560 1896.970 910.620 ;
        RECT 1895.730 821.340 1896.050 821.400 ;
        RECT 1896.650 821.340 1896.970 821.400 ;
        RECT 1895.730 821.200 1896.970 821.340 ;
        RECT 1895.730 821.140 1896.050 821.200 ;
        RECT 1896.650 821.140 1896.970 821.200 ;
        RECT 1895.270 814.200 1895.590 814.260 ;
        RECT 1895.075 814.060 1895.590 814.200 ;
        RECT 1895.270 814.000 1895.590 814.060 ;
        RECT 1895.270 786.660 1895.590 786.720 ;
        RECT 1895.075 786.520 1895.590 786.660 ;
        RECT 1895.270 786.460 1895.590 786.520 ;
        RECT 1895.730 724.580 1896.050 724.840 ;
        RECT 1895.820 724.160 1895.960 724.580 ;
        RECT 1895.730 723.900 1896.050 724.160 ;
        RECT 1895.730 710.500 1896.050 710.560 ;
        RECT 1895.535 710.360 1896.050 710.500 ;
        RECT 1895.730 710.300 1896.050 710.360 ;
        RECT 1895.745 662.560 1896.035 662.605 ;
        RECT 1896.190 662.560 1896.510 662.620 ;
        RECT 1895.745 662.420 1896.510 662.560 ;
        RECT 1895.745 662.375 1896.035 662.420 ;
        RECT 1896.190 662.360 1896.510 662.420 ;
        RECT 1895.745 661.880 1896.035 661.925 ;
        RECT 1896.190 661.880 1896.510 661.940 ;
        RECT 1895.745 661.740 1896.510 661.880 ;
        RECT 1895.745 661.695 1896.035 661.740 ;
        RECT 1896.190 661.680 1896.510 661.740 ;
        RECT 1895.730 614.280 1896.050 614.340 ;
        RECT 1895.535 614.140 1896.050 614.280 ;
        RECT 1895.730 614.080 1896.050 614.140 ;
        RECT 1895.730 500.380 1896.050 500.440 ;
        RECT 1895.535 500.240 1896.050 500.380 ;
        RECT 1895.730 500.180 1896.050 500.240 ;
        RECT 1895.730 447.000 1896.050 447.060 ;
        RECT 1895.535 446.860 1896.050 447.000 ;
        RECT 1895.730 446.800 1896.050 446.860 ;
        RECT 1895.730 331.060 1896.050 331.120 ;
        RECT 1895.535 330.920 1896.050 331.060 ;
        RECT 1895.730 330.860 1896.050 330.920 ;
        RECT 1895.730 283.460 1896.050 283.520 ;
        RECT 1895.535 283.320 1896.050 283.460 ;
        RECT 1895.730 283.260 1896.050 283.320 ;
        RECT 1895.730 282.780 1896.050 282.840 ;
        RECT 1895.535 282.640 1896.050 282.780 ;
        RECT 1895.730 282.580 1896.050 282.640 ;
        RECT 1895.745 234.840 1896.035 234.885 ;
        RECT 1896.190 234.840 1896.510 234.900 ;
        RECT 1895.745 234.700 1896.510 234.840 ;
        RECT 1895.745 234.655 1896.035 234.700 ;
        RECT 1896.190 234.640 1896.510 234.700 ;
        RECT 1895.730 186.560 1896.050 186.620 ;
        RECT 1896.190 186.560 1896.510 186.620 ;
        RECT 1895.730 186.420 1896.510 186.560 ;
        RECT 1895.730 186.360 1896.050 186.420 ;
        RECT 1896.190 186.360 1896.510 186.420 ;
        RECT 1896.650 159.020 1896.970 159.080 ;
        RECT 1896.280 158.880 1896.970 159.020 ;
        RECT 1896.280 158.400 1896.420 158.880 ;
        RECT 1896.650 158.820 1896.970 158.880 ;
        RECT 1896.190 158.140 1896.510 158.400 ;
        RECT 1896.190 137.600 1896.510 137.660 ;
        RECT 1895.995 137.460 1896.510 137.600 ;
        RECT 1896.190 137.400 1896.510 137.460 ;
        RECT 1896.205 110.400 1896.495 110.445 ;
        RECT 1896.650 110.400 1896.970 110.460 ;
        RECT 1896.205 110.260 1896.970 110.400 ;
        RECT 1896.205 110.215 1896.495 110.260 ;
        RECT 1896.650 110.200 1896.970 110.260 ;
        RECT 1896.190 34.920 1896.510 34.980 ;
        RECT 2226.930 34.920 2227.250 34.980 ;
        RECT 1896.190 34.780 2227.250 34.920 ;
        RECT 1896.190 34.720 1896.510 34.780 ;
        RECT 2226.930 34.720 2227.250 34.780 ;
      LAYER via ;
        RECT 1895.300 1104.020 1895.560 1104.280 ;
        RECT 1896.220 1104.020 1896.480 1104.280 ;
        RECT 1895.760 1103.680 1896.020 1103.940 ;
        RECT 1896.680 1103.680 1896.940 1103.940 ;
        RECT 1895.760 1055.400 1896.020 1055.660 ;
        RECT 1896.220 1055.400 1896.480 1055.660 ;
        RECT 1894.380 918.040 1894.640 918.300 ;
        RECT 1895.300 918.040 1895.560 918.300 ;
        RECT 1895.300 910.560 1895.560 910.820 ;
        RECT 1896.680 910.560 1896.940 910.820 ;
        RECT 1895.760 821.140 1896.020 821.400 ;
        RECT 1896.680 821.140 1896.940 821.400 ;
        RECT 1895.300 814.000 1895.560 814.260 ;
        RECT 1895.300 786.460 1895.560 786.720 ;
        RECT 1895.760 724.580 1896.020 724.840 ;
        RECT 1895.760 723.900 1896.020 724.160 ;
        RECT 1895.760 710.300 1896.020 710.560 ;
        RECT 1896.220 662.360 1896.480 662.620 ;
        RECT 1896.220 661.680 1896.480 661.940 ;
        RECT 1895.760 614.080 1896.020 614.340 ;
        RECT 1895.760 500.180 1896.020 500.440 ;
        RECT 1895.760 446.800 1896.020 447.060 ;
        RECT 1895.760 330.860 1896.020 331.120 ;
        RECT 1895.760 283.260 1896.020 283.520 ;
        RECT 1895.760 282.580 1896.020 282.840 ;
        RECT 1896.220 234.640 1896.480 234.900 ;
        RECT 1895.760 186.360 1896.020 186.620 ;
        RECT 1896.220 186.360 1896.480 186.620 ;
        RECT 1896.680 158.820 1896.940 159.080 ;
        RECT 1896.220 158.140 1896.480 158.400 ;
        RECT 1896.220 137.400 1896.480 137.660 ;
        RECT 1896.680 110.200 1896.940 110.460 ;
        RECT 1896.220 34.720 1896.480 34.980 ;
        RECT 2226.960 34.720 2227.220 34.980 ;
      LAYER met2 ;
        RECT 1893.470 1220.330 1894.030 1228.680 ;
        RECT 1893.470 1220.190 1895.040 1220.330 ;
        RECT 1893.470 1219.680 1894.030 1220.190 ;
        RECT 1894.900 1177.490 1895.040 1220.190 ;
        RECT 1894.440 1177.350 1895.040 1177.490 ;
        RECT 1894.440 1153.805 1894.580 1177.350 ;
        RECT 1894.370 1153.435 1894.650 1153.805 ;
        RECT 1896.210 1152.075 1896.490 1152.445 ;
        RECT 1895.360 1104.310 1895.500 1104.465 ;
        RECT 1896.280 1104.310 1896.420 1152.075 ;
        RECT 1895.300 1104.050 1895.560 1104.310 ;
        RECT 1895.300 1103.990 1895.960 1104.050 ;
        RECT 1896.220 1103.990 1896.480 1104.310 ;
        RECT 1895.360 1103.970 1895.960 1103.990 ;
        RECT 1895.360 1103.910 1896.020 1103.970 ;
        RECT 1895.760 1103.650 1896.020 1103.910 ;
        RECT 1896.680 1103.650 1896.940 1103.970 ;
        RECT 1896.740 1055.770 1896.880 1103.650 ;
        RECT 1895.820 1055.690 1896.880 1055.770 ;
        RECT 1895.760 1055.630 1896.880 1055.690 ;
        RECT 1895.760 1055.370 1896.020 1055.630 ;
        RECT 1896.220 1055.370 1896.480 1055.630 ;
        RECT 1895.820 1055.215 1895.960 1055.370 ;
        RECT 1896.280 1007.605 1896.420 1055.370 ;
        RECT 1895.290 1007.235 1895.570 1007.605 ;
        RECT 1896.210 1007.235 1896.490 1007.605 ;
        RECT 1895.360 966.010 1895.500 1007.235 ;
        RECT 1894.440 965.870 1895.500 966.010 ;
        RECT 1894.440 918.330 1894.580 965.870 ;
        RECT 1894.380 918.010 1894.640 918.330 ;
        RECT 1895.300 918.010 1895.560 918.330 ;
        RECT 1895.360 910.850 1895.500 918.010 ;
        RECT 1895.300 910.530 1895.560 910.850 ;
        RECT 1896.680 910.530 1896.940 910.850 ;
        RECT 1896.740 821.430 1896.880 910.530 ;
        RECT 1895.760 821.170 1896.020 821.430 ;
        RECT 1895.360 821.110 1896.020 821.170 ;
        RECT 1896.680 821.110 1896.940 821.430 ;
        RECT 1895.360 821.030 1895.960 821.110 ;
        RECT 1895.360 814.290 1895.500 821.030 ;
        RECT 1895.300 813.970 1895.560 814.290 ;
        RECT 1895.300 786.430 1895.560 786.750 ;
        RECT 1895.360 766.090 1895.500 786.430 ;
        RECT 1895.360 765.950 1895.960 766.090 ;
        RECT 1895.820 724.870 1895.960 765.950 ;
        RECT 1895.760 724.550 1896.020 724.870 ;
        RECT 1895.760 723.870 1896.020 724.190 ;
        RECT 1895.820 710.590 1895.960 723.870 ;
        RECT 1895.760 710.270 1896.020 710.590 ;
        RECT 1896.220 662.330 1896.480 662.650 ;
        RECT 1896.280 661.970 1896.420 662.330 ;
        RECT 1896.220 661.650 1896.480 661.970 ;
        RECT 1895.760 614.050 1896.020 614.370 ;
        RECT 1895.820 500.470 1895.960 614.050 ;
        RECT 1895.760 500.150 1896.020 500.470 ;
        RECT 1895.760 446.770 1896.020 447.090 ;
        RECT 1895.820 331.150 1895.960 446.770 ;
        RECT 1895.760 330.830 1896.020 331.150 ;
        RECT 1895.760 283.230 1896.020 283.550 ;
        RECT 1895.820 282.870 1895.960 283.230 ;
        RECT 1895.760 282.550 1896.020 282.870 ;
        RECT 1896.220 234.610 1896.480 234.930 ;
        RECT 1896.280 186.650 1896.420 234.610 ;
        RECT 1895.760 186.330 1896.020 186.650 ;
        RECT 1896.220 186.330 1896.480 186.650 ;
        RECT 1895.820 186.165 1895.960 186.330 ;
        RECT 1895.750 185.795 1896.030 186.165 ;
        RECT 1896.670 185.795 1896.950 186.165 ;
        RECT 1896.740 159.110 1896.880 185.795 ;
        RECT 1896.680 158.790 1896.940 159.110 ;
        RECT 1896.220 158.110 1896.480 158.430 ;
        RECT 1896.280 137.690 1896.420 158.110 ;
        RECT 1896.220 137.370 1896.480 137.690 ;
        RECT 1896.680 110.170 1896.940 110.490 ;
        RECT 1896.740 72.490 1896.880 110.170 ;
        RECT 1896.280 72.350 1896.880 72.490 ;
        RECT 1896.280 35.010 1896.420 72.350 ;
        RECT 1896.220 34.690 1896.480 35.010 ;
        RECT 2226.960 34.690 2227.220 35.010 ;
        RECT 2227.020 2.400 2227.160 34.690 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
      LAYER via2 ;
        RECT 1894.370 1153.480 1894.650 1153.760 ;
        RECT 1896.210 1152.120 1896.490 1152.400 ;
        RECT 1895.290 1007.280 1895.570 1007.560 ;
        RECT 1896.210 1007.280 1896.490 1007.560 ;
        RECT 1895.750 185.840 1896.030 186.120 ;
        RECT 1896.670 185.840 1896.950 186.120 ;
      LAYER met3 ;
        RECT 1894.345 1153.770 1894.675 1153.785 ;
        RECT 1894.345 1153.470 1896.730 1153.770 ;
        RECT 1894.345 1153.455 1894.675 1153.470 ;
        RECT 1896.430 1152.425 1896.730 1153.470 ;
        RECT 1896.185 1152.110 1896.730 1152.425 ;
        RECT 1896.185 1152.095 1896.515 1152.110 ;
        RECT 1895.265 1007.570 1895.595 1007.585 ;
        RECT 1896.185 1007.570 1896.515 1007.585 ;
        RECT 1895.265 1007.270 1896.515 1007.570 ;
        RECT 1895.265 1007.255 1895.595 1007.270 ;
        RECT 1896.185 1007.255 1896.515 1007.270 ;
        RECT 1895.725 186.130 1896.055 186.145 ;
        RECT 1896.645 186.130 1896.975 186.145 ;
        RECT 1895.725 185.830 1896.975 186.130 ;
        RECT 1895.725 185.815 1896.055 185.830 ;
        RECT 1896.645 185.815 1896.975 185.830 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1146.850 1159.300 1147.170 1159.360 ;
        RECT 1149.150 1159.300 1149.470 1159.360 ;
        RECT 1146.850 1159.160 1149.470 1159.300 ;
        RECT 1146.850 1159.100 1147.170 1159.160 ;
        RECT 1149.150 1159.100 1149.470 1159.160 ;
        RECT 1146.390 1014.460 1146.710 1014.520 ;
        RECT 1146.850 1014.460 1147.170 1014.520 ;
        RECT 1146.390 1014.320 1147.170 1014.460 ;
        RECT 1146.390 1014.260 1146.710 1014.320 ;
        RECT 1146.850 1014.260 1147.170 1014.320 ;
        RECT 1146.850 1007.320 1147.170 1007.380 ;
        RECT 1147.310 1007.320 1147.630 1007.380 ;
        RECT 1146.850 1007.180 1147.630 1007.320 ;
        RECT 1146.850 1007.120 1147.170 1007.180 ;
        RECT 1147.310 1007.120 1147.630 1007.180 ;
        RECT 1146.390 869.620 1146.710 869.680 ;
        RECT 1147.310 869.620 1147.630 869.680 ;
        RECT 1146.390 869.480 1147.630 869.620 ;
        RECT 1146.390 869.420 1146.710 869.480 ;
        RECT 1147.310 869.420 1147.630 869.480 ;
        RECT 1145.930 773.060 1146.250 773.120 ;
        RECT 1146.390 773.060 1146.710 773.120 ;
        RECT 1145.930 772.920 1146.710 773.060 ;
        RECT 1145.930 772.860 1146.250 772.920 ;
        RECT 1146.390 772.860 1146.710 772.920 ;
        RECT 1145.930 435.100 1146.250 435.160 ;
        RECT 1146.390 435.100 1146.710 435.160 ;
        RECT 1145.930 434.960 1146.710 435.100 ;
        RECT 1145.930 434.900 1146.250 434.960 ;
        RECT 1146.390 434.900 1146.710 434.960 ;
        RECT 1145.930 427.420 1146.250 427.680 ;
        RECT 1146.020 427.280 1146.160 427.420 ;
        RECT 1146.850 427.280 1147.170 427.340 ;
        RECT 1146.020 427.140 1147.170 427.280 ;
        RECT 1146.850 427.080 1147.170 427.140 ;
        RECT 1146.390 289.920 1146.710 289.980 ;
        RECT 1146.850 289.920 1147.170 289.980 ;
        RECT 1146.390 289.780 1147.170 289.920 ;
        RECT 1146.390 289.720 1146.710 289.780 ;
        RECT 1146.850 289.720 1147.170 289.780 ;
        RECT 1146.850 145.080 1147.170 145.140 ;
        RECT 1147.310 145.080 1147.630 145.140 ;
        RECT 1146.850 144.940 1147.630 145.080 ;
        RECT 1146.850 144.880 1147.170 144.940 ;
        RECT 1147.310 144.880 1147.630 144.940 ;
        RECT 1146.390 96.800 1146.710 96.860 ;
        RECT 1146.850 96.800 1147.170 96.860 ;
        RECT 1146.390 96.660 1147.170 96.800 ;
        RECT 1146.390 96.600 1146.710 96.660 ;
        RECT 1146.850 96.600 1147.170 96.660 ;
        RECT 781.610 41.720 781.930 41.780 ;
        RECT 1146.390 41.720 1146.710 41.780 ;
        RECT 781.610 41.580 1146.710 41.720 ;
        RECT 781.610 41.520 781.930 41.580 ;
        RECT 1146.390 41.520 1146.710 41.580 ;
      LAYER via ;
        RECT 1146.880 1159.100 1147.140 1159.360 ;
        RECT 1149.180 1159.100 1149.440 1159.360 ;
        RECT 1146.420 1014.260 1146.680 1014.520 ;
        RECT 1146.880 1014.260 1147.140 1014.520 ;
        RECT 1146.880 1007.120 1147.140 1007.380 ;
        RECT 1147.340 1007.120 1147.600 1007.380 ;
        RECT 1146.420 869.420 1146.680 869.680 ;
        RECT 1147.340 869.420 1147.600 869.680 ;
        RECT 1145.960 772.860 1146.220 773.120 ;
        RECT 1146.420 772.860 1146.680 773.120 ;
        RECT 1145.960 434.900 1146.220 435.160 ;
        RECT 1146.420 434.900 1146.680 435.160 ;
        RECT 1145.960 427.420 1146.220 427.680 ;
        RECT 1146.880 427.080 1147.140 427.340 ;
        RECT 1146.420 289.720 1146.680 289.980 ;
        RECT 1146.880 289.720 1147.140 289.980 ;
        RECT 1146.880 144.880 1147.140 145.140 ;
        RECT 1147.340 144.880 1147.600 145.140 ;
        RECT 1146.420 96.600 1146.680 96.860 ;
        RECT 1146.880 96.600 1147.140 96.860 ;
        RECT 781.640 41.520 781.900 41.780 ;
        RECT 1146.420 41.520 1146.680 41.780 ;
      LAYER met2 ;
        RECT 1151.490 1221.010 1152.050 1228.680 ;
        RECT 1149.240 1220.870 1152.050 1221.010 ;
        RECT 1149.240 1159.390 1149.380 1220.870 ;
        RECT 1151.490 1219.680 1152.050 1220.870 ;
        RECT 1146.880 1159.070 1147.140 1159.390 ;
        RECT 1149.180 1159.070 1149.440 1159.390 ;
        RECT 1146.940 1076.850 1147.080 1159.070 ;
        RECT 1146.480 1076.710 1147.080 1076.850 ;
        RECT 1146.480 1014.550 1146.620 1076.710 ;
        RECT 1146.420 1014.230 1146.680 1014.550 ;
        RECT 1146.880 1014.230 1147.140 1014.550 ;
        RECT 1146.940 1007.410 1147.080 1014.230 ;
        RECT 1146.880 1007.090 1147.140 1007.410 ;
        RECT 1147.340 1007.090 1147.600 1007.410 ;
        RECT 1147.400 869.710 1147.540 1007.090 ;
        RECT 1146.420 869.390 1146.680 869.710 ;
        RECT 1147.340 869.390 1147.600 869.710 ;
        RECT 1146.480 787.850 1146.620 869.390 ;
        RECT 1146.020 787.710 1146.620 787.850 ;
        RECT 1146.020 773.150 1146.160 787.710 ;
        RECT 1145.960 772.830 1146.220 773.150 ;
        RECT 1146.420 772.830 1146.680 773.150 ;
        RECT 1146.480 748.410 1146.620 772.830 ;
        RECT 1146.480 748.270 1147.540 748.410 ;
        RECT 1147.400 676.445 1147.540 748.270 ;
        RECT 1146.410 676.075 1146.690 676.445 ;
        RECT 1147.330 676.075 1147.610 676.445 ;
        RECT 1146.480 628.050 1146.620 676.075 ;
        RECT 1146.480 627.910 1147.080 628.050 ;
        RECT 1146.940 507.010 1147.080 627.910 ;
        RECT 1146.480 506.870 1147.080 507.010 ;
        RECT 1146.480 435.190 1146.620 506.870 ;
        RECT 1145.960 434.870 1146.220 435.190 ;
        RECT 1146.420 434.870 1146.680 435.190 ;
        RECT 1146.020 427.710 1146.160 434.870 ;
        RECT 1145.960 427.390 1146.220 427.710 ;
        RECT 1146.880 427.050 1147.140 427.370 ;
        RECT 1146.940 290.010 1147.080 427.050 ;
        RECT 1146.420 289.690 1146.680 290.010 ;
        RECT 1146.880 289.690 1147.140 290.010 ;
        RECT 1146.480 266.290 1146.620 289.690 ;
        RECT 1146.480 266.150 1147.540 266.290 ;
        RECT 1147.400 198.970 1147.540 266.150 ;
        RECT 1146.940 198.830 1147.540 198.970 ;
        RECT 1146.940 193.020 1147.080 198.830 ;
        RECT 1146.940 192.880 1147.540 193.020 ;
        RECT 1147.400 145.170 1147.540 192.880 ;
        RECT 1146.880 144.850 1147.140 145.170 ;
        RECT 1147.340 144.850 1147.600 145.170 ;
        RECT 1146.940 96.890 1147.080 144.850 ;
        RECT 1146.420 96.570 1146.680 96.890 ;
        RECT 1146.880 96.570 1147.140 96.890 ;
        RECT 1146.480 41.810 1146.620 96.570 ;
        RECT 781.640 41.490 781.900 41.810 ;
        RECT 1146.420 41.490 1146.680 41.810 ;
        RECT 781.700 2.400 781.840 41.490 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 1146.410 676.120 1146.690 676.400 ;
        RECT 1147.330 676.120 1147.610 676.400 ;
      LAYER met3 ;
        RECT 1146.385 676.410 1146.715 676.425 ;
        RECT 1147.305 676.410 1147.635 676.425 ;
        RECT 1146.385 676.110 1147.635 676.410 ;
        RECT 1146.385 676.095 1146.715 676.110 ;
        RECT 1147.305 676.095 1147.635 676.110 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1903.550 47.160 1903.870 47.220 ;
        RECT 2244.870 47.160 2245.190 47.220 ;
        RECT 1903.550 47.020 2245.190 47.160 ;
        RECT 1903.550 46.960 1903.870 47.020 ;
        RECT 2244.870 46.960 2245.190 47.020 ;
      LAYER via ;
        RECT 1903.580 46.960 1903.840 47.220 ;
        RECT 2244.900 46.960 2245.160 47.220 ;
      LAYER met2 ;
        RECT 1902.670 1220.330 1903.230 1228.680 ;
        RECT 1902.670 1220.190 1903.780 1220.330 ;
        RECT 1902.670 1219.680 1903.230 1220.190 ;
        RECT 1903.640 47.250 1903.780 1220.190 ;
        RECT 1903.580 46.930 1903.840 47.250 ;
        RECT 2244.900 46.930 2245.160 47.250 ;
        RECT 2244.960 2.400 2245.100 46.930 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1911.830 1207.580 1912.150 1207.640 ;
        RECT 1917.810 1207.580 1918.130 1207.640 ;
        RECT 1911.830 1207.440 1918.130 1207.580 ;
        RECT 1911.830 1207.380 1912.150 1207.440 ;
        RECT 1917.810 1207.380 1918.130 1207.440 ;
        RECT 1917.810 47.500 1918.130 47.560 ;
        RECT 2262.350 47.500 2262.670 47.560 ;
        RECT 1917.810 47.360 2262.670 47.500 ;
        RECT 1917.810 47.300 1918.130 47.360 ;
        RECT 2262.350 47.300 2262.670 47.360 ;
      LAYER via ;
        RECT 1911.860 1207.380 1912.120 1207.640 ;
        RECT 1917.840 1207.380 1918.100 1207.640 ;
        RECT 1917.840 47.300 1918.100 47.560 ;
        RECT 2262.380 47.300 2262.640 47.560 ;
      LAYER met2 ;
        RECT 1911.870 1219.680 1912.430 1228.680 ;
        RECT 1911.920 1207.670 1912.060 1219.680 ;
        RECT 1911.860 1207.350 1912.120 1207.670 ;
        RECT 1917.840 1207.350 1918.100 1207.670 ;
        RECT 1917.900 47.590 1918.040 1207.350 ;
        RECT 1917.840 47.270 1918.100 47.590 ;
        RECT 2262.380 47.270 2262.640 47.590 ;
        RECT 2262.440 2.400 2262.580 47.270 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1923.405 1027.905 1923.575 1055.615 ;
        RECT 1922.945 883.065 1923.115 910.775 ;
        RECT 1922.945 766.105 1923.115 814.215 ;
        RECT 1923.405 638.945 1923.575 669.375 ;
        RECT 1922.945 524.365 1923.115 572.135 ;
        RECT 1923.405 331.245 1923.575 379.355 ;
        RECT 1922.945 89.845 1923.115 137.955 ;
      LAYER mcon ;
        RECT 1923.405 1055.445 1923.575 1055.615 ;
        RECT 1922.945 910.605 1923.115 910.775 ;
        RECT 1922.945 814.045 1923.115 814.215 ;
        RECT 1923.405 669.205 1923.575 669.375 ;
        RECT 1922.945 571.965 1923.115 572.135 ;
        RECT 1923.405 379.185 1923.575 379.355 ;
        RECT 1922.945 137.785 1923.115 137.955 ;
      LAYER met1 ;
        RECT 1922.870 1104.220 1923.190 1104.280 ;
        RECT 1924.250 1104.220 1924.570 1104.280 ;
        RECT 1922.870 1104.080 1924.570 1104.220 ;
        RECT 1922.870 1104.020 1923.190 1104.080 ;
        RECT 1924.250 1104.020 1924.570 1104.080 ;
        RECT 1923.330 1055.600 1923.650 1055.660 ;
        RECT 1923.135 1055.460 1923.650 1055.600 ;
        RECT 1923.330 1055.400 1923.650 1055.460 ;
        RECT 1923.330 1028.060 1923.650 1028.120 ;
        RECT 1923.135 1027.920 1923.650 1028.060 ;
        RECT 1923.330 1027.860 1923.650 1027.920 ;
        RECT 1922.870 918.240 1923.190 918.300 ;
        RECT 1923.330 918.240 1923.650 918.300 ;
        RECT 1922.870 918.100 1923.650 918.240 ;
        RECT 1922.870 918.040 1923.190 918.100 ;
        RECT 1923.330 918.040 1923.650 918.100 ;
        RECT 1922.870 910.760 1923.190 910.820 ;
        RECT 1922.675 910.620 1923.190 910.760 ;
        RECT 1922.870 910.560 1923.190 910.620 ;
        RECT 1922.870 883.220 1923.190 883.280 ;
        RECT 1922.675 883.080 1923.190 883.220 ;
        RECT 1922.870 883.020 1923.190 883.080 ;
        RECT 1922.870 814.200 1923.190 814.260 ;
        RECT 1922.675 814.060 1923.190 814.200 ;
        RECT 1922.870 814.000 1923.190 814.060 ;
        RECT 1922.870 766.260 1923.190 766.320 ;
        RECT 1922.675 766.120 1923.190 766.260 ;
        RECT 1922.870 766.060 1923.190 766.120 ;
        RECT 1922.870 724.100 1923.190 724.160 ;
        RECT 1924.250 724.100 1924.570 724.160 ;
        RECT 1922.870 723.960 1924.570 724.100 ;
        RECT 1922.870 723.900 1923.190 723.960 ;
        RECT 1924.250 723.900 1924.570 723.960 ;
        RECT 1923.330 669.360 1923.650 669.420 ;
        RECT 1923.135 669.220 1923.650 669.360 ;
        RECT 1923.330 669.160 1923.650 669.220 ;
        RECT 1923.330 639.100 1923.650 639.160 ;
        RECT 1923.135 638.960 1923.650 639.100 ;
        RECT 1923.330 638.900 1923.650 638.960 ;
        RECT 1922.870 572.800 1923.190 572.860 ;
        RECT 1923.330 572.800 1923.650 572.860 ;
        RECT 1922.870 572.660 1923.650 572.800 ;
        RECT 1922.870 572.600 1923.190 572.660 ;
        RECT 1923.330 572.600 1923.650 572.660 ;
        RECT 1922.870 572.120 1923.190 572.180 ;
        RECT 1922.675 571.980 1923.190 572.120 ;
        RECT 1922.870 571.920 1923.190 571.980 ;
        RECT 1922.885 524.520 1923.175 524.565 ;
        RECT 1924.250 524.520 1924.570 524.580 ;
        RECT 1922.885 524.380 1924.570 524.520 ;
        RECT 1922.885 524.335 1923.175 524.380 ;
        RECT 1924.250 524.320 1924.570 524.380 ;
        RECT 1923.330 483.040 1923.650 483.100 ;
        RECT 1924.250 483.040 1924.570 483.100 ;
        RECT 1923.330 482.900 1924.570 483.040 ;
        RECT 1923.330 482.840 1923.650 482.900 ;
        RECT 1924.250 482.840 1924.570 482.900 ;
        RECT 1923.330 379.340 1923.650 379.400 ;
        RECT 1923.135 379.200 1923.650 379.340 ;
        RECT 1923.330 379.140 1923.650 379.200 ;
        RECT 1923.345 331.400 1923.635 331.445 ;
        RECT 1923.790 331.400 1924.110 331.460 ;
        RECT 1923.345 331.260 1924.110 331.400 ;
        RECT 1923.345 331.215 1923.635 331.260 ;
        RECT 1923.790 331.200 1924.110 331.260 ;
        RECT 1923.790 241.640 1924.110 241.700 ;
        RECT 1924.250 241.640 1924.570 241.700 ;
        RECT 1923.790 241.500 1924.570 241.640 ;
        RECT 1923.790 241.440 1924.110 241.500 ;
        RECT 1924.250 241.440 1924.570 241.500 ;
        RECT 1923.330 193.360 1923.650 193.420 ;
        RECT 1923.790 193.360 1924.110 193.420 ;
        RECT 1923.330 193.220 1924.110 193.360 ;
        RECT 1923.330 193.160 1923.650 193.220 ;
        RECT 1923.790 193.160 1924.110 193.220 ;
        RECT 1923.330 158.680 1923.650 158.740 ;
        RECT 1924.250 158.680 1924.570 158.740 ;
        RECT 1923.330 158.540 1924.570 158.680 ;
        RECT 1923.330 158.480 1923.650 158.540 ;
        RECT 1924.250 158.480 1924.570 158.540 ;
        RECT 1922.885 137.940 1923.175 137.985 ;
        RECT 1924.250 137.940 1924.570 138.000 ;
        RECT 1922.885 137.800 1924.570 137.940 ;
        RECT 1922.885 137.755 1923.175 137.800 ;
        RECT 1924.250 137.740 1924.570 137.800 ;
        RECT 1922.870 90.000 1923.190 90.060 ;
        RECT 1922.675 89.860 1923.190 90.000 ;
        RECT 1922.870 89.800 1923.190 89.860 ;
        RECT 1922.870 48.520 1923.190 48.580 ;
        RECT 1924.250 48.520 1924.570 48.580 ;
        RECT 1922.870 48.380 1924.570 48.520 ;
        RECT 1922.870 48.320 1923.190 48.380 ;
        RECT 1924.250 48.320 1924.570 48.380 ;
        RECT 1924.250 46.820 1924.570 46.880 ;
        RECT 2280.290 46.820 2280.610 46.880 ;
        RECT 1924.250 46.680 2280.610 46.820 ;
        RECT 1924.250 46.620 1924.570 46.680 ;
        RECT 2280.290 46.620 2280.610 46.680 ;
      LAYER via ;
        RECT 1922.900 1104.020 1923.160 1104.280 ;
        RECT 1924.280 1104.020 1924.540 1104.280 ;
        RECT 1923.360 1055.400 1923.620 1055.660 ;
        RECT 1923.360 1027.860 1923.620 1028.120 ;
        RECT 1922.900 918.040 1923.160 918.300 ;
        RECT 1923.360 918.040 1923.620 918.300 ;
        RECT 1922.900 910.560 1923.160 910.820 ;
        RECT 1922.900 883.020 1923.160 883.280 ;
        RECT 1922.900 814.000 1923.160 814.260 ;
        RECT 1922.900 766.060 1923.160 766.320 ;
        RECT 1922.900 723.900 1923.160 724.160 ;
        RECT 1924.280 723.900 1924.540 724.160 ;
        RECT 1923.360 669.160 1923.620 669.420 ;
        RECT 1923.360 638.900 1923.620 639.160 ;
        RECT 1922.900 572.600 1923.160 572.860 ;
        RECT 1923.360 572.600 1923.620 572.860 ;
        RECT 1922.900 571.920 1923.160 572.180 ;
        RECT 1924.280 524.320 1924.540 524.580 ;
        RECT 1923.360 482.840 1923.620 483.100 ;
        RECT 1924.280 482.840 1924.540 483.100 ;
        RECT 1923.360 379.140 1923.620 379.400 ;
        RECT 1923.820 331.200 1924.080 331.460 ;
        RECT 1923.820 241.440 1924.080 241.700 ;
        RECT 1924.280 241.440 1924.540 241.700 ;
        RECT 1923.360 193.160 1923.620 193.420 ;
        RECT 1923.820 193.160 1924.080 193.420 ;
        RECT 1923.360 158.480 1923.620 158.740 ;
        RECT 1924.280 158.480 1924.540 158.740 ;
        RECT 1924.280 137.740 1924.540 138.000 ;
        RECT 1922.900 89.800 1923.160 90.060 ;
        RECT 1922.900 48.320 1923.160 48.580 ;
        RECT 1924.280 48.320 1924.540 48.580 ;
        RECT 1924.280 46.620 1924.540 46.880 ;
        RECT 2280.320 46.620 2280.580 46.880 ;
      LAYER met2 ;
        RECT 1921.070 1220.330 1921.630 1228.680 ;
        RECT 1921.070 1220.190 1923.100 1220.330 ;
        RECT 1921.070 1219.680 1921.630 1220.190 ;
        RECT 1922.960 1186.330 1923.100 1220.190 ;
        RECT 1922.960 1186.190 1923.560 1186.330 ;
        RECT 1923.420 1152.445 1923.560 1186.190 ;
        RECT 1923.350 1152.075 1923.630 1152.445 ;
        RECT 1924.270 1152.075 1924.550 1152.445 ;
        RECT 1922.960 1104.310 1923.100 1104.465 ;
        RECT 1924.340 1104.310 1924.480 1152.075 ;
        RECT 1922.900 1104.050 1923.160 1104.310 ;
        RECT 1922.900 1103.990 1923.560 1104.050 ;
        RECT 1924.280 1103.990 1924.540 1104.310 ;
        RECT 1922.960 1103.910 1923.560 1103.990 ;
        RECT 1923.420 1103.370 1923.560 1103.910 ;
        RECT 1922.960 1103.230 1923.560 1103.370 ;
        RECT 1922.960 1055.770 1923.100 1103.230 ;
        RECT 1922.960 1055.690 1923.560 1055.770 ;
        RECT 1922.960 1055.630 1923.620 1055.690 ;
        RECT 1923.360 1055.370 1923.620 1055.630 ;
        RECT 1923.420 1055.215 1923.560 1055.370 ;
        RECT 1923.360 1027.830 1923.620 1028.150 ;
        RECT 1923.420 918.330 1923.560 1027.830 ;
        RECT 1922.900 918.010 1923.160 918.330 ;
        RECT 1923.360 918.010 1923.620 918.330 ;
        RECT 1922.960 910.850 1923.100 918.010 ;
        RECT 1922.900 910.530 1923.160 910.850 ;
        RECT 1922.900 882.990 1923.160 883.310 ;
        RECT 1922.960 821.850 1923.100 882.990 ;
        RECT 1922.960 821.710 1923.560 821.850 ;
        RECT 1923.420 821.170 1923.560 821.710 ;
        RECT 1922.960 821.030 1923.560 821.170 ;
        RECT 1922.960 814.290 1923.100 821.030 ;
        RECT 1922.900 813.970 1923.160 814.290 ;
        RECT 1922.900 766.030 1923.160 766.350 ;
        RECT 1922.960 724.190 1923.100 766.030 ;
        RECT 1922.900 723.870 1923.160 724.190 ;
        RECT 1924.280 723.870 1924.540 724.190 ;
        RECT 1924.340 676.445 1924.480 723.870 ;
        RECT 1923.350 676.075 1923.630 676.445 ;
        RECT 1924.270 676.075 1924.550 676.445 ;
        RECT 1923.420 669.450 1923.560 676.075 ;
        RECT 1923.360 669.130 1923.620 669.450 ;
        RECT 1923.360 638.870 1923.620 639.190 ;
        RECT 1923.420 572.890 1923.560 638.870 ;
        RECT 1922.900 572.570 1923.160 572.890 ;
        RECT 1923.360 572.570 1923.620 572.890 ;
        RECT 1922.960 572.210 1923.100 572.570 ;
        RECT 1922.900 571.890 1923.160 572.210 ;
        RECT 1924.280 524.290 1924.540 524.610 ;
        RECT 1924.340 483.325 1924.480 524.290 ;
        RECT 1923.350 482.955 1923.630 483.325 ;
        RECT 1924.270 482.955 1924.550 483.325 ;
        RECT 1923.360 482.810 1923.620 482.955 ;
        RECT 1924.280 482.810 1924.540 482.955 ;
        RECT 1924.340 435.045 1924.480 482.810 ;
        RECT 1923.350 434.675 1923.630 435.045 ;
        RECT 1924.270 434.675 1924.550 435.045 ;
        RECT 1923.420 379.430 1923.560 434.675 ;
        RECT 1923.360 379.110 1923.620 379.430 ;
        RECT 1923.820 331.170 1924.080 331.490 ;
        RECT 1923.880 307.090 1924.020 331.170 ;
        RECT 1923.880 306.950 1924.480 307.090 ;
        RECT 1924.340 241.730 1924.480 306.950 ;
        RECT 1923.820 241.410 1924.080 241.730 ;
        RECT 1924.280 241.410 1924.540 241.730 ;
        RECT 1923.880 193.450 1924.020 241.410 ;
        RECT 1923.360 193.130 1923.620 193.450 ;
        RECT 1923.820 193.130 1924.080 193.450 ;
        RECT 1923.420 158.770 1923.560 193.130 ;
        RECT 1923.360 158.450 1923.620 158.770 ;
        RECT 1924.280 158.450 1924.540 158.770 ;
        RECT 1924.340 138.030 1924.480 158.450 ;
        RECT 1924.280 137.710 1924.540 138.030 ;
        RECT 1922.900 89.770 1923.160 90.090 ;
        RECT 1922.960 48.610 1923.100 89.770 ;
        RECT 1922.900 48.290 1923.160 48.610 ;
        RECT 1924.280 48.290 1924.540 48.610 ;
        RECT 1924.340 46.910 1924.480 48.290 ;
        RECT 1924.280 46.590 1924.540 46.910 ;
        RECT 2280.320 46.590 2280.580 46.910 ;
        RECT 2280.380 2.400 2280.520 46.590 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
      LAYER via2 ;
        RECT 1923.350 1152.120 1923.630 1152.400 ;
        RECT 1924.270 1152.120 1924.550 1152.400 ;
        RECT 1923.350 676.120 1923.630 676.400 ;
        RECT 1924.270 676.120 1924.550 676.400 ;
        RECT 1923.350 483.000 1923.630 483.280 ;
        RECT 1924.270 483.000 1924.550 483.280 ;
        RECT 1923.350 434.720 1923.630 435.000 ;
        RECT 1924.270 434.720 1924.550 435.000 ;
      LAYER met3 ;
        RECT 1923.325 1152.410 1923.655 1152.425 ;
        RECT 1924.245 1152.410 1924.575 1152.425 ;
        RECT 1923.325 1152.110 1924.575 1152.410 ;
        RECT 1923.325 1152.095 1923.655 1152.110 ;
        RECT 1924.245 1152.095 1924.575 1152.110 ;
        RECT 1923.325 676.410 1923.655 676.425 ;
        RECT 1924.245 676.410 1924.575 676.425 ;
        RECT 1923.325 676.110 1924.575 676.410 ;
        RECT 1923.325 676.095 1923.655 676.110 ;
        RECT 1924.245 676.095 1924.575 676.110 ;
        RECT 1923.325 483.290 1923.655 483.305 ;
        RECT 1924.245 483.290 1924.575 483.305 ;
        RECT 1923.325 482.990 1924.575 483.290 ;
        RECT 1923.325 482.975 1923.655 482.990 ;
        RECT 1924.245 482.975 1924.575 482.990 ;
        RECT 1923.325 435.010 1923.655 435.025 ;
        RECT 1924.245 435.010 1924.575 435.025 ;
        RECT 1923.325 434.710 1924.575 435.010 ;
        RECT 1923.325 434.695 1923.655 434.710 ;
        RECT 1924.245 434.695 1924.575 434.710 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1931.150 46.480 1931.470 46.540 ;
        RECT 2298.230 46.480 2298.550 46.540 ;
        RECT 1931.150 46.340 2298.550 46.480 ;
        RECT 1931.150 46.280 1931.470 46.340 ;
        RECT 2298.230 46.280 2298.550 46.340 ;
      LAYER via ;
        RECT 1931.180 46.280 1931.440 46.540 ;
        RECT 2298.260 46.280 2298.520 46.540 ;
      LAYER met2 ;
        RECT 1930.270 1220.330 1930.830 1228.680 ;
        RECT 1930.270 1220.190 1931.380 1220.330 ;
        RECT 1930.270 1219.680 1930.830 1220.190 ;
        RECT 1931.240 46.570 1931.380 1220.190 ;
        RECT 1931.180 46.250 1931.440 46.570 ;
        RECT 2298.260 46.250 2298.520 46.570 ;
        RECT 2298.320 2.400 2298.460 46.250 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1939.430 1207.580 1939.750 1207.640 ;
        RECT 1944.950 1207.580 1945.270 1207.640 ;
        RECT 1939.430 1207.440 1945.270 1207.580 ;
        RECT 1939.430 1207.380 1939.750 1207.440 ;
        RECT 1944.950 1207.380 1945.270 1207.440 ;
        RECT 1944.950 46.140 1945.270 46.200 ;
        RECT 2316.170 46.140 2316.490 46.200 ;
        RECT 1944.950 46.000 2316.490 46.140 ;
        RECT 1944.950 45.940 1945.270 46.000 ;
        RECT 2316.170 45.940 2316.490 46.000 ;
      LAYER via ;
        RECT 1939.460 1207.380 1939.720 1207.640 ;
        RECT 1944.980 1207.380 1945.240 1207.640 ;
        RECT 1944.980 45.940 1945.240 46.200 ;
        RECT 2316.200 45.940 2316.460 46.200 ;
      LAYER met2 ;
        RECT 1939.470 1219.680 1940.030 1228.680 ;
        RECT 1939.520 1207.670 1939.660 1219.680 ;
        RECT 1939.460 1207.350 1939.720 1207.670 ;
        RECT 1944.980 1207.350 1945.240 1207.670 ;
        RECT 1945.040 46.230 1945.180 1207.350 ;
        RECT 1944.980 45.910 1945.240 46.230 ;
        RECT 2316.200 45.910 2316.460 46.230 ;
        RECT 2316.260 2.400 2316.400 45.910 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1971.245 1208.785 1971.415 1212.015 ;
      LAYER mcon ;
        RECT 1971.245 1211.845 1971.415 1212.015 ;
      LAYER met1 ;
        RECT 1948.630 1212.000 1948.950 1212.060 ;
        RECT 1971.185 1212.000 1971.475 1212.045 ;
        RECT 1948.630 1211.860 1971.475 1212.000 ;
        RECT 1948.630 1211.800 1948.950 1211.860 ;
        RECT 1971.185 1211.815 1971.475 1211.860 ;
        RECT 1971.185 1208.940 1971.475 1208.985 ;
        RECT 2332.270 1208.940 2332.590 1209.000 ;
        RECT 1971.185 1208.800 2332.590 1208.940 ;
        RECT 1971.185 1208.755 1971.475 1208.800 ;
        RECT 2332.270 1208.740 2332.590 1208.800 ;
      LAYER via ;
        RECT 1948.660 1211.800 1948.920 1212.060 ;
        RECT 2332.300 1208.740 2332.560 1209.000 ;
      LAYER met2 ;
        RECT 1948.670 1219.680 1949.230 1228.680 ;
        RECT 1948.720 1212.090 1948.860 1219.680 ;
        RECT 1948.660 1211.770 1948.920 1212.090 ;
        RECT 2332.300 1208.710 2332.560 1209.030 ;
        RECT 2332.360 16.730 2332.500 1208.710 ;
        RECT 2332.360 16.590 2334.340 16.730 ;
        RECT 2334.200 2.400 2334.340 16.590 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1958.750 45.800 1959.070 45.860 ;
        RECT 2351.590 45.800 2351.910 45.860 ;
        RECT 1958.750 45.660 2351.910 45.800 ;
        RECT 1958.750 45.600 1959.070 45.660 ;
        RECT 2351.590 45.600 2351.910 45.660 ;
      LAYER via ;
        RECT 1958.780 45.600 1959.040 45.860 ;
        RECT 2351.620 45.600 2351.880 45.860 ;
      LAYER met2 ;
        RECT 1957.870 1220.330 1958.430 1228.680 ;
        RECT 1957.870 1220.190 1958.980 1220.330 ;
        RECT 1957.870 1219.680 1958.430 1220.190 ;
        RECT 1958.840 45.890 1958.980 1220.190 ;
        RECT 1958.780 45.570 1959.040 45.890 ;
        RECT 2351.620 45.570 2351.880 45.890 ;
        RECT 2351.680 2.400 2351.820 45.570 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1967.030 1209.620 1967.350 1209.680 ;
        RECT 2366.770 1209.620 2367.090 1209.680 ;
        RECT 1967.030 1209.480 2367.090 1209.620 ;
        RECT 1967.030 1209.420 1967.350 1209.480 ;
        RECT 2366.770 1209.420 2367.090 1209.480 ;
        RECT 2366.770 2.960 2367.090 3.020 ;
        RECT 2369.530 2.960 2369.850 3.020 ;
        RECT 2366.770 2.820 2369.850 2.960 ;
        RECT 2366.770 2.760 2367.090 2.820 ;
        RECT 2369.530 2.760 2369.850 2.820 ;
      LAYER via ;
        RECT 1967.060 1209.420 1967.320 1209.680 ;
        RECT 2366.800 1209.420 2367.060 1209.680 ;
        RECT 2366.800 2.760 2367.060 3.020 ;
        RECT 2369.560 2.760 2369.820 3.020 ;
      LAYER met2 ;
        RECT 1967.070 1219.680 1967.630 1228.680 ;
        RECT 1967.120 1209.710 1967.260 1219.680 ;
        RECT 1967.060 1209.390 1967.320 1209.710 ;
        RECT 2366.800 1209.390 2367.060 1209.710 ;
        RECT 2366.860 3.050 2367.000 1209.390 ;
        RECT 2366.800 2.730 2367.060 3.050 ;
        RECT 2369.560 2.730 2369.820 3.050 ;
        RECT 2369.620 2.400 2369.760 2.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1976.230 1212.000 1976.550 1212.060 ;
        RECT 2100.890 1212.000 2101.210 1212.060 ;
        RECT 1976.230 1211.860 2101.210 1212.000 ;
        RECT 1976.230 1211.800 1976.550 1211.860 ;
        RECT 2100.890 1211.800 2101.210 1211.860 ;
        RECT 2100.890 14.520 2101.210 14.580 ;
        RECT 2387.470 14.520 2387.790 14.580 ;
        RECT 2100.890 14.380 2387.790 14.520 ;
        RECT 2100.890 14.320 2101.210 14.380 ;
        RECT 2387.470 14.320 2387.790 14.380 ;
      LAYER via ;
        RECT 1976.260 1211.800 1976.520 1212.060 ;
        RECT 2100.920 1211.800 2101.180 1212.060 ;
        RECT 2100.920 14.320 2101.180 14.580 ;
        RECT 2387.500 14.320 2387.760 14.580 ;
      LAYER met2 ;
        RECT 1976.270 1219.680 1976.830 1228.680 ;
        RECT 1976.320 1212.090 1976.460 1219.680 ;
        RECT 1976.260 1211.770 1976.520 1212.090 ;
        RECT 2100.920 1211.770 2101.180 1212.090 ;
        RECT 2100.980 14.610 2101.120 1211.770 ;
        RECT 2100.920 14.290 2101.180 14.610 ;
        RECT 2387.500 14.290 2387.760 14.610 ;
        RECT 2387.560 2.400 2387.700 14.290 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2063.705 1212.185 2064.795 1212.355 ;
      LAYER mcon ;
        RECT 2064.625 1212.185 2064.795 1212.355 ;
      LAYER met1 ;
        RECT 1985.430 1212.340 1985.750 1212.400 ;
        RECT 2063.645 1212.340 2063.935 1212.385 ;
        RECT 1985.430 1212.200 2063.935 1212.340 ;
        RECT 1985.430 1212.140 1985.750 1212.200 ;
        RECT 2063.645 1212.155 2063.935 1212.200 ;
        RECT 2064.565 1212.340 2064.855 1212.385 ;
        RECT 2107.790 1212.340 2108.110 1212.400 ;
        RECT 2064.565 1212.200 2108.110 1212.340 ;
        RECT 2064.565 1212.155 2064.855 1212.200 ;
        RECT 2107.790 1212.140 2108.110 1212.200 ;
        RECT 2107.330 14.860 2107.650 14.920 ;
        RECT 2405.410 14.860 2405.730 14.920 ;
        RECT 2107.330 14.720 2405.730 14.860 ;
        RECT 2107.330 14.660 2107.650 14.720 ;
        RECT 2405.410 14.660 2405.730 14.720 ;
      LAYER via ;
        RECT 1985.460 1212.140 1985.720 1212.400 ;
        RECT 2107.820 1212.140 2108.080 1212.400 ;
        RECT 2107.360 14.660 2107.620 14.920 ;
        RECT 2405.440 14.660 2405.700 14.920 ;
      LAYER met2 ;
        RECT 1985.470 1219.680 1986.030 1228.680 ;
        RECT 1985.520 1212.430 1985.660 1219.680 ;
        RECT 1985.460 1212.110 1985.720 1212.430 ;
        RECT 2107.820 1212.110 2108.080 1212.430 ;
        RECT 2107.880 38.490 2108.020 1212.110 ;
        RECT 2107.420 38.350 2108.020 38.490 ;
        RECT 2107.420 14.950 2107.560 38.350 ;
        RECT 2107.360 14.630 2107.620 14.950 ;
        RECT 2405.440 14.630 2405.700 14.950 ;
        RECT 2405.500 2.400 2405.640 14.630 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 799.550 31.520 799.870 31.580 ;
        RECT 1159.730 31.520 1160.050 31.580 ;
        RECT 799.550 31.380 1160.050 31.520 ;
        RECT 799.550 31.320 799.870 31.380 ;
        RECT 1159.730 31.320 1160.050 31.380 ;
      LAYER via ;
        RECT 799.580 31.320 799.840 31.580 ;
        RECT 1159.760 31.320 1160.020 31.580 ;
      LAYER met2 ;
        RECT 1160.230 1220.330 1160.790 1228.680 ;
        RECT 1159.820 1220.190 1160.790 1220.330 ;
        RECT 1159.820 31.610 1159.960 1220.190 ;
        RECT 1160.230 1219.680 1160.790 1220.190 ;
        RECT 799.580 31.290 799.840 31.610 ;
        RECT 1159.760 31.290 1160.020 31.610 ;
        RECT 799.640 2.400 799.780 31.290 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.470 1196.700 1076.790 1196.760 ;
        RECT 1079.230 1196.700 1079.550 1196.760 ;
        RECT 1076.470 1196.560 1079.550 1196.700 ;
        RECT 1076.470 1196.500 1076.790 1196.560 ;
        RECT 1079.230 1196.500 1079.550 1196.560 ;
        RECT 644.990 30.500 645.310 30.560 ;
        RECT 1076.470 30.500 1076.790 30.560 ;
        RECT 644.990 30.360 1076.790 30.500 ;
        RECT 644.990 30.300 645.310 30.360 ;
        RECT 1076.470 30.300 1076.790 30.360 ;
      LAYER via ;
        RECT 1076.500 1196.500 1076.760 1196.760 ;
        RECT 1079.260 1196.500 1079.520 1196.760 ;
        RECT 645.020 30.300 645.280 30.560 ;
        RECT 1076.500 30.300 1076.760 30.560 ;
      LAYER met2 ;
        RECT 1081.110 1220.330 1081.670 1228.680 ;
        RECT 1079.320 1220.190 1081.670 1220.330 ;
        RECT 1079.320 1196.790 1079.460 1220.190 ;
        RECT 1081.110 1219.680 1081.670 1220.190 ;
        RECT 1076.500 1196.470 1076.760 1196.790 ;
        RECT 1079.260 1196.470 1079.520 1196.790 ;
        RECT 1076.560 30.590 1076.700 1196.470 ;
        RECT 645.020 30.270 645.280 30.590 ;
        RECT 1076.500 30.270 1076.760 30.590 ;
        RECT 645.080 2.400 645.220 30.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1997.390 1214.380 1997.710 1214.440 ;
        RECT 2428.870 1214.380 2429.190 1214.440 ;
        RECT 1997.390 1214.240 2429.190 1214.380 ;
        RECT 1997.390 1214.180 1997.710 1214.240 ;
        RECT 2428.870 1214.180 2429.190 1214.240 ;
      LAYER via ;
        RECT 1997.420 1214.180 1997.680 1214.440 ;
        RECT 2428.900 1214.180 2429.160 1214.440 ;
      LAYER met2 ;
        RECT 1997.430 1219.680 1997.990 1228.680 ;
        RECT 1997.480 1214.470 1997.620 1219.680 ;
        RECT 1997.420 1214.150 1997.680 1214.470 ;
        RECT 2428.900 1214.150 2429.160 1214.470 ;
        RECT 2428.960 2.400 2429.100 1214.150 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2114.765 1212.185 2114.935 1213.035 ;
      LAYER mcon ;
        RECT 2114.765 1212.865 2114.935 1213.035 ;
      LAYER met1 ;
        RECT 2006.590 1213.020 2006.910 1213.080 ;
        RECT 2114.705 1213.020 2114.995 1213.065 ;
        RECT 2006.590 1212.880 2114.995 1213.020 ;
        RECT 2006.590 1212.820 2006.910 1212.880 ;
        RECT 2114.705 1212.835 2114.995 1212.880 ;
        RECT 2114.705 1212.340 2114.995 1212.385 ;
        RECT 2156.090 1212.340 2156.410 1212.400 ;
        RECT 2114.705 1212.200 2156.410 1212.340 ;
        RECT 2114.705 1212.155 2114.995 1212.200 ;
        RECT 2156.090 1212.140 2156.410 1212.200 ;
        RECT 2156.090 14.180 2156.410 14.240 ;
        RECT 2446.810 14.180 2447.130 14.240 ;
        RECT 2156.090 14.040 2447.130 14.180 ;
        RECT 2156.090 13.980 2156.410 14.040 ;
        RECT 2446.810 13.980 2447.130 14.040 ;
      LAYER via ;
        RECT 2006.620 1212.820 2006.880 1213.080 ;
        RECT 2156.120 1212.140 2156.380 1212.400 ;
        RECT 2156.120 13.980 2156.380 14.240 ;
        RECT 2446.840 13.980 2447.100 14.240 ;
      LAYER met2 ;
        RECT 2006.630 1219.680 2007.190 1228.680 ;
        RECT 2006.680 1213.110 2006.820 1219.680 ;
        RECT 2006.620 1212.790 2006.880 1213.110 ;
        RECT 2156.120 1212.110 2156.380 1212.430 ;
        RECT 2156.180 14.270 2156.320 1212.110 ;
        RECT 2156.120 13.950 2156.380 14.270 ;
        RECT 2446.840 13.950 2447.100 14.270 ;
        RECT 2446.900 2.400 2447.040 13.950 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2015.790 1213.360 2016.110 1213.420 ;
        RECT 2463.370 1213.360 2463.690 1213.420 ;
        RECT 2015.790 1213.220 2463.690 1213.360 ;
        RECT 2015.790 1213.160 2016.110 1213.220 ;
        RECT 2463.370 1213.160 2463.690 1213.220 ;
      LAYER via ;
        RECT 2015.820 1213.160 2016.080 1213.420 ;
        RECT 2463.400 1213.160 2463.660 1213.420 ;
      LAYER met2 ;
        RECT 2015.830 1219.680 2016.390 1228.680 ;
        RECT 2015.880 1213.450 2016.020 1219.680 ;
        RECT 2015.820 1213.130 2016.080 1213.450 ;
        RECT 2463.400 1213.130 2463.660 1213.450 ;
        RECT 2463.460 3.130 2463.600 1213.130 ;
        RECT 2463.460 2.990 2464.520 3.130 ;
        RECT 2464.380 2.960 2464.520 2.990 ;
        RECT 2464.380 2.820 2464.980 2.960 ;
        RECT 2464.840 2.400 2464.980 2.820 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2024.990 1213.700 2025.310 1213.760 ;
        RECT 2176.790 1213.700 2177.110 1213.760 ;
        RECT 2024.990 1213.560 2177.110 1213.700 ;
        RECT 2024.990 1213.500 2025.310 1213.560 ;
        RECT 2176.790 1213.500 2177.110 1213.560 ;
        RECT 2176.790 15.200 2177.110 15.260 ;
        RECT 2482.690 15.200 2483.010 15.260 ;
        RECT 2176.790 15.060 2483.010 15.200 ;
        RECT 2176.790 15.000 2177.110 15.060 ;
        RECT 2482.690 15.000 2483.010 15.060 ;
      LAYER via ;
        RECT 2025.020 1213.500 2025.280 1213.760 ;
        RECT 2176.820 1213.500 2177.080 1213.760 ;
        RECT 2176.820 15.000 2177.080 15.260 ;
        RECT 2482.720 15.000 2482.980 15.260 ;
      LAYER met2 ;
        RECT 2025.030 1219.680 2025.590 1228.680 ;
        RECT 2025.080 1213.790 2025.220 1219.680 ;
        RECT 2025.020 1213.470 2025.280 1213.790 ;
        RECT 2176.820 1213.470 2177.080 1213.790 ;
        RECT 2176.880 15.290 2177.020 1213.470 ;
        RECT 2176.820 14.970 2177.080 15.290 ;
        RECT 2482.720 14.970 2482.980 15.290 ;
        RECT 2482.780 2.400 2482.920 14.970 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2034.190 1210.980 2034.510 1211.040 ;
        RECT 2497.870 1210.980 2498.190 1211.040 ;
        RECT 2034.190 1210.840 2498.190 1210.980 ;
        RECT 2034.190 1210.780 2034.510 1210.840 ;
        RECT 2497.870 1210.780 2498.190 1210.840 ;
        RECT 2497.870 2.960 2498.190 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2497.870 2.820 2500.950 2.960 ;
        RECT 2497.870 2.760 2498.190 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 2034.220 1210.780 2034.480 1211.040 ;
        RECT 2497.900 1210.780 2498.160 1211.040 ;
        RECT 2497.900 2.760 2498.160 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 2034.230 1219.680 2034.790 1228.680 ;
        RECT 2034.280 1211.070 2034.420 1219.680 ;
        RECT 2034.220 1210.750 2034.480 1211.070 ;
        RECT 2497.900 1210.750 2498.160 1211.070 ;
        RECT 2497.960 3.050 2498.100 1210.750 ;
        RECT 2497.900 2.730 2498.160 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2064.165 1210.485 2064.335 1211.335 ;
        RECT 2091.305 1210.485 2091.475 1211.335 ;
        RECT 2097.745 1207.425 2097.915 1210.655 ;
      LAYER mcon ;
        RECT 2064.165 1211.165 2064.335 1211.335 ;
        RECT 2091.305 1211.165 2091.475 1211.335 ;
        RECT 2097.745 1210.485 2097.915 1210.655 ;
      LAYER met1 ;
        RECT 2064.105 1211.320 2064.395 1211.365 ;
        RECT 2091.245 1211.320 2091.535 1211.365 ;
        RECT 2064.105 1211.180 2091.535 1211.320 ;
        RECT 2064.105 1211.135 2064.395 1211.180 ;
        RECT 2091.245 1211.135 2091.535 1211.180 ;
        RECT 2043.390 1210.640 2043.710 1210.700 ;
        RECT 2064.105 1210.640 2064.395 1210.685 ;
        RECT 2043.390 1210.500 2064.395 1210.640 ;
        RECT 2043.390 1210.440 2043.710 1210.500 ;
        RECT 2064.105 1210.455 2064.395 1210.500 ;
        RECT 2091.245 1210.640 2091.535 1210.685 ;
        RECT 2097.685 1210.640 2097.975 1210.685 ;
        RECT 2091.245 1210.500 2097.975 1210.640 ;
        RECT 2091.245 1210.455 2091.535 1210.500 ;
        RECT 2097.685 1210.455 2097.975 1210.500 ;
        RECT 2097.685 1207.580 2097.975 1207.625 ;
        RECT 2119.290 1207.580 2119.610 1207.640 ;
        RECT 2097.685 1207.440 2104.340 1207.580 ;
        RECT 2097.685 1207.395 2097.975 1207.440 ;
        RECT 2104.200 1207.240 2104.340 1207.440 ;
        RECT 2111.100 1207.440 2119.610 1207.580 ;
        RECT 2111.100 1207.240 2111.240 1207.440 ;
        RECT 2119.290 1207.380 2119.610 1207.440 ;
        RECT 2104.200 1207.100 2111.240 1207.240 ;
        RECT 2121.590 16.560 2121.910 16.620 ;
        RECT 2518.110 16.560 2518.430 16.620 ;
        RECT 2121.590 16.420 2518.430 16.560 ;
        RECT 2121.590 16.360 2121.910 16.420 ;
        RECT 2518.110 16.360 2518.430 16.420 ;
      LAYER via ;
        RECT 2043.420 1210.440 2043.680 1210.700 ;
        RECT 2119.320 1207.380 2119.580 1207.640 ;
        RECT 2121.620 16.360 2121.880 16.620 ;
        RECT 2518.140 16.360 2518.400 16.620 ;
      LAYER met2 ;
        RECT 2043.430 1219.680 2043.990 1228.680 ;
        RECT 2043.480 1210.730 2043.620 1219.680 ;
        RECT 2043.420 1210.410 2043.680 1210.730 ;
        RECT 2119.320 1207.350 2119.580 1207.670 ;
        RECT 2119.380 1193.130 2119.520 1207.350 ;
        RECT 2119.380 1192.990 2121.820 1193.130 ;
        RECT 2121.680 16.650 2121.820 1192.990 ;
        RECT 2121.620 16.330 2121.880 16.650 ;
        RECT 2518.140 16.330 2518.400 16.650 ;
        RECT 2518.200 2.400 2518.340 16.330 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2070.145 1211.505 2070.315 1212.695 ;
      LAYER mcon ;
        RECT 2070.145 1212.525 2070.315 1212.695 ;
      LAYER met1 ;
        RECT 2070.085 1212.680 2070.375 1212.725 ;
        RECT 2514.890 1212.680 2515.210 1212.740 ;
        RECT 2070.085 1212.540 2515.210 1212.680 ;
        RECT 2070.085 1212.495 2070.375 1212.540 ;
        RECT 2514.890 1212.480 2515.210 1212.540 ;
        RECT 2052.590 1211.660 2052.910 1211.720 ;
        RECT 2070.085 1211.660 2070.375 1211.705 ;
        RECT 2052.590 1211.520 2070.375 1211.660 ;
        RECT 2052.590 1211.460 2052.910 1211.520 ;
        RECT 2070.085 1211.475 2070.375 1211.520 ;
        RECT 2514.890 15.200 2515.210 15.260 ;
        RECT 2536.050 15.200 2536.370 15.260 ;
        RECT 2514.890 15.060 2536.370 15.200 ;
        RECT 2514.890 15.000 2515.210 15.060 ;
        RECT 2536.050 15.000 2536.370 15.060 ;
      LAYER via ;
        RECT 2514.920 1212.480 2515.180 1212.740 ;
        RECT 2052.620 1211.460 2052.880 1211.720 ;
        RECT 2514.920 15.000 2515.180 15.260 ;
        RECT 2536.080 15.000 2536.340 15.260 ;
      LAYER met2 ;
        RECT 2052.630 1219.680 2053.190 1228.680 ;
        RECT 2052.680 1211.750 2052.820 1219.680 ;
        RECT 2514.920 1212.450 2515.180 1212.770 ;
        RECT 2052.620 1211.430 2052.880 1211.750 ;
        RECT 2514.980 15.290 2515.120 1212.450 ;
        RECT 2514.920 14.970 2515.180 15.290 ;
        RECT 2536.080 14.970 2536.340 15.290 ;
        RECT 2536.140 2.400 2536.280 14.970 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2091.765 1207.425 2091.935 1211.335 ;
      LAYER mcon ;
        RECT 2091.765 1211.165 2091.935 1211.335 ;
      LAYER met1 ;
        RECT 2091.705 1211.320 2091.995 1211.365 ;
        RECT 2114.690 1211.320 2115.010 1211.380 ;
        RECT 2091.705 1211.180 2115.010 1211.320 ;
        RECT 2091.705 1211.135 2091.995 1211.180 ;
        RECT 2114.690 1211.120 2115.010 1211.180 ;
        RECT 2061.790 1207.580 2062.110 1207.640 ;
        RECT 2091.705 1207.580 2091.995 1207.625 ;
        RECT 2061.790 1207.440 2091.995 1207.580 ;
        RECT 2061.790 1207.380 2062.110 1207.440 ;
        RECT 2091.705 1207.395 2091.995 1207.440 ;
        RECT 2116.070 20.300 2116.390 20.360 ;
        RECT 2553.990 20.300 2554.310 20.360 ;
        RECT 2116.070 20.160 2554.310 20.300 ;
        RECT 2116.070 20.100 2116.390 20.160 ;
        RECT 2553.990 20.100 2554.310 20.160 ;
      LAYER via ;
        RECT 2114.720 1211.120 2114.980 1211.380 ;
        RECT 2061.820 1207.380 2062.080 1207.640 ;
        RECT 2116.100 20.100 2116.360 20.360 ;
        RECT 2554.020 20.100 2554.280 20.360 ;
      LAYER met2 ;
        RECT 2061.830 1219.680 2062.390 1228.680 ;
        RECT 2061.880 1207.670 2062.020 1219.680 ;
        RECT 2114.720 1211.090 2114.980 1211.410 ;
        RECT 2061.820 1207.350 2062.080 1207.670 ;
        RECT 2114.780 41.210 2114.920 1211.090 ;
        RECT 2114.780 41.070 2116.300 41.210 ;
        RECT 2116.160 20.390 2116.300 41.070 ;
        RECT 2116.100 20.070 2116.360 20.390 ;
        RECT 2554.020 20.070 2554.280 20.390 ;
        RECT 2554.080 2.400 2554.220 20.070 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2090.845 1211.505 2091.015 1214.735 ;
      LAYER mcon ;
        RECT 2090.845 1214.565 2091.015 1214.735 ;
      LAYER met1 ;
        RECT 2072.370 1214.720 2072.690 1214.780 ;
        RECT 2090.785 1214.720 2091.075 1214.765 ;
        RECT 2072.370 1214.580 2091.075 1214.720 ;
        RECT 2072.370 1214.520 2072.690 1214.580 ;
        RECT 2090.785 1214.535 2091.075 1214.580 ;
        RECT 2090.785 1211.660 2091.075 1211.705 ;
        RECT 2535.590 1211.660 2535.910 1211.720 ;
        RECT 2090.785 1211.520 2535.910 1211.660 ;
        RECT 2090.785 1211.475 2091.075 1211.520 ;
        RECT 2535.590 1211.460 2535.910 1211.520 ;
        RECT 2535.590 20.640 2535.910 20.700 ;
        RECT 2571.930 20.640 2572.250 20.700 ;
        RECT 2535.590 20.500 2572.250 20.640 ;
        RECT 2535.590 20.440 2535.910 20.500 ;
        RECT 2571.930 20.440 2572.250 20.500 ;
      LAYER via ;
        RECT 2072.400 1214.520 2072.660 1214.780 ;
        RECT 2535.620 1211.460 2535.880 1211.720 ;
        RECT 2535.620 20.440 2535.880 20.700 ;
        RECT 2571.960 20.440 2572.220 20.700 ;
      LAYER met2 ;
        RECT 2071.030 1220.330 2071.590 1228.680 ;
        RECT 2071.030 1220.190 2072.600 1220.330 ;
        RECT 2071.030 1219.680 2071.590 1220.190 ;
        RECT 2072.460 1214.810 2072.600 1220.190 ;
        RECT 2072.400 1214.490 2072.660 1214.810 ;
        RECT 2535.620 1211.430 2535.880 1211.750 ;
        RECT 2535.680 20.730 2535.820 1211.430 ;
        RECT 2535.620 20.410 2535.880 20.730 ;
        RECT 2571.960 20.410 2572.220 20.730 ;
        RECT 2572.020 2.400 2572.160 20.410 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2080.190 1211.660 2080.510 1211.720 ;
        RECT 2083.410 1211.660 2083.730 1211.720 ;
        RECT 2080.190 1211.520 2083.730 1211.660 ;
        RECT 2080.190 1211.460 2080.510 1211.520 ;
        RECT 2083.410 1211.460 2083.730 1211.520 ;
        RECT 2083.410 19.960 2083.730 20.020 ;
        RECT 2589.410 19.960 2589.730 20.020 ;
        RECT 2083.410 19.820 2589.730 19.960 ;
        RECT 2083.410 19.760 2083.730 19.820 ;
        RECT 2589.410 19.760 2589.730 19.820 ;
      LAYER via ;
        RECT 2080.220 1211.460 2080.480 1211.720 ;
        RECT 2083.440 1211.460 2083.700 1211.720 ;
        RECT 2083.440 19.760 2083.700 20.020 ;
        RECT 2589.440 19.760 2589.700 20.020 ;
      LAYER met2 ;
        RECT 2080.230 1219.680 2080.790 1228.680 ;
        RECT 2080.280 1211.750 2080.420 1219.680 ;
        RECT 2080.220 1211.430 2080.480 1211.750 ;
        RECT 2083.440 1211.430 2083.700 1211.750 ;
        RECT 2083.500 20.050 2083.640 1211.430 ;
        RECT 2083.440 19.730 2083.700 20.050 ;
        RECT 2589.440 19.730 2589.700 20.050 ;
        RECT 2589.500 2.400 2589.640 19.730 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.630 1196.700 1166.950 1196.760 ;
        RECT 1171.230 1196.700 1171.550 1196.760 ;
        RECT 1166.630 1196.560 1171.550 1196.700 ;
        RECT 1166.630 1196.500 1166.950 1196.560 ;
        RECT 1171.230 1196.500 1171.550 1196.560 ;
        RECT 823.470 28.120 823.790 28.180 ;
        RECT 1166.630 28.120 1166.950 28.180 ;
        RECT 823.470 27.980 1166.950 28.120 ;
        RECT 823.470 27.920 823.790 27.980 ;
        RECT 1166.630 27.920 1166.950 27.980 ;
      LAYER via ;
        RECT 1166.660 1196.500 1166.920 1196.760 ;
        RECT 1171.260 1196.500 1171.520 1196.760 ;
        RECT 823.500 27.920 823.760 28.180 ;
        RECT 1166.660 27.920 1166.920 28.180 ;
      LAYER met2 ;
        RECT 1172.650 1220.330 1173.210 1228.680 ;
        RECT 1171.320 1220.190 1173.210 1220.330 ;
        RECT 1171.320 1196.790 1171.460 1220.190 ;
        RECT 1172.650 1219.680 1173.210 1220.190 ;
        RECT 1166.660 1196.470 1166.920 1196.790 ;
        RECT 1171.260 1196.470 1171.520 1196.790 ;
        RECT 1166.720 28.210 1166.860 1196.470 ;
        RECT 823.500 27.890 823.760 28.210 ;
        RECT 1166.660 27.890 1166.920 28.210 ;
        RECT 823.560 2.400 823.700 27.890 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2556.290 20.300 2556.610 20.360 ;
        RECT 2607.350 20.300 2607.670 20.360 ;
        RECT 2556.290 20.160 2607.670 20.300 ;
        RECT 2556.290 20.100 2556.610 20.160 ;
        RECT 2607.350 20.100 2607.670 20.160 ;
      LAYER via ;
        RECT 2556.320 20.100 2556.580 20.360 ;
        RECT 2607.380 20.100 2607.640 20.360 ;
      LAYER met2 ;
        RECT 2088.970 1219.680 2089.530 1228.680 ;
        RECT 2089.020 1210.925 2089.160 1219.680 ;
        RECT 2088.950 1210.555 2089.230 1210.925 ;
        RECT 2556.310 1210.555 2556.590 1210.925 ;
        RECT 2556.380 20.390 2556.520 1210.555 ;
        RECT 2556.320 20.070 2556.580 20.390 ;
        RECT 2607.380 20.070 2607.640 20.390 ;
        RECT 2607.440 2.400 2607.580 20.070 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
      LAYER via2 ;
        RECT 2088.950 1210.600 2089.230 1210.880 ;
        RECT 2556.310 1210.600 2556.590 1210.880 ;
      LAYER met3 ;
        RECT 2088.925 1210.890 2089.255 1210.905 ;
        RECT 2556.285 1210.890 2556.615 1210.905 ;
        RECT 2088.925 1210.590 2556.615 1210.890 ;
        RECT 2088.925 1210.575 2089.255 1210.590 ;
        RECT 2556.285 1210.575 2556.615 1210.590 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2098.130 1210.640 2098.450 1210.700 ;
        RECT 2108.250 1210.640 2108.570 1210.700 ;
        RECT 2098.130 1210.500 2108.570 1210.640 ;
        RECT 2098.130 1210.440 2098.450 1210.500 ;
        RECT 2108.250 1210.440 2108.570 1210.500 ;
        RECT 2108.250 19.620 2108.570 19.680 ;
        RECT 2625.290 19.620 2625.610 19.680 ;
        RECT 2108.250 19.480 2625.610 19.620 ;
        RECT 2108.250 19.420 2108.570 19.480 ;
        RECT 2625.290 19.420 2625.610 19.480 ;
      LAYER via ;
        RECT 2098.160 1210.440 2098.420 1210.700 ;
        RECT 2108.280 1210.440 2108.540 1210.700 ;
        RECT 2108.280 19.420 2108.540 19.680 ;
        RECT 2625.320 19.420 2625.580 19.680 ;
      LAYER met2 ;
        RECT 2098.170 1219.680 2098.730 1228.680 ;
        RECT 2098.220 1210.730 2098.360 1219.680 ;
        RECT 2098.160 1210.410 2098.420 1210.730 ;
        RECT 2108.280 1210.410 2108.540 1210.730 ;
        RECT 2108.340 19.710 2108.480 1210.410 ;
        RECT 2108.280 19.390 2108.540 19.710 ;
        RECT 2625.320 19.390 2625.580 19.710 ;
        RECT 2625.380 2.400 2625.520 19.390 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2107.330 1212.000 2107.650 1212.060 ;
        RECT 2570.090 1212.000 2570.410 1212.060 ;
        RECT 2107.330 1211.860 2570.410 1212.000 ;
        RECT 2107.330 1211.800 2107.650 1211.860 ;
        RECT 2570.090 1211.800 2570.410 1211.860 ;
        RECT 2570.090 15.880 2570.410 15.940 ;
        RECT 2643.230 15.880 2643.550 15.940 ;
        RECT 2570.090 15.740 2643.550 15.880 ;
        RECT 2570.090 15.680 2570.410 15.740 ;
        RECT 2643.230 15.680 2643.550 15.740 ;
      LAYER via ;
        RECT 2107.360 1211.800 2107.620 1212.060 ;
        RECT 2570.120 1211.800 2570.380 1212.060 ;
        RECT 2570.120 15.680 2570.380 15.940 ;
        RECT 2643.260 15.680 2643.520 15.940 ;
      LAYER met2 ;
        RECT 2107.370 1219.680 2107.930 1228.680 ;
        RECT 2107.420 1212.090 2107.560 1219.680 ;
        RECT 2107.360 1211.770 2107.620 1212.090 ;
        RECT 2570.120 1211.770 2570.380 1212.090 ;
        RECT 2570.180 15.970 2570.320 1211.770 ;
        RECT 2570.120 15.650 2570.380 15.970 ;
        RECT 2643.260 15.650 2643.520 15.970 ;
        RECT 2643.320 2.400 2643.460 15.650 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 19.280 2118.230 19.340 ;
        RECT 2661.170 19.280 2661.490 19.340 ;
        RECT 2117.910 19.140 2661.490 19.280 ;
        RECT 2117.910 19.080 2118.230 19.140 ;
        RECT 2661.170 19.080 2661.490 19.140 ;
      LAYER via ;
        RECT 2117.940 19.080 2118.200 19.340 ;
        RECT 2661.200 19.080 2661.460 19.340 ;
      LAYER met2 ;
        RECT 2116.570 1220.330 2117.130 1228.680 ;
        RECT 2116.570 1220.190 2118.140 1220.330 ;
        RECT 2116.570 1219.680 2117.130 1220.190 ;
        RECT 2118.000 19.370 2118.140 1220.190 ;
        RECT 2117.940 19.050 2118.200 19.370 ;
        RECT 2661.200 19.050 2661.460 19.370 ;
        RECT 2661.260 2.400 2661.400 19.050 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2159.385 1212.865 2160.015 1213.035 ;
        RECT 2159.845 1212.185 2160.015 1212.865 ;
      LAYER met1 ;
        RECT 2125.730 1213.020 2126.050 1213.080 ;
        RECT 2159.325 1213.020 2159.615 1213.065 ;
        RECT 2125.730 1212.880 2159.615 1213.020 ;
        RECT 2125.730 1212.820 2126.050 1212.880 ;
        RECT 2159.325 1212.835 2159.615 1212.880 ;
        RECT 2159.785 1212.340 2160.075 1212.385 ;
        RECT 2590.790 1212.340 2591.110 1212.400 ;
        RECT 2159.785 1212.200 2591.110 1212.340 ;
        RECT 2159.785 1212.155 2160.075 1212.200 ;
        RECT 2590.790 1212.140 2591.110 1212.200 ;
        RECT 2590.790 16.220 2591.110 16.280 ;
        RECT 2678.650 16.220 2678.970 16.280 ;
        RECT 2590.790 16.080 2678.970 16.220 ;
        RECT 2590.790 16.020 2591.110 16.080 ;
        RECT 2678.650 16.020 2678.970 16.080 ;
      LAYER via ;
        RECT 2125.760 1212.820 2126.020 1213.080 ;
        RECT 2590.820 1212.140 2591.080 1212.400 ;
        RECT 2590.820 16.020 2591.080 16.280 ;
        RECT 2678.680 16.020 2678.940 16.280 ;
      LAYER met2 ;
        RECT 2125.770 1219.680 2126.330 1228.680 ;
        RECT 2125.820 1213.110 2125.960 1219.680 ;
        RECT 2125.760 1212.790 2126.020 1213.110 ;
        RECT 2590.820 1212.110 2591.080 1212.430 ;
        RECT 2590.880 16.310 2591.020 1212.110 ;
        RECT 2590.820 15.990 2591.080 16.310 ;
        RECT 2678.680 15.990 2678.940 16.310 ;
        RECT 2678.740 2.400 2678.880 15.990 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2134.930 1207.580 2135.250 1207.640 ;
        RECT 2138.610 1207.580 2138.930 1207.640 ;
        RECT 2134.930 1207.440 2138.930 1207.580 ;
        RECT 2134.930 1207.380 2135.250 1207.440 ;
        RECT 2138.610 1207.380 2138.930 1207.440 ;
        RECT 2138.610 18.940 2138.930 19.000 ;
        RECT 2696.590 18.940 2696.910 19.000 ;
        RECT 2138.610 18.800 2696.910 18.940 ;
        RECT 2138.610 18.740 2138.930 18.800 ;
        RECT 2696.590 18.740 2696.910 18.800 ;
      LAYER via ;
        RECT 2134.960 1207.380 2135.220 1207.640 ;
        RECT 2138.640 1207.380 2138.900 1207.640 ;
        RECT 2138.640 18.740 2138.900 19.000 ;
        RECT 2696.620 18.740 2696.880 19.000 ;
      LAYER met2 ;
        RECT 2134.970 1219.680 2135.530 1228.680 ;
        RECT 2135.020 1207.670 2135.160 1219.680 ;
        RECT 2134.960 1207.350 2135.220 1207.670 ;
        RECT 2138.640 1207.350 2138.900 1207.670 ;
        RECT 2138.700 19.030 2138.840 1207.350 ;
        RECT 2138.640 18.710 2138.900 19.030 ;
        RECT 2696.620 18.710 2696.880 19.030 ;
        RECT 2696.680 2.400 2696.820 18.710 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2144.130 1211.320 2144.450 1211.380 ;
        RECT 2604.590 1211.320 2604.910 1211.380 ;
        RECT 2144.130 1211.180 2604.910 1211.320 ;
        RECT 2144.130 1211.120 2144.450 1211.180 ;
        RECT 2604.590 1211.120 2604.910 1211.180 ;
        RECT 2604.590 16.560 2604.910 16.620 ;
        RECT 2714.530 16.560 2714.850 16.620 ;
        RECT 2604.590 16.420 2714.850 16.560 ;
        RECT 2604.590 16.360 2604.910 16.420 ;
        RECT 2714.530 16.360 2714.850 16.420 ;
      LAYER via ;
        RECT 2144.160 1211.120 2144.420 1211.380 ;
        RECT 2604.620 1211.120 2604.880 1211.380 ;
        RECT 2604.620 16.360 2604.880 16.620 ;
        RECT 2714.560 16.360 2714.820 16.620 ;
      LAYER met2 ;
        RECT 2144.170 1219.680 2144.730 1228.680 ;
        RECT 2144.220 1211.410 2144.360 1219.680 ;
        RECT 2144.160 1211.090 2144.420 1211.410 ;
        RECT 2604.620 1211.090 2604.880 1211.410 ;
        RECT 2604.680 16.650 2604.820 1211.090 ;
        RECT 2604.620 16.330 2604.880 16.650 ;
        RECT 2714.560 16.330 2714.820 16.650 ;
        RECT 2714.620 2.400 2714.760 16.330 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2153.330 1207.580 2153.650 1207.640 ;
        RECT 2153.330 1207.440 2158.160 1207.580 ;
        RECT 2153.330 1207.380 2153.650 1207.440 ;
        RECT 2158.020 1206.900 2158.160 1207.440 ;
        RECT 2159.310 1206.900 2159.630 1206.960 ;
        RECT 2158.020 1206.760 2159.630 1206.900 ;
        RECT 2159.310 1206.700 2159.630 1206.760 ;
        RECT 2159.310 18.600 2159.630 18.660 ;
        RECT 2732.470 18.600 2732.790 18.660 ;
        RECT 2159.310 18.460 2732.790 18.600 ;
        RECT 2159.310 18.400 2159.630 18.460 ;
        RECT 2732.470 18.400 2732.790 18.460 ;
      LAYER via ;
        RECT 2153.360 1207.380 2153.620 1207.640 ;
        RECT 2159.340 1206.700 2159.600 1206.960 ;
        RECT 2159.340 18.400 2159.600 18.660 ;
        RECT 2732.500 18.400 2732.760 18.660 ;
      LAYER met2 ;
        RECT 2153.370 1219.680 2153.930 1228.680 ;
        RECT 2153.420 1207.670 2153.560 1219.680 ;
        RECT 2153.360 1207.350 2153.620 1207.670 ;
        RECT 2159.340 1206.670 2159.600 1206.990 ;
        RECT 2159.400 18.690 2159.540 1206.670 ;
        RECT 2159.340 18.370 2159.600 18.690 ;
        RECT 2732.500 18.370 2732.760 18.690 ;
        RECT 2732.560 2.400 2732.700 18.370 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2162.530 1213.020 2162.850 1213.080 ;
        RECT 2618.390 1213.020 2618.710 1213.080 ;
        RECT 2162.530 1212.880 2618.710 1213.020 ;
        RECT 2162.530 1212.820 2162.850 1212.880 ;
        RECT 2618.390 1212.820 2618.710 1212.880 ;
        RECT 2618.390 16.900 2618.710 16.960 ;
        RECT 2750.410 16.900 2750.730 16.960 ;
        RECT 2618.390 16.760 2750.730 16.900 ;
        RECT 2618.390 16.700 2618.710 16.760 ;
        RECT 2750.410 16.700 2750.730 16.760 ;
      LAYER via ;
        RECT 2162.560 1212.820 2162.820 1213.080 ;
        RECT 2618.420 1212.820 2618.680 1213.080 ;
        RECT 2618.420 16.700 2618.680 16.960 ;
        RECT 2750.440 16.700 2750.700 16.960 ;
      LAYER met2 ;
        RECT 2162.570 1219.680 2163.130 1228.680 ;
        RECT 2162.620 1213.110 2162.760 1219.680 ;
        RECT 2162.560 1212.790 2162.820 1213.110 ;
        RECT 2618.420 1212.790 2618.680 1213.110 ;
        RECT 2618.480 16.990 2618.620 1212.790 ;
        RECT 2618.420 16.670 2618.680 16.990 ;
        RECT 2750.440 16.670 2750.700 16.990 ;
        RECT 2750.500 2.400 2750.640 16.670 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.110 18.260 2173.430 18.320 ;
        RECT 2767.890 18.260 2768.210 18.320 ;
        RECT 2173.110 18.120 2768.210 18.260 ;
        RECT 2173.110 18.060 2173.430 18.120 ;
        RECT 2767.890 18.060 2768.210 18.120 ;
      LAYER via ;
        RECT 2173.140 18.060 2173.400 18.320 ;
        RECT 2767.920 18.060 2768.180 18.320 ;
      LAYER met2 ;
        RECT 2171.770 1220.330 2172.330 1228.680 ;
        RECT 2171.770 1220.190 2173.340 1220.330 ;
        RECT 2171.770 1219.680 2172.330 1220.190 ;
        RECT 2173.200 18.350 2173.340 1220.190 ;
        RECT 2173.140 18.030 2173.400 18.350 ;
        RECT 2767.920 18.030 2768.180 18.350 ;
        RECT 2767.980 2.400 2768.120 18.030 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 27.780 841.270 27.840 ;
        RECT 1180.430 27.780 1180.750 27.840 ;
        RECT 840.950 27.640 1180.750 27.780 ;
        RECT 840.950 27.580 841.270 27.640 ;
        RECT 1180.430 27.580 1180.750 27.640 ;
      LAYER via ;
        RECT 840.980 27.580 841.240 27.840 ;
        RECT 1180.460 27.580 1180.720 27.840 ;
      LAYER met2 ;
        RECT 1181.850 1220.330 1182.410 1228.680 ;
        RECT 1180.520 1220.190 1182.410 1220.330 ;
        RECT 1180.520 27.870 1180.660 1220.190 ;
        RECT 1181.850 1219.680 1182.410 1220.190 ;
        RECT 840.980 27.550 841.240 27.870 ;
        RECT 1180.460 27.550 1180.720 27.870 ;
        RECT 841.040 2.400 841.180 27.550 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.930 1213.700 2181.250 1213.760 ;
        RECT 2625.290 1213.700 2625.610 1213.760 ;
        RECT 2180.930 1213.560 2625.610 1213.700 ;
        RECT 2180.930 1213.500 2181.250 1213.560 ;
        RECT 2625.290 1213.500 2625.610 1213.560 ;
        RECT 2625.290 20.640 2625.610 20.700 ;
        RECT 2785.830 20.640 2786.150 20.700 ;
        RECT 2625.290 20.500 2786.150 20.640 ;
        RECT 2625.290 20.440 2625.610 20.500 ;
        RECT 2785.830 20.440 2786.150 20.500 ;
      LAYER via ;
        RECT 2180.960 1213.500 2181.220 1213.760 ;
        RECT 2625.320 1213.500 2625.580 1213.760 ;
        RECT 2625.320 20.440 2625.580 20.700 ;
        RECT 2785.860 20.440 2786.120 20.700 ;
      LAYER met2 ;
        RECT 2180.970 1219.680 2181.530 1228.680 ;
        RECT 2181.020 1213.790 2181.160 1219.680 ;
        RECT 2180.960 1213.470 2181.220 1213.790 ;
        RECT 2625.320 1213.470 2625.580 1213.790 ;
        RECT 2625.380 20.730 2625.520 1213.470 ;
        RECT 2625.320 20.410 2625.580 20.730 ;
        RECT 2785.860 20.410 2786.120 20.730 ;
        RECT 2785.920 2.400 2786.060 20.410 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2190.130 1207.580 2190.450 1207.640 ;
        RECT 2193.810 1207.580 2194.130 1207.640 ;
        RECT 2190.130 1207.440 2194.130 1207.580 ;
        RECT 2190.130 1207.380 2190.450 1207.440 ;
        RECT 2193.810 1207.380 2194.130 1207.440 ;
        RECT 2193.810 17.920 2194.130 17.980 ;
        RECT 2803.770 17.920 2804.090 17.980 ;
        RECT 2193.810 17.780 2804.090 17.920 ;
        RECT 2193.810 17.720 2194.130 17.780 ;
        RECT 2803.770 17.720 2804.090 17.780 ;
      LAYER via ;
        RECT 2190.160 1207.380 2190.420 1207.640 ;
        RECT 2193.840 1207.380 2194.100 1207.640 ;
        RECT 2193.840 17.720 2194.100 17.980 ;
        RECT 2803.800 17.720 2804.060 17.980 ;
      LAYER met2 ;
        RECT 2190.170 1219.680 2190.730 1228.680 ;
        RECT 2190.220 1207.670 2190.360 1219.680 ;
        RECT 2190.160 1207.350 2190.420 1207.670 ;
        RECT 2193.840 1207.350 2194.100 1207.670 ;
        RECT 2193.900 18.010 2194.040 1207.350 ;
        RECT 2193.840 17.690 2194.100 18.010 ;
        RECT 2803.800 17.690 2804.060 18.010 ;
        RECT 2803.860 2.400 2804.000 17.690 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2201.170 1207.580 2201.490 1207.640 ;
        RECT 2639.090 1207.580 2639.410 1207.640 ;
        RECT 2201.170 1207.440 2639.410 1207.580 ;
        RECT 2201.170 1207.380 2201.490 1207.440 ;
        RECT 2639.090 1207.380 2639.410 1207.440 ;
        RECT 2639.090 20.300 2639.410 20.360 ;
        RECT 2821.710 20.300 2822.030 20.360 ;
        RECT 2639.090 20.160 2822.030 20.300 ;
        RECT 2639.090 20.100 2639.410 20.160 ;
        RECT 2821.710 20.100 2822.030 20.160 ;
      LAYER via ;
        RECT 2201.200 1207.380 2201.460 1207.640 ;
        RECT 2639.120 1207.380 2639.380 1207.640 ;
        RECT 2639.120 20.100 2639.380 20.360 ;
        RECT 2821.740 20.100 2822.000 20.360 ;
      LAYER met2 ;
        RECT 2199.370 1220.330 2199.930 1228.680 ;
        RECT 2199.370 1220.190 2200.940 1220.330 ;
        RECT 2199.370 1219.680 2199.930 1220.190 ;
        RECT 2200.800 1208.090 2200.940 1220.190 ;
        RECT 2200.800 1207.950 2201.400 1208.090 ;
        RECT 2201.260 1207.670 2201.400 1207.950 ;
        RECT 2201.200 1207.350 2201.460 1207.670 ;
        RECT 2639.120 1207.350 2639.380 1207.670 ;
        RECT 2639.180 20.390 2639.320 1207.350 ;
        RECT 2639.120 20.070 2639.380 20.390 ;
        RECT 2821.740 20.070 2822.000 20.390 ;
        RECT 2821.800 2.400 2821.940 20.070 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2208.530 1210.640 2208.850 1210.700 ;
        RECT 2214.970 1210.640 2215.290 1210.700 ;
        RECT 2208.530 1210.500 2215.290 1210.640 ;
        RECT 2208.530 1210.440 2208.850 1210.500 ;
        RECT 2214.970 1210.440 2215.290 1210.500 ;
        RECT 2214.510 17.580 2214.830 17.640 ;
        RECT 2839.190 17.580 2839.510 17.640 ;
        RECT 2214.510 17.440 2839.510 17.580 ;
        RECT 2214.510 17.380 2214.830 17.440 ;
        RECT 2839.190 17.380 2839.510 17.440 ;
      LAYER via ;
        RECT 2208.560 1210.440 2208.820 1210.700 ;
        RECT 2215.000 1210.440 2215.260 1210.700 ;
        RECT 2214.540 17.380 2214.800 17.640 ;
        RECT 2839.220 17.380 2839.480 17.640 ;
      LAYER met2 ;
        RECT 2208.570 1219.680 2209.130 1228.680 ;
        RECT 2208.620 1210.730 2208.760 1219.680 ;
        RECT 2208.560 1210.410 2208.820 1210.730 ;
        RECT 2215.000 1210.410 2215.260 1210.730 ;
        RECT 2215.060 1209.450 2215.200 1210.410 ;
        RECT 2214.600 1209.310 2215.200 1209.450 ;
        RECT 2214.600 17.670 2214.740 1209.310 ;
        RECT 2214.540 17.350 2214.800 17.670 ;
        RECT 2839.220 17.350 2839.480 17.670 ;
        RECT 2839.280 2.400 2839.420 17.350 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2250.005 1210.485 2250.175 1214.055 ;
      LAYER mcon ;
        RECT 2250.005 1213.885 2250.175 1214.055 ;
      LAYER met1 ;
        RECT 2217.270 1214.040 2217.590 1214.100 ;
        RECT 2249.945 1214.040 2250.235 1214.085 ;
        RECT 2217.270 1213.900 2250.235 1214.040 ;
        RECT 2217.270 1213.840 2217.590 1213.900 ;
        RECT 2249.945 1213.855 2250.235 1213.900 ;
        RECT 2249.945 1210.640 2250.235 1210.685 ;
        RECT 2645.990 1210.640 2646.310 1210.700 ;
        RECT 2249.945 1210.500 2646.310 1210.640 ;
        RECT 2249.945 1210.455 2250.235 1210.500 ;
        RECT 2645.990 1210.440 2646.310 1210.500 ;
        RECT 2645.990 19.960 2646.310 20.020 ;
        RECT 2857.130 19.960 2857.450 20.020 ;
        RECT 2645.990 19.820 2857.450 19.960 ;
        RECT 2645.990 19.760 2646.310 19.820 ;
        RECT 2857.130 19.760 2857.450 19.820 ;
      LAYER via ;
        RECT 2217.300 1213.840 2217.560 1214.100 ;
        RECT 2646.020 1210.440 2646.280 1210.700 ;
        RECT 2646.020 19.760 2646.280 20.020 ;
        RECT 2857.160 19.760 2857.420 20.020 ;
      LAYER met2 ;
        RECT 2217.310 1219.680 2217.870 1228.680 ;
        RECT 2217.360 1214.130 2217.500 1219.680 ;
        RECT 2217.300 1213.810 2217.560 1214.130 ;
        RECT 2646.020 1210.410 2646.280 1210.730 ;
        RECT 2646.080 20.050 2646.220 1210.410 ;
        RECT 2646.020 19.730 2646.280 20.050 ;
        RECT 2857.160 19.730 2857.420 20.050 ;
        RECT 2857.220 2.400 2857.360 19.730 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2228.310 17.240 2228.630 17.300 ;
        RECT 2875.070 17.240 2875.390 17.300 ;
        RECT 2228.310 17.100 2875.390 17.240 ;
        RECT 2228.310 17.040 2228.630 17.100 ;
        RECT 2875.070 17.040 2875.390 17.100 ;
      LAYER via ;
        RECT 2228.340 17.040 2228.600 17.300 ;
        RECT 2875.100 17.040 2875.360 17.300 ;
      LAYER met2 ;
        RECT 2226.510 1220.330 2227.070 1228.680 ;
        RECT 2226.510 1220.190 2228.540 1220.330 ;
        RECT 2226.510 1219.680 2227.070 1220.190 ;
        RECT 2228.400 17.330 2228.540 1220.190 ;
        RECT 2228.340 17.010 2228.600 17.330 ;
        RECT 2875.100 17.010 2875.360 17.330 ;
        RECT 2875.160 2.400 2875.300 17.010 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2235.670 1210.640 2235.990 1210.700 ;
        RECT 2235.670 1210.500 2249.700 1210.640 ;
        RECT 2235.670 1210.440 2235.990 1210.500 ;
        RECT 2249.560 1210.300 2249.700 1210.500 ;
        RECT 2652.890 1210.300 2653.210 1210.360 ;
        RECT 2249.560 1210.160 2653.210 1210.300 ;
        RECT 2652.890 1210.100 2653.210 1210.160 ;
        RECT 2652.890 19.620 2653.210 19.680 ;
        RECT 2893.010 19.620 2893.330 19.680 ;
        RECT 2652.890 19.480 2893.330 19.620 ;
        RECT 2652.890 19.420 2653.210 19.480 ;
        RECT 2893.010 19.420 2893.330 19.480 ;
      LAYER via ;
        RECT 2235.700 1210.440 2235.960 1210.700 ;
        RECT 2652.920 1210.100 2653.180 1210.360 ;
        RECT 2652.920 19.420 2653.180 19.680 ;
        RECT 2893.040 19.420 2893.300 19.680 ;
      LAYER met2 ;
        RECT 2235.710 1219.680 2236.270 1228.680 ;
        RECT 2235.760 1210.730 2235.900 1219.680 ;
        RECT 2235.700 1210.410 2235.960 1210.730 ;
        RECT 2652.920 1210.070 2653.180 1210.390 ;
        RECT 2652.980 19.710 2653.120 1210.070 ;
        RECT 2652.920 19.390 2653.180 19.710 ;
        RECT 2893.040 19.390 2893.300 19.710 ;
        RECT 2893.100 2.400 2893.240 19.390 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2244.870 1210.300 2245.190 1210.360 ;
        RECT 2249.010 1210.300 2249.330 1210.360 ;
        RECT 2244.870 1210.160 2249.330 1210.300 ;
        RECT 2244.870 1210.100 2245.190 1210.160 ;
        RECT 2249.010 1210.100 2249.330 1210.160 ;
      LAYER via ;
        RECT 2244.900 1210.100 2245.160 1210.360 ;
        RECT 2249.040 1210.100 2249.300 1210.360 ;
      LAYER met2 ;
        RECT 2244.910 1219.680 2245.470 1228.680 ;
        RECT 2244.960 1210.390 2245.100 1219.680 ;
        RECT 2244.900 1210.070 2245.160 1210.390 ;
        RECT 2249.040 1210.070 2249.300 1210.390 ;
        RECT 2249.100 16.845 2249.240 1210.070 ;
        RECT 2249.030 16.475 2249.310 16.845 ;
        RECT 2910.970 16.475 2911.250 16.845 ;
        RECT 2911.040 2.400 2911.180 16.475 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 2249.030 16.520 2249.310 16.800 ;
        RECT 2910.970 16.520 2911.250 16.800 ;
      LAYER met3 ;
        RECT 2249.005 16.810 2249.335 16.825 ;
        RECT 2910.945 16.810 2911.275 16.825 ;
        RECT 2249.005 16.510 2911.275 16.810 ;
        RECT 2249.005 16.495 2249.335 16.510 ;
        RECT 2910.945 16.495 2911.275 16.510 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1188.325 1159.145 1188.495 1197.055 ;
        RECT 1187.865 786.165 1188.035 821.015 ;
      LAYER mcon ;
        RECT 1188.325 1196.885 1188.495 1197.055 ;
        RECT 1187.865 820.845 1188.035 821.015 ;
      LAYER met1 ;
        RECT 1188.265 1197.040 1188.555 1197.085 ;
        RECT 1188.710 1197.040 1189.030 1197.100 ;
        RECT 1188.265 1196.900 1189.030 1197.040 ;
        RECT 1188.265 1196.855 1188.555 1196.900 ;
        RECT 1188.710 1196.840 1189.030 1196.900 ;
        RECT 1188.250 1159.300 1188.570 1159.360 ;
        RECT 1188.055 1159.160 1188.570 1159.300 ;
        RECT 1188.250 1159.100 1188.570 1159.160 ;
        RECT 1187.790 966.180 1188.110 966.240 ;
        RECT 1188.710 966.180 1189.030 966.240 ;
        RECT 1187.790 966.040 1189.030 966.180 ;
        RECT 1187.790 965.980 1188.110 966.040 ;
        RECT 1188.710 965.980 1189.030 966.040 ;
        RECT 1187.790 869.620 1188.110 869.680 ;
        RECT 1188.710 869.620 1189.030 869.680 ;
        RECT 1187.790 869.480 1189.030 869.620 ;
        RECT 1187.790 869.420 1188.110 869.480 ;
        RECT 1188.710 869.420 1189.030 869.480 ;
        RECT 1187.790 821.000 1188.110 821.060 ;
        RECT 1187.595 820.860 1188.110 821.000 ;
        RECT 1187.790 820.800 1188.110 820.860 ;
        RECT 1187.790 786.320 1188.110 786.380 ;
        RECT 1187.595 786.180 1188.110 786.320 ;
        RECT 1187.790 786.120 1188.110 786.180 ;
        RECT 1187.790 724.440 1188.110 724.500 ;
        RECT 1188.250 724.440 1188.570 724.500 ;
        RECT 1187.790 724.300 1188.570 724.440 ;
        RECT 1187.790 724.240 1188.110 724.300 ;
        RECT 1188.250 724.240 1188.570 724.300 ;
        RECT 1187.790 579.400 1188.110 579.660 ;
        RECT 1187.880 579.260 1188.020 579.400 ;
        RECT 1188.250 579.260 1188.570 579.320 ;
        RECT 1187.880 579.120 1188.570 579.260 ;
        RECT 1188.250 579.060 1188.570 579.120 ;
        RECT 1187.330 386.480 1187.650 386.540 ;
        RECT 1187.790 386.480 1188.110 386.540 ;
        RECT 1187.330 386.340 1188.110 386.480 ;
        RECT 1187.330 386.280 1187.650 386.340 ;
        RECT 1187.790 386.280 1188.110 386.340 ;
        RECT 1187.790 337.860 1188.110 337.920 ;
        RECT 1188.250 337.860 1188.570 337.920 ;
        RECT 1187.790 337.720 1188.570 337.860 ;
        RECT 1187.790 337.660 1188.110 337.720 ;
        RECT 1188.250 337.660 1188.570 337.720 ;
        RECT 1187.790 241.300 1188.110 241.360 ;
        RECT 1188.250 241.300 1188.570 241.360 ;
        RECT 1187.790 241.160 1188.570 241.300 ;
        RECT 1187.790 241.100 1188.110 241.160 ;
        RECT 1188.250 241.100 1188.570 241.160 ;
        RECT 1187.330 96.800 1187.650 96.860 ;
        RECT 1187.790 96.800 1188.110 96.860 ;
        RECT 1187.330 96.660 1188.110 96.800 ;
        RECT 1187.330 96.600 1187.650 96.660 ;
        RECT 1187.790 96.600 1188.110 96.660 ;
        RECT 858.890 32.200 859.210 32.260 ;
        RECT 1187.790 32.200 1188.110 32.260 ;
        RECT 858.890 32.060 1188.110 32.200 ;
        RECT 858.890 32.000 859.210 32.060 ;
        RECT 1187.790 32.000 1188.110 32.060 ;
      LAYER via ;
        RECT 1188.740 1196.840 1189.000 1197.100 ;
        RECT 1188.280 1159.100 1188.540 1159.360 ;
        RECT 1187.820 965.980 1188.080 966.240 ;
        RECT 1188.740 965.980 1189.000 966.240 ;
        RECT 1187.820 869.420 1188.080 869.680 ;
        RECT 1188.740 869.420 1189.000 869.680 ;
        RECT 1187.820 820.800 1188.080 821.060 ;
        RECT 1187.820 786.120 1188.080 786.380 ;
        RECT 1187.820 724.240 1188.080 724.500 ;
        RECT 1188.280 724.240 1188.540 724.500 ;
        RECT 1187.820 579.400 1188.080 579.660 ;
        RECT 1188.280 579.060 1188.540 579.320 ;
        RECT 1187.360 386.280 1187.620 386.540 ;
        RECT 1187.820 386.280 1188.080 386.540 ;
        RECT 1187.820 337.660 1188.080 337.920 ;
        RECT 1188.280 337.660 1188.540 337.920 ;
        RECT 1187.820 241.100 1188.080 241.360 ;
        RECT 1188.280 241.100 1188.540 241.360 ;
        RECT 1187.360 96.600 1187.620 96.860 ;
        RECT 1187.820 96.600 1188.080 96.860 ;
        RECT 858.920 32.000 859.180 32.260 ;
        RECT 1187.820 32.000 1188.080 32.260 ;
      LAYER met2 ;
        RECT 1191.050 1221.010 1191.610 1228.680 ;
        RECT 1188.800 1220.870 1191.610 1221.010 ;
        RECT 1188.800 1197.130 1188.940 1220.870 ;
        RECT 1191.050 1219.680 1191.610 1220.870 ;
        RECT 1188.740 1196.810 1189.000 1197.130 ;
        RECT 1188.280 1159.070 1188.540 1159.390 ;
        RECT 1188.340 1076.850 1188.480 1159.070 ;
        RECT 1187.880 1076.710 1188.480 1076.850 ;
        RECT 1187.880 1038.770 1188.020 1076.710 ;
        RECT 1187.880 1038.630 1188.480 1038.770 ;
        RECT 1188.340 990.490 1188.480 1038.630 ;
        RECT 1188.340 990.350 1188.940 990.490 ;
        RECT 1188.800 966.270 1188.940 990.350 ;
        RECT 1187.820 966.010 1188.080 966.270 ;
        RECT 1187.820 965.950 1188.480 966.010 ;
        RECT 1188.740 965.950 1189.000 966.270 ;
        RECT 1187.880 965.870 1188.480 965.950 ;
        RECT 1188.340 893.930 1188.480 965.870 ;
        RECT 1188.340 893.790 1188.940 893.930 ;
        RECT 1188.800 869.710 1188.940 893.790 ;
        RECT 1187.820 869.390 1188.080 869.710 ;
        RECT 1188.740 869.390 1189.000 869.710 ;
        RECT 1187.880 821.090 1188.020 869.390 ;
        RECT 1187.820 820.770 1188.080 821.090 ;
        RECT 1187.820 786.090 1188.080 786.410 ;
        RECT 1187.880 748.410 1188.020 786.090 ;
        RECT 1187.880 748.270 1188.480 748.410 ;
        RECT 1188.340 724.530 1188.480 748.270 ;
        RECT 1187.820 724.210 1188.080 724.530 ;
        RECT 1188.280 724.210 1188.540 724.530 ;
        RECT 1187.880 651.850 1188.020 724.210 ;
        RECT 1187.880 651.710 1188.480 651.850 ;
        RECT 1188.340 580.565 1188.480 651.710 ;
        RECT 1188.270 580.195 1188.550 580.565 ;
        RECT 1187.810 579.515 1188.090 579.885 ;
        RECT 1187.820 579.370 1188.080 579.515 ;
        RECT 1188.280 579.030 1188.540 579.350 ;
        RECT 1188.340 507.010 1188.480 579.030 ;
        RECT 1187.880 506.870 1188.480 507.010 ;
        RECT 1187.880 435.725 1188.020 506.870 ;
        RECT 1187.810 435.355 1188.090 435.725 ;
        RECT 1187.350 434.675 1187.630 435.045 ;
        RECT 1187.420 386.570 1187.560 434.675 ;
        RECT 1187.360 386.250 1187.620 386.570 ;
        RECT 1187.820 386.250 1188.080 386.570 ;
        RECT 1187.880 337.950 1188.020 386.250 ;
        RECT 1187.820 337.630 1188.080 337.950 ;
        RECT 1188.280 337.630 1188.540 337.950 ;
        RECT 1188.340 241.390 1188.480 337.630 ;
        RECT 1187.820 241.070 1188.080 241.390 ;
        RECT 1188.280 241.070 1188.540 241.390 ;
        RECT 1187.880 169.050 1188.020 241.070 ;
        RECT 1187.420 168.910 1188.020 169.050 ;
        RECT 1187.420 96.890 1187.560 168.910 ;
        RECT 1187.360 96.570 1187.620 96.890 ;
        RECT 1187.820 96.570 1188.080 96.890 ;
        RECT 1187.880 32.290 1188.020 96.570 ;
        RECT 858.920 31.970 859.180 32.290 ;
        RECT 1187.820 31.970 1188.080 32.290 ;
        RECT 858.980 2.400 859.120 31.970 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 1188.270 580.240 1188.550 580.520 ;
        RECT 1187.810 579.560 1188.090 579.840 ;
        RECT 1187.810 435.400 1188.090 435.680 ;
        RECT 1187.350 434.720 1187.630 435.000 ;
      LAYER met3 ;
        RECT 1188.245 580.530 1188.575 580.545 ;
        RECT 1188.030 580.215 1188.575 580.530 ;
        RECT 1188.030 579.865 1188.330 580.215 ;
        RECT 1187.785 579.550 1188.330 579.865 ;
        RECT 1187.785 579.535 1188.115 579.550 ;
        RECT 1187.785 435.690 1188.115 435.705 ;
        RECT 1187.110 435.390 1188.115 435.690 ;
        RECT 1187.110 435.025 1187.410 435.390 ;
        RECT 1187.785 435.375 1188.115 435.390 ;
        RECT 1187.110 434.710 1187.655 435.025 ;
        RECT 1187.325 434.695 1187.655 434.710 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1195.610 1159.300 1195.930 1159.360 ;
        RECT 1198.370 1159.300 1198.690 1159.360 ;
        RECT 1195.610 1159.160 1198.690 1159.300 ;
        RECT 1195.610 1159.100 1195.930 1159.160 ;
        RECT 1198.370 1159.100 1198.690 1159.160 ;
        RECT 1195.150 966.180 1195.470 966.240 ;
        RECT 1196.070 966.180 1196.390 966.240 ;
        RECT 1195.150 966.040 1196.390 966.180 ;
        RECT 1195.150 965.980 1195.470 966.040 ;
        RECT 1196.070 965.980 1196.390 966.040 ;
        RECT 1195.150 869.620 1195.470 869.680 ;
        RECT 1196.070 869.620 1196.390 869.680 ;
        RECT 1195.150 869.480 1196.390 869.620 ;
        RECT 1195.150 869.420 1195.470 869.480 ;
        RECT 1196.070 869.420 1196.390 869.480 ;
        RECT 1195.150 821.000 1195.470 821.060 ;
        RECT 1195.610 821.000 1195.930 821.060 ;
        RECT 1195.150 820.860 1195.930 821.000 ;
        RECT 1195.150 820.800 1195.470 820.860 ;
        RECT 1195.610 820.800 1195.930 820.860 ;
        RECT 1195.150 772.520 1195.470 772.780 ;
        RECT 1195.240 772.380 1195.380 772.520 ;
        RECT 1195.610 772.380 1195.930 772.440 ;
        RECT 1195.240 772.240 1195.930 772.380 ;
        RECT 1195.610 772.180 1195.930 772.240 ;
        RECT 1195.150 724.440 1195.470 724.500 ;
        RECT 1195.610 724.440 1195.930 724.500 ;
        RECT 1195.150 724.300 1195.930 724.440 ;
        RECT 1195.150 724.240 1195.470 724.300 ;
        RECT 1195.610 724.240 1195.930 724.300 ;
        RECT 1194.690 627.880 1195.010 627.940 ;
        RECT 1195.610 627.880 1195.930 627.940 ;
        RECT 1194.690 627.740 1195.930 627.880 ;
        RECT 1194.690 627.680 1195.010 627.740 ;
        RECT 1195.610 627.680 1195.930 627.740 ;
        RECT 1195.150 96.800 1195.470 96.860 ;
        RECT 1195.610 96.800 1195.930 96.860 ;
        RECT 1195.150 96.660 1195.930 96.800 ;
        RECT 1195.150 96.600 1195.470 96.660 ;
        RECT 1195.610 96.600 1195.930 96.660 ;
        RECT 876.830 32.540 877.150 32.600 ;
        RECT 1195.150 32.540 1195.470 32.600 ;
        RECT 876.830 32.400 1195.470 32.540 ;
        RECT 876.830 32.340 877.150 32.400 ;
        RECT 1195.150 32.340 1195.470 32.400 ;
      LAYER via ;
        RECT 1195.640 1159.100 1195.900 1159.360 ;
        RECT 1198.400 1159.100 1198.660 1159.360 ;
        RECT 1195.180 965.980 1195.440 966.240 ;
        RECT 1196.100 965.980 1196.360 966.240 ;
        RECT 1195.180 869.420 1195.440 869.680 ;
        RECT 1196.100 869.420 1196.360 869.680 ;
        RECT 1195.180 820.800 1195.440 821.060 ;
        RECT 1195.640 820.800 1195.900 821.060 ;
        RECT 1195.180 772.520 1195.440 772.780 ;
        RECT 1195.640 772.180 1195.900 772.440 ;
        RECT 1195.180 724.240 1195.440 724.500 ;
        RECT 1195.640 724.240 1195.900 724.500 ;
        RECT 1194.720 627.680 1194.980 627.940 ;
        RECT 1195.640 627.680 1195.900 627.940 ;
        RECT 1195.180 96.600 1195.440 96.860 ;
        RECT 1195.640 96.600 1195.900 96.860 ;
        RECT 876.860 32.340 877.120 32.600 ;
        RECT 1195.180 32.340 1195.440 32.600 ;
      LAYER met2 ;
        RECT 1200.250 1220.330 1200.810 1228.680 ;
        RECT 1198.460 1220.190 1200.810 1220.330 ;
        RECT 1198.460 1159.390 1198.600 1220.190 ;
        RECT 1200.250 1219.680 1200.810 1220.190 ;
        RECT 1195.640 1159.070 1195.900 1159.390 ;
        RECT 1198.400 1159.070 1198.660 1159.390 ;
        RECT 1195.700 1076.850 1195.840 1159.070 ;
        RECT 1195.240 1076.710 1195.840 1076.850 ;
        RECT 1195.240 1027.890 1195.380 1076.710 ;
        RECT 1195.240 1027.750 1195.840 1027.890 ;
        RECT 1195.700 990.490 1195.840 1027.750 ;
        RECT 1195.700 990.350 1196.300 990.490 ;
        RECT 1196.160 966.270 1196.300 990.350 ;
        RECT 1195.180 966.125 1195.440 966.270 ;
        RECT 1196.100 966.125 1196.360 966.270 ;
        RECT 1195.170 965.755 1195.450 966.125 ;
        RECT 1196.090 965.755 1196.370 966.125 ;
        RECT 1196.160 931.330 1196.300 965.755 ;
        RECT 1195.700 931.190 1196.300 931.330 ;
        RECT 1195.700 893.930 1195.840 931.190 ;
        RECT 1195.700 893.790 1196.300 893.930 ;
        RECT 1196.160 869.710 1196.300 893.790 ;
        RECT 1195.180 869.390 1195.440 869.710 ;
        RECT 1196.100 869.390 1196.360 869.710 ;
        RECT 1195.240 821.090 1195.380 869.390 ;
        RECT 1195.180 820.770 1195.440 821.090 ;
        RECT 1195.640 820.770 1195.900 821.090 ;
        RECT 1195.700 796.010 1195.840 820.770 ;
        RECT 1195.240 795.870 1195.840 796.010 ;
        RECT 1195.240 772.810 1195.380 795.870 ;
        RECT 1195.180 772.490 1195.440 772.810 ;
        RECT 1195.640 772.150 1195.900 772.470 ;
        RECT 1195.700 724.530 1195.840 772.150 ;
        RECT 1195.180 724.210 1195.440 724.530 ;
        RECT 1195.640 724.210 1195.900 724.530 ;
        RECT 1195.240 651.850 1195.380 724.210 ;
        RECT 1195.240 651.710 1196.300 651.850 ;
        RECT 1196.160 641.650 1196.300 651.710 ;
        RECT 1195.700 641.510 1196.300 641.650 ;
        RECT 1195.700 627.970 1195.840 641.510 ;
        RECT 1194.720 627.650 1194.980 627.970 ;
        RECT 1195.640 627.650 1195.900 627.970 ;
        RECT 1194.780 593.370 1194.920 627.650 ;
        RECT 1194.780 593.230 1195.380 593.370 ;
        RECT 1195.240 555.290 1195.380 593.230 ;
        RECT 1195.240 555.150 1195.840 555.290 ;
        RECT 1195.700 507.010 1195.840 555.150 ;
        RECT 1195.240 506.870 1195.840 507.010 ;
        RECT 1195.240 254.730 1195.380 506.870 ;
        RECT 1195.240 254.590 1195.840 254.730 ;
        RECT 1195.700 96.890 1195.840 254.590 ;
        RECT 1195.180 96.570 1195.440 96.890 ;
        RECT 1195.640 96.570 1195.900 96.890 ;
        RECT 1195.240 32.630 1195.380 96.570 ;
        RECT 876.860 32.310 877.120 32.630 ;
        RECT 1195.180 32.310 1195.440 32.630 ;
        RECT 876.920 2.400 877.060 32.310 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1195.170 965.800 1195.450 966.080 ;
        RECT 1196.090 965.800 1196.370 966.080 ;
      LAYER met3 ;
        RECT 1195.145 966.090 1195.475 966.105 ;
        RECT 1196.065 966.090 1196.395 966.105 ;
        RECT 1195.145 965.790 1196.395 966.090 ;
        RECT 1195.145 965.775 1195.475 965.790 ;
        RECT 1196.065 965.775 1196.395 965.790 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 32.880 895.090 32.940 ;
        RECT 1208.030 32.880 1208.350 32.940 ;
        RECT 894.770 32.740 1208.350 32.880 ;
        RECT 894.770 32.680 895.090 32.740 ;
        RECT 1208.030 32.680 1208.350 32.740 ;
      LAYER via ;
        RECT 894.800 32.680 895.060 32.940 ;
        RECT 1208.060 32.680 1208.320 32.940 ;
      LAYER met2 ;
        RECT 1209.450 1220.330 1210.010 1228.680 ;
        RECT 1208.120 1220.190 1210.010 1220.330 ;
        RECT 1208.120 32.970 1208.260 1220.190 ;
        RECT 1209.450 1219.680 1210.010 1220.190 ;
        RECT 894.800 32.650 895.060 32.970 ;
        RECT 1208.060 32.650 1208.320 32.970 ;
        RECT 894.860 2.400 895.000 32.650 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1010.690 1210.300 1011.010 1210.360 ;
        RECT 1218.610 1210.300 1218.930 1210.360 ;
        RECT 1010.690 1210.160 1218.930 1210.300 ;
        RECT 1010.690 1210.100 1011.010 1210.160 ;
        RECT 1218.610 1210.100 1218.930 1210.160 ;
        RECT 912.710 19.620 913.030 19.680 ;
        RECT 1010.690 19.620 1011.010 19.680 ;
        RECT 912.710 19.480 1011.010 19.620 ;
        RECT 912.710 19.420 913.030 19.480 ;
        RECT 1010.690 19.420 1011.010 19.480 ;
      LAYER via ;
        RECT 1010.720 1210.100 1010.980 1210.360 ;
        RECT 1218.640 1210.100 1218.900 1210.360 ;
        RECT 912.740 19.420 913.000 19.680 ;
        RECT 1010.720 19.420 1010.980 19.680 ;
      LAYER met2 ;
        RECT 1218.650 1219.680 1219.210 1228.680 ;
        RECT 1218.700 1210.390 1218.840 1219.680 ;
        RECT 1010.720 1210.070 1010.980 1210.390 ;
        RECT 1218.640 1210.070 1218.900 1210.390 ;
        RECT 1010.780 19.710 1010.920 1210.070 ;
        RECT 912.740 19.390 913.000 19.710 ;
        RECT 1010.720 19.390 1010.980 19.710 ;
        RECT 912.800 2.400 912.940 19.390 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 996.890 1213.700 997.210 1213.760 ;
        RECT 1227.810 1213.700 1228.130 1213.760 ;
        RECT 996.890 1213.560 1228.130 1213.700 ;
        RECT 996.890 1213.500 997.210 1213.560 ;
        RECT 1227.810 1213.500 1228.130 1213.560 ;
        RECT 930.190 19.960 930.510 20.020 ;
        RECT 996.890 19.960 997.210 20.020 ;
        RECT 930.190 19.820 997.210 19.960 ;
        RECT 930.190 19.760 930.510 19.820 ;
        RECT 996.890 19.760 997.210 19.820 ;
      LAYER via ;
        RECT 996.920 1213.500 997.180 1213.760 ;
        RECT 1227.840 1213.500 1228.100 1213.760 ;
        RECT 930.220 19.760 930.480 20.020 ;
        RECT 996.920 19.760 997.180 20.020 ;
      LAYER met2 ;
        RECT 1227.850 1219.680 1228.410 1228.680 ;
        RECT 1227.900 1213.790 1228.040 1219.680 ;
        RECT 996.920 1213.470 997.180 1213.790 ;
        RECT 1227.840 1213.470 1228.100 1213.790 ;
        RECT 996.980 20.050 997.120 1213.470 ;
        RECT 930.220 19.730 930.480 20.050 ;
        RECT 996.920 19.730 997.180 20.050 ;
        RECT 930.280 2.400 930.420 19.730 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 991.445 1159.145 991.615 1207.255 ;
        RECT 991.445 745.365 991.615 793.475 ;
        RECT 990.985 269.025 991.155 317.475 ;
      LAYER mcon ;
        RECT 991.445 1207.085 991.615 1207.255 ;
        RECT 991.445 793.305 991.615 793.475 ;
        RECT 990.985 317.305 991.155 317.475 ;
      LAYER met1 ;
        RECT 991.370 1212.340 991.690 1212.400 ;
        RECT 1237.010 1212.340 1237.330 1212.400 ;
        RECT 991.370 1212.200 1237.330 1212.340 ;
        RECT 991.370 1212.140 991.690 1212.200 ;
        RECT 1237.010 1212.140 1237.330 1212.200 ;
        RECT 991.370 1207.240 991.690 1207.300 ;
        RECT 991.175 1207.100 991.690 1207.240 ;
        RECT 991.370 1207.040 991.690 1207.100 ;
        RECT 991.370 1159.300 991.690 1159.360 ;
        RECT 991.175 1159.160 991.690 1159.300 ;
        RECT 991.370 1159.100 991.690 1159.160 ;
        RECT 991.370 1124.760 991.690 1125.020 ;
        RECT 991.460 1124.280 991.600 1124.760 ;
        RECT 991.830 1124.280 992.150 1124.340 ;
        RECT 991.460 1124.140 992.150 1124.280 ;
        RECT 991.830 1124.080 992.150 1124.140 ;
        RECT 990.910 1055.600 991.230 1055.660 ;
        RECT 991.830 1055.600 992.150 1055.660 ;
        RECT 990.910 1055.460 992.150 1055.600 ;
        RECT 990.910 1055.400 991.230 1055.460 ;
        RECT 991.830 1055.400 992.150 1055.460 ;
        RECT 991.830 1007.800 992.150 1008.060 ;
        RECT 991.920 1007.380 992.060 1007.800 ;
        RECT 991.830 1007.120 992.150 1007.380 ;
        RECT 991.370 945.440 991.690 945.500 ;
        RECT 991.830 945.440 992.150 945.500 ;
        RECT 991.370 945.300 992.150 945.440 ;
        RECT 991.370 945.240 991.690 945.300 ;
        RECT 991.830 945.240 992.150 945.300 ;
        RECT 991.370 814.200 991.690 814.260 ;
        RECT 991.830 814.200 992.150 814.260 ;
        RECT 991.370 814.060 992.150 814.200 ;
        RECT 991.370 814.000 991.690 814.060 ;
        RECT 991.830 814.000 992.150 814.060 ;
        RECT 991.385 793.460 991.675 793.505 ;
        RECT 991.830 793.460 992.150 793.520 ;
        RECT 991.385 793.320 992.150 793.460 ;
        RECT 991.385 793.275 991.675 793.320 ;
        RECT 991.830 793.260 992.150 793.320 ;
        RECT 991.370 745.520 991.690 745.580 ;
        RECT 991.175 745.380 991.690 745.520 ;
        RECT 991.370 745.320 991.690 745.380 ;
        RECT 991.370 690.240 991.690 690.500 ;
        RECT 991.460 689.820 991.600 690.240 ;
        RECT 991.370 689.560 991.690 689.820 ;
        RECT 991.370 493.380 991.690 493.640 ;
        RECT 991.460 492.960 991.600 493.380 ;
        RECT 991.370 492.700 991.690 492.960 ;
        RECT 991.370 380.020 991.690 380.080 ;
        RECT 991.000 379.880 991.690 380.020 ;
        RECT 991.000 379.740 991.140 379.880 ;
        RECT 991.370 379.820 991.690 379.880 ;
        RECT 990.910 379.480 991.230 379.740 ;
        RECT 990.910 372.540 991.230 372.600 ;
        RECT 991.370 372.540 991.690 372.600 ;
        RECT 990.910 372.400 991.690 372.540 ;
        RECT 990.910 372.340 991.230 372.400 ;
        RECT 991.370 372.340 991.690 372.400 ;
        RECT 990.910 317.460 991.230 317.520 ;
        RECT 990.715 317.320 991.230 317.460 ;
        RECT 990.910 317.260 991.230 317.320 ;
        RECT 990.910 269.180 991.230 269.240 ;
        RECT 990.715 269.040 991.230 269.180 ;
        RECT 990.910 268.980 991.230 269.040 ;
        RECT 990.910 138.280 991.230 138.340 ;
        RECT 991.370 138.280 991.690 138.340 ;
        RECT 990.910 138.140 991.690 138.280 ;
        RECT 990.910 138.080 991.230 138.140 ;
        RECT 991.370 138.080 991.690 138.140 ;
        RECT 991.370 110.740 991.690 110.800 ;
        RECT 991.000 110.600 991.690 110.740 ;
        RECT 991.000 110.460 991.140 110.600 ;
        RECT 991.370 110.540 991.690 110.600 ;
        RECT 990.910 110.200 991.230 110.460 ;
        RECT 948.130 20.300 948.450 20.360 ;
        RECT 990.910 20.300 991.230 20.360 ;
        RECT 948.130 20.160 991.230 20.300 ;
        RECT 948.130 20.100 948.450 20.160 ;
        RECT 990.910 20.100 991.230 20.160 ;
      LAYER via ;
        RECT 991.400 1212.140 991.660 1212.400 ;
        RECT 1237.040 1212.140 1237.300 1212.400 ;
        RECT 991.400 1207.040 991.660 1207.300 ;
        RECT 991.400 1159.100 991.660 1159.360 ;
        RECT 991.400 1124.760 991.660 1125.020 ;
        RECT 991.860 1124.080 992.120 1124.340 ;
        RECT 990.940 1055.400 991.200 1055.660 ;
        RECT 991.860 1055.400 992.120 1055.660 ;
        RECT 991.860 1007.800 992.120 1008.060 ;
        RECT 991.860 1007.120 992.120 1007.380 ;
        RECT 991.400 945.240 991.660 945.500 ;
        RECT 991.860 945.240 992.120 945.500 ;
        RECT 991.400 814.000 991.660 814.260 ;
        RECT 991.860 814.000 992.120 814.260 ;
        RECT 991.860 793.260 992.120 793.520 ;
        RECT 991.400 745.320 991.660 745.580 ;
        RECT 991.400 690.240 991.660 690.500 ;
        RECT 991.400 689.560 991.660 689.820 ;
        RECT 991.400 493.380 991.660 493.640 ;
        RECT 991.400 492.700 991.660 492.960 ;
        RECT 991.400 379.820 991.660 380.080 ;
        RECT 990.940 379.480 991.200 379.740 ;
        RECT 990.940 372.340 991.200 372.600 ;
        RECT 991.400 372.340 991.660 372.600 ;
        RECT 990.940 317.260 991.200 317.520 ;
        RECT 990.940 268.980 991.200 269.240 ;
        RECT 990.940 138.080 991.200 138.340 ;
        RECT 991.400 138.080 991.660 138.340 ;
        RECT 991.400 110.540 991.660 110.800 ;
        RECT 990.940 110.200 991.200 110.460 ;
        RECT 948.160 20.100 948.420 20.360 ;
        RECT 990.940 20.100 991.200 20.360 ;
      LAYER met2 ;
        RECT 1237.050 1219.680 1237.610 1228.680 ;
        RECT 1237.100 1212.430 1237.240 1219.680 ;
        RECT 991.400 1212.110 991.660 1212.430 ;
        RECT 1237.040 1212.110 1237.300 1212.430 ;
        RECT 991.460 1207.330 991.600 1212.110 ;
        RECT 991.400 1207.010 991.660 1207.330 ;
        RECT 991.400 1159.070 991.660 1159.390 ;
        RECT 991.460 1125.050 991.600 1159.070 ;
        RECT 991.400 1124.730 991.660 1125.050 ;
        RECT 991.860 1124.050 992.120 1124.370 ;
        RECT 991.920 1055.885 992.060 1124.050 ;
        RECT 990.930 1055.515 991.210 1055.885 ;
        RECT 991.850 1055.515 992.130 1055.885 ;
        RECT 990.940 1055.370 991.200 1055.515 ;
        RECT 991.860 1055.370 992.120 1055.515 ;
        RECT 991.920 1008.090 992.060 1055.370 ;
        RECT 991.860 1007.770 992.120 1008.090 ;
        RECT 991.860 1007.090 992.120 1007.410 ;
        RECT 991.920 945.530 992.060 1007.090 ;
        RECT 991.400 945.210 991.660 945.530 ;
        RECT 991.860 945.210 992.120 945.530 ;
        RECT 991.460 814.290 991.600 945.210 ;
        RECT 991.400 813.970 991.660 814.290 ;
        RECT 991.860 813.970 992.120 814.290 ;
        RECT 991.920 793.550 992.060 813.970 ;
        RECT 991.860 793.230 992.120 793.550 ;
        RECT 991.400 745.290 991.660 745.610 ;
        RECT 991.460 690.530 991.600 745.290 ;
        RECT 991.400 690.210 991.660 690.530 ;
        RECT 991.400 689.530 991.660 689.850 ;
        RECT 991.460 566.170 991.600 689.530 ;
        RECT 991.000 566.030 991.600 566.170 ;
        RECT 991.000 545.770 991.140 566.030 ;
        RECT 991.000 545.630 992.060 545.770 ;
        RECT 991.920 544.410 992.060 545.630 ;
        RECT 991.460 544.270 992.060 544.410 ;
        RECT 991.460 493.670 991.600 544.270 ;
        RECT 991.400 493.350 991.660 493.670 ;
        RECT 991.400 492.670 991.660 492.990 ;
        RECT 991.460 380.110 991.600 492.670 ;
        RECT 991.400 379.790 991.660 380.110 ;
        RECT 990.940 379.450 991.200 379.770 ;
        RECT 991.000 372.630 991.140 379.450 ;
        RECT 990.940 372.310 991.200 372.630 ;
        RECT 991.400 372.310 991.660 372.630 ;
        RECT 991.460 324.770 991.600 372.310 ;
        RECT 991.000 324.630 991.600 324.770 ;
        RECT 991.000 317.550 991.140 324.630 ;
        RECT 990.940 317.230 991.200 317.550 ;
        RECT 990.940 268.950 991.200 269.270 ;
        RECT 991.000 252.010 991.140 268.950 ;
        RECT 991.000 251.870 991.600 252.010 ;
        RECT 991.460 203.730 991.600 251.870 ;
        RECT 991.000 203.590 991.600 203.730 ;
        RECT 991.000 138.370 991.140 203.590 ;
        RECT 990.940 138.050 991.200 138.370 ;
        RECT 991.400 138.050 991.660 138.370 ;
        RECT 991.460 110.830 991.600 138.050 ;
        RECT 991.400 110.510 991.660 110.830 ;
        RECT 990.940 110.170 991.200 110.490 ;
        RECT 991.000 73.170 991.140 110.170 ;
        RECT 991.000 73.030 991.600 73.170 ;
        RECT 991.460 71.810 991.600 73.030 ;
        RECT 991.000 71.670 991.600 71.810 ;
        RECT 991.000 20.390 991.140 71.670 ;
        RECT 948.160 20.070 948.420 20.390 ;
        RECT 990.940 20.070 991.200 20.390 ;
        RECT 948.220 2.400 948.360 20.070 ;
        RECT 948.010 -4.800 948.570 2.400 ;
      LAYER via2 ;
        RECT 990.930 1055.560 991.210 1055.840 ;
        RECT 991.850 1055.560 992.130 1055.840 ;
      LAYER met3 ;
        RECT 990.905 1055.850 991.235 1055.865 ;
        RECT 991.825 1055.850 992.155 1055.865 ;
        RECT 990.905 1055.550 992.155 1055.850 ;
        RECT 990.905 1055.535 991.235 1055.550 ;
        RECT 991.825 1055.535 992.155 1055.550 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1192.465 1210.825 1192.635 1211.675 ;
      LAYER mcon ;
        RECT 1192.465 1211.505 1192.635 1211.675 ;
      LAYER met1 ;
        RECT 990.910 1211.660 991.230 1211.720 ;
        RECT 1192.405 1211.660 1192.695 1211.705 ;
        RECT 990.910 1211.520 1192.695 1211.660 ;
        RECT 990.910 1211.460 991.230 1211.520 ;
        RECT 1192.405 1211.475 1192.695 1211.520 ;
        RECT 1192.405 1210.980 1192.695 1211.025 ;
        RECT 1245.750 1210.980 1246.070 1211.040 ;
        RECT 1192.405 1210.840 1246.070 1210.980 ;
        RECT 1192.405 1210.795 1192.695 1210.840 ;
        RECT 1245.750 1210.780 1246.070 1210.840 ;
        RECT 966.070 15.200 966.390 15.260 ;
        RECT 989.990 15.200 990.310 15.260 ;
        RECT 966.070 15.060 990.310 15.200 ;
        RECT 966.070 15.000 966.390 15.060 ;
        RECT 989.990 15.000 990.310 15.060 ;
      LAYER via ;
        RECT 990.940 1211.460 991.200 1211.720 ;
        RECT 1245.780 1210.780 1246.040 1211.040 ;
        RECT 966.100 15.000 966.360 15.260 ;
        RECT 990.020 15.000 990.280 15.260 ;
      LAYER met2 ;
        RECT 1245.790 1219.680 1246.350 1228.680 ;
        RECT 990.940 1211.430 991.200 1211.750 ;
        RECT 991.000 1192.450 991.140 1211.430 ;
        RECT 1245.840 1211.070 1245.980 1219.680 ;
        RECT 1245.780 1210.750 1246.040 1211.070 ;
        RECT 990.080 1192.310 991.140 1192.450 ;
        RECT 990.080 15.290 990.220 1192.310 ;
        RECT 966.100 14.970 966.360 15.290 ;
        RECT 990.020 14.970 990.280 15.290 ;
        RECT 966.160 2.400 966.300 14.970 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1192.005 1207.765 1192.175 1210.995 ;
      LAYER mcon ;
        RECT 1192.005 1210.825 1192.175 1210.995 ;
      LAYER met1 ;
        RECT 986.310 1210.980 986.630 1211.040 ;
        RECT 1191.945 1210.980 1192.235 1211.025 ;
        RECT 986.310 1210.840 1192.235 1210.980 ;
        RECT 986.310 1210.780 986.630 1210.840 ;
        RECT 1191.945 1210.795 1192.235 1210.840 ;
        RECT 1191.945 1207.920 1192.235 1207.965 ;
        RECT 1254.950 1207.920 1255.270 1207.980 ;
        RECT 1191.945 1207.780 1255.270 1207.920 ;
        RECT 1191.945 1207.735 1192.235 1207.780 ;
        RECT 1254.950 1207.720 1255.270 1207.780 ;
        RECT 984.010 20.640 984.330 20.700 ;
        RECT 986.310 20.640 986.630 20.700 ;
        RECT 984.010 20.500 986.630 20.640 ;
        RECT 984.010 20.440 984.330 20.500 ;
        RECT 986.310 20.440 986.630 20.500 ;
      LAYER via ;
        RECT 986.340 1210.780 986.600 1211.040 ;
        RECT 1254.980 1207.720 1255.240 1207.980 ;
        RECT 984.040 20.440 984.300 20.700 ;
        RECT 986.340 20.440 986.600 20.700 ;
      LAYER met2 ;
        RECT 1254.990 1219.680 1255.550 1228.680 ;
        RECT 986.340 1210.750 986.600 1211.070 ;
        RECT 986.400 20.730 986.540 1210.750 ;
        RECT 1255.040 1208.010 1255.180 1219.680 ;
        RECT 1254.980 1207.690 1255.240 1208.010 ;
        RECT 984.040 20.410 984.300 20.730 ;
        RECT 986.340 20.410 986.600 20.730 ;
        RECT 984.100 2.400 984.240 20.410 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 30.160 663.250 30.220 ;
        RECT 1090.270 30.160 1090.590 30.220 ;
        RECT 662.930 30.020 1090.590 30.160 ;
        RECT 662.930 29.960 663.250 30.020 ;
        RECT 1090.270 29.960 1090.590 30.020 ;
      LAYER via ;
        RECT 662.960 29.960 663.220 30.220 ;
        RECT 1090.300 29.960 1090.560 30.220 ;
      LAYER met2 ;
        RECT 1090.310 1219.680 1090.870 1228.680 ;
        RECT 1090.360 30.250 1090.500 1219.680 ;
        RECT 662.960 29.930 663.220 30.250 ;
        RECT 1090.300 29.930 1090.560 30.250 ;
        RECT 663.020 2.400 663.160 29.930 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 1211.320 1007.330 1211.380 ;
        RECT 1264.150 1211.320 1264.470 1211.380 ;
        RECT 1007.010 1211.180 1264.470 1211.320 ;
        RECT 1007.010 1211.120 1007.330 1211.180 ;
        RECT 1264.150 1211.120 1264.470 1211.180 ;
        RECT 1001.950 16.900 1002.270 16.960 ;
        RECT 1007.010 16.900 1007.330 16.960 ;
        RECT 1001.950 16.760 1007.330 16.900 ;
        RECT 1001.950 16.700 1002.270 16.760 ;
        RECT 1007.010 16.700 1007.330 16.760 ;
      LAYER via ;
        RECT 1007.040 1211.120 1007.300 1211.380 ;
        RECT 1264.180 1211.120 1264.440 1211.380 ;
        RECT 1001.980 16.700 1002.240 16.960 ;
        RECT 1007.040 16.700 1007.300 16.960 ;
      LAYER met2 ;
        RECT 1264.190 1219.680 1264.750 1228.680 ;
        RECT 1264.240 1211.410 1264.380 1219.680 ;
        RECT 1007.040 1211.090 1007.300 1211.410 ;
        RECT 1264.180 1211.090 1264.440 1211.410 ;
        RECT 1007.100 16.990 1007.240 1211.090 ;
        RECT 1001.980 16.670 1002.240 16.990 ;
        RECT 1007.040 16.670 1007.300 16.990 ;
        RECT 1002.040 2.400 1002.180 16.670 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1020.810 1212.000 1021.130 1212.060 ;
        RECT 1273.350 1212.000 1273.670 1212.060 ;
        RECT 1020.810 1211.860 1273.670 1212.000 ;
        RECT 1020.810 1211.800 1021.130 1211.860 ;
        RECT 1273.350 1211.800 1273.670 1211.860 ;
      LAYER via ;
        RECT 1020.840 1211.800 1021.100 1212.060 ;
        RECT 1273.380 1211.800 1273.640 1212.060 ;
      LAYER met2 ;
        RECT 1273.390 1219.680 1273.950 1228.680 ;
        RECT 1273.440 1212.090 1273.580 1219.680 ;
        RECT 1020.840 1211.770 1021.100 1212.090 ;
        RECT 1273.380 1211.770 1273.640 1212.090 ;
        RECT 1020.900 3.130 1021.040 1211.770 ;
        RECT 1019.520 2.990 1021.040 3.130 ;
        RECT 1019.520 2.400 1019.660 2.990 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 1213.020 1041.830 1213.080 ;
        RECT 1282.550 1213.020 1282.870 1213.080 ;
        RECT 1041.510 1212.880 1282.870 1213.020 ;
        RECT 1041.510 1212.820 1041.830 1212.880 ;
        RECT 1282.550 1212.820 1282.870 1212.880 ;
        RECT 1037.370 20.640 1037.690 20.700 ;
        RECT 1041.510 20.640 1041.830 20.700 ;
        RECT 1037.370 20.500 1041.830 20.640 ;
        RECT 1037.370 20.440 1037.690 20.500 ;
        RECT 1041.510 20.440 1041.830 20.500 ;
      LAYER via ;
        RECT 1041.540 1212.820 1041.800 1213.080 ;
        RECT 1282.580 1212.820 1282.840 1213.080 ;
        RECT 1037.400 20.440 1037.660 20.700 ;
        RECT 1041.540 20.440 1041.800 20.700 ;
      LAYER met2 ;
        RECT 1282.590 1219.680 1283.150 1228.680 ;
        RECT 1282.640 1213.110 1282.780 1219.680 ;
        RECT 1041.540 1212.790 1041.800 1213.110 ;
        RECT 1282.580 1212.790 1282.840 1213.110 ;
        RECT 1041.600 20.730 1041.740 1212.790 ;
        RECT 1037.400 20.410 1037.660 20.730 ;
        RECT 1041.540 20.410 1041.800 20.730 ;
        RECT 1037.460 2.400 1037.600 20.410 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1058.990 1213.360 1059.310 1213.420 ;
        RECT 1291.750 1213.360 1292.070 1213.420 ;
        RECT 1058.990 1213.220 1292.070 1213.360 ;
        RECT 1058.990 1213.160 1059.310 1213.220 ;
        RECT 1291.750 1213.160 1292.070 1213.220 ;
        RECT 1055.310 20.640 1055.630 20.700 ;
        RECT 1058.990 20.640 1059.310 20.700 ;
        RECT 1055.310 20.500 1059.310 20.640 ;
        RECT 1055.310 20.440 1055.630 20.500 ;
        RECT 1058.990 20.440 1059.310 20.500 ;
      LAYER via ;
        RECT 1059.020 1213.160 1059.280 1213.420 ;
        RECT 1291.780 1213.160 1292.040 1213.420 ;
        RECT 1055.340 20.440 1055.600 20.700 ;
        RECT 1059.020 20.440 1059.280 20.700 ;
      LAYER met2 ;
        RECT 1291.790 1219.680 1292.350 1228.680 ;
        RECT 1291.840 1213.450 1291.980 1219.680 ;
        RECT 1059.020 1213.130 1059.280 1213.450 ;
        RECT 1291.780 1213.130 1292.040 1213.450 ;
        RECT 1059.080 20.730 1059.220 1213.130 ;
        RECT 1055.340 20.410 1055.600 20.730 ;
        RECT 1059.020 20.410 1059.280 20.730 ;
        RECT 1055.400 2.400 1055.540 20.410 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1100.465 1210.485 1100.635 1214.055 ;
      LAYER mcon ;
        RECT 1100.465 1213.885 1100.635 1214.055 ;
      LAYER met1 ;
        RECT 1100.405 1214.040 1100.695 1214.085 ;
        RECT 1300.950 1214.040 1301.270 1214.100 ;
        RECT 1100.405 1213.900 1301.270 1214.040 ;
        RECT 1100.405 1213.855 1100.695 1213.900 ;
        RECT 1300.950 1213.840 1301.270 1213.900 ;
        RECT 1076.010 1210.640 1076.330 1210.700 ;
        RECT 1100.405 1210.640 1100.695 1210.685 ;
        RECT 1076.010 1210.500 1100.695 1210.640 ;
        RECT 1076.010 1210.440 1076.330 1210.500 ;
        RECT 1100.405 1210.455 1100.695 1210.500 ;
        RECT 1073.250 20.640 1073.570 20.700 ;
        RECT 1076.010 20.640 1076.330 20.700 ;
        RECT 1073.250 20.500 1076.330 20.640 ;
        RECT 1073.250 20.440 1073.570 20.500 ;
        RECT 1076.010 20.440 1076.330 20.500 ;
      LAYER via ;
        RECT 1300.980 1213.840 1301.240 1214.100 ;
        RECT 1076.040 1210.440 1076.300 1210.700 ;
        RECT 1073.280 20.440 1073.540 20.700 ;
        RECT 1076.040 20.440 1076.300 20.700 ;
      LAYER met2 ;
        RECT 1300.990 1219.680 1301.550 1228.680 ;
        RECT 1301.040 1214.130 1301.180 1219.680 ;
        RECT 1300.980 1213.810 1301.240 1214.130 ;
        RECT 1076.040 1210.410 1076.300 1210.730 ;
        RECT 1076.100 20.730 1076.240 1210.410 ;
        RECT 1073.280 20.410 1073.540 20.730 ;
        RECT 1076.040 20.410 1076.300 20.730 ;
        RECT 1073.340 2.400 1073.480 20.410 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1252.725 13.685 1252.895 16.235 ;
      LAYER mcon ;
        RECT 1252.725 16.065 1252.895 16.235 ;
      LAYER met1 ;
        RECT 1310.150 1213.020 1310.470 1213.080 ;
        RECT 1283.100 1212.880 1310.470 1213.020 ;
        RECT 1272.890 1212.680 1273.210 1212.740 ;
        RECT 1283.100 1212.680 1283.240 1212.880 ;
        RECT 1310.150 1212.820 1310.470 1212.880 ;
        RECT 1272.890 1212.540 1283.240 1212.680 ;
        RECT 1272.890 1212.480 1273.210 1212.540 ;
        RECT 1252.665 16.220 1252.955 16.265 ;
        RECT 1272.890 16.220 1273.210 16.280 ;
        RECT 1252.665 16.080 1273.210 16.220 ;
        RECT 1252.665 16.035 1252.955 16.080 ;
        RECT 1272.890 16.020 1273.210 16.080 ;
        RECT 1090.730 14.180 1091.050 14.240 ;
        RECT 1090.730 14.040 1245.060 14.180 ;
        RECT 1090.730 13.980 1091.050 14.040 ;
        RECT 1244.920 13.840 1245.060 14.040 ;
        RECT 1252.665 13.840 1252.955 13.885 ;
        RECT 1244.920 13.700 1252.955 13.840 ;
        RECT 1252.665 13.655 1252.955 13.700 ;
      LAYER via ;
        RECT 1272.920 1212.480 1273.180 1212.740 ;
        RECT 1310.180 1212.820 1310.440 1213.080 ;
        RECT 1272.920 16.020 1273.180 16.280 ;
        RECT 1090.760 13.980 1091.020 14.240 ;
      LAYER met2 ;
        RECT 1310.190 1219.680 1310.750 1228.680 ;
        RECT 1310.240 1213.110 1310.380 1219.680 ;
        RECT 1310.180 1212.790 1310.440 1213.110 ;
        RECT 1272.920 1212.450 1273.180 1212.770 ;
        RECT 1272.980 16.310 1273.120 1212.450 ;
        RECT 1272.920 15.990 1273.180 16.310 ;
        RECT 1090.760 13.950 1091.020 14.270 ;
        RECT 1090.820 2.400 1090.960 13.950 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1160.265 15.385 1160.435 16.915 ;
      LAYER mcon ;
        RECT 1160.265 16.745 1160.435 16.915 ;
      LAYER met1 ;
        RECT 1307.850 1209.620 1308.170 1209.680 ;
        RECT 1319.350 1209.620 1319.670 1209.680 ;
        RECT 1307.850 1209.480 1319.670 1209.620 ;
        RECT 1307.850 1209.420 1308.170 1209.480 ;
        RECT 1319.350 1209.420 1319.670 1209.480 ;
        RECT 1160.205 16.900 1160.495 16.945 ;
        RECT 1307.850 16.900 1308.170 16.960 ;
        RECT 1160.205 16.760 1292.900 16.900 ;
        RECT 1160.205 16.715 1160.495 16.760 ;
        RECT 1292.760 16.560 1292.900 16.760 ;
        RECT 1297.360 16.760 1308.170 16.900 ;
        RECT 1297.360 16.560 1297.500 16.760 ;
        RECT 1307.850 16.700 1308.170 16.760 ;
        RECT 1292.760 16.420 1297.500 16.560 ;
        RECT 1108.670 15.540 1108.990 15.600 ;
        RECT 1160.205 15.540 1160.495 15.585 ;
        RECT 1108.670 15.400 1160.495 15.540 ;
        RECT 1108.670 15.340 1108.990 15.400 ;
        RECT 1160.205 15.355 1160.495 15.400 ;
      LAYER via ;
        RECT 1307.880 1209.420 1308.140 1209.680 ;
        RECT 1319.380 1209.420 1319.640 1209.680 ;
        RECT 1307.880 16.700 1308.140 16.960 ;
        RECT 1108.700 15.340 1108.960 15.600 ;
      LAYER met2 ;
        RECT 1319.390 1219.680 1319.950 1228.680 ;
        RECT 1319.440 1209.710 1319.580 1219.680 ;
        RECT 1307.880 1209.390 1308.140 1209.710 ;
        RECT 1319.380 1209.390 1319.640 1209.710 ;
        RECT 1307.940 16.990 1308.080 1209.390 ;
        RECT 1307.880 16.670 1308.140 16.990 ;
        RECT 1108.700 15.310 1108.960 15.630 ;
        RECT 1108.760 2.400 1108.900 15.310 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 1210.640 1131.530 1210.700 ;
        RECT 1328.550 1210.640 1328.870 1210.700 ;
        RECT 1131.210 1210.500 1328.870 1210.640 ;
        RECT 1131.210 1210.440 1131.530 1210.500 ;
        RECT 1328.550 1210.440 1328.870 1210.500 ;
        RECT 1126.610 18.260 1126.930 18.320 ;
        RECT 1131.210 18.260 1131.530 18.320 ;
        RECT 1126.610 18.120 1131.530 18.260 ;
        RECT 1126.610 18.060 1126.930 18.120 ;
        RECT 1131.210 18.060 1131.530 18.120 ;
      LAYER via ;
        RECT 1131.240 1210.440 1131.500 1210.700 ;
        RECT 1328.580 1210.440 1328.840 1210.700 ;
        RECT 1126.640 18.060 1126.900 18.320 ;
        RECT 1131.240 18.060 1131.500 18.320 ;
      LAYER met2 ;
        RECT 1328.590 1219.680 1329.150 1228.680 ;
        RECT 1328.640 1210.730 1328.780 1219.680 ;
        RECT 1131.240 1210.410 1131.500 1210.730 ;
        RECT 1328.580 1210.410 1328.840 1210.730 ;
        RECT 1131.300 18.350 1131.440 1210.410 ;
        RECT 1126.640 18.030 1126.900 18.350 ;
        RECT 1131.240 18.030 1131.500 18.350 ;
        RECT 1126.700 2.400 1126.840 18.030 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1307.465 1209.465 1307.635 1214.055 ;
      LAYER mcon ;
        RECT 1307.465 1213.885 1307.635 1214.055 ;
      LAYER met1 ;
        RECT 1307.405 1214.040 1307.695 1214.085 ;
        RECT 1337.750 1214.040 1338.070 1214.100 ;
        RECT 1307.405 1213.900 1338.070 1214.040 ;
        RECT 1307.405 1213.855 1307.695 1213.900 ;
        RECT 1337.750 1213.840 1338.070 1213.900 ;
        RECT 1162.490 1209.620 1162.810 1209.680 ;
        RECT 1307.405 1209.620 1307.695 1209.665 ;
        RECT 1162.490 1209.480 1307.695 1209.620 ;
        RECT 1162.490 1209.420 1162.810 1209.480 ;
        RECT 1307.405 1209.435 1307.695 1209.480 ;
        RECT 1144.550 18.260 1144.870 18.320 ;
        RECT 1156.050 18.260 1156.370 18.320 ;
        RECT 1144.550 18.120 1156.370 18.260 ;
        RECT 1144.550 18.060 1144.870 18.120 ;
        RECT 1156.050 18.060 1156.370 18.120 ;
      LAYER via ;
        RECT 1337.780 1213.840 1338.040 1214.100 ;
        RECT 1162.520 1209.420 1162.780 1209.680 ;
        RECT 1144.580 18.060 1144.840 18.320 ;
        RECT 1156.080 18.060 1156.340 18.320 ;
      LAYER met2 ;
        RECT 1337.790 1219.680 1338.350 1228.680 ;
        RECT 1337.840 1214.130 1337.980 1219.680 ;
        RECT 1337.780 1213.810 1338.040 1214.130 ;
        RECT 1162.520 1209.390 1162.780 1209.710 ;
        RECT 1144.580 18.030 1144.840 18.350 ;
        RECT 1156.080 18.205 1156.340 18.350 ;
        RECT 1162.580 18.205 1162.720 1209.390 ;
        RECT 1144.640 2.400 1144.780 18.030 ;
        RECT 1156.070 17.835 1156.350 18.205 ;
        RECT 1162.510 17.835 1162.790 18.205 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 1156.070 17.880 1156.350 18.160 ;
        RECT 1162.510 17.880 1162.790 18.160 ;
      LAYER met3 ;
        RECT 1156.045 18.170 1156.375 18.185 ;
        RECT 1162.485 18.170 1162.815 18.185 ;
        RECT 1156.045 17.870 1162.815 18.170 ;
        RECT 1156.045 17.855 1156.375 17.870 ;
        RECT 1162.485 17.855 1162.815 17.870 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 14.520 1162.810 14.580 ;
        RECT 1346.030 14.520 1346.350 14.580 ;
        RECT 1162.490 14.380 1346.350 14.520 ;
        RECT 1162.490 14.320 1162.810 14.380 ;
        RECT 1346.030 14.320 1346.350 14.380 ;
      LAYER via ;
        RECT 1162.520 14.320 1162.780 14.580 ;
        RECT 1346.060 14.320 1346.320 14.580 ;
      LAYER met2 ;
        RECT 1346.990 1220.330 1347.550 1228.680 ;
        RECT 1346.580 1220.190 1347.550 1220.330 ;
        RECT 1346.580 21.490 1346.720 1220.190 ;
        RECT 1346.990 1219.680 1347.550 1220.190 ;
        RECT 1346.120 21.350 1346.720 21.490 ;
        RECT 1346.120 14.610 1346.260 21.350 ;
        RECT 1162.520 14.290 1162.780 14.610 ;
        RECT 1346.060 14.290 1346.320 14.610 ;
        RECT 1162.580 2.400 1162.720 14.290 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 680.410 29.820 680.730 29.880 ;
        RECT 1097.170 29.820 1097.490 29.880 ;
        RECT 680.410 29.680 1097.490 29.820 ;
        RECT 680.410 29.620 680.730 29.680 ;
        RECT 1097.170 29.620 1097.490 29.680 ;
      LAYER via ;
        RECT 680.440 29.620 680.700 29.880 ;
        RECT 1097.200 29.620 1097.460 29.880 ;
      LAYER met2 ;
        RECT 1099.510 1220.330 1100.070 1228.680 ;
        RECT 1097.260 1220.190 1100.070 1220.330 ;
        RECT 1097.260 29.910 1097.400 1220.190 ;
        RECT 1099.510 1219.680 1100.070 1220.190 ;
        RECT 680.440 29.590 680.700 29.910 ;
        RECT 1097.200 29.590 1097.460 29.910 ;
        RECT 680.500 2.400 680.640 29.590 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1217.690 1208.260 1218.010 1208.320 ;
        RECT 1356.150 1208.260 1356.470 1208.320 ;
        RECT 1217.690 1208.120 1356.470 1208.260 ;
        RECT 1217.690 1208.060 1218.010 1208.120 ;
        RECT 1356.150 1208.060 1356.470 1208.120 ;
        RECT 1179.970 18.260 1180.290 18.320 ;
        RECT 1217.690 18.260 1218.010 18.320 ;
        RECT 1179.970 18.120 1218.010 18.260 ;
        RECT 1179.970 18.060 1180.290 18.120 ;
        RECT 1217.690 18.060 1218.010 18.120 ;
      LAYER via ;
        RECT 1217.720 1208.060 1217.980 1208.320 ;
        RECT 1356.180 1208.060 1356.440 1208.320 ;
        RECT 1180.000 18.060 1180.260 18.320 ;
        RECT 1217.720 18.060 1217.980 18.320 ;
      LAYER met2 ;
        RECT 1356.190 1219.680 1356.750 1228.680 ;
        RECT 1356.240 1208.350 1356.380 1219.680 ;
        RECT 1217.720 1208.030 1217.980 1208.350 ;
        RECT 1356.180 1208.030 1356.440 1208.350 ;
        RECT 1217.780 18.350 1217.920 1208.030 ;
        RECT 1180.000 18.030 1180.260 18.350 ;
        RECT 1217.720 18.030 1217.980 18.350 ;
        RECT 1180.060 2.400 1180.200 18.030 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1360.365 1062.585 1360.535 1076.355 ;
        RECT 1360.365 469.285 1360.535 517.395 ;
        RECT 1360.365 379.525 1360.535 427.635 ;
        RECT 1359.445 241.485 1359.615 255.595 ;
      LAYER mcon ;
        RECT 1360.365 1076.185 1360.535 1076.355 ;
        RECT 1360.365 517.225 1360.535 517.395 ;
        RECT 1360.365 427.465 1360.535 427.635 ;
        RECT 1359.445 255.425 1359.615 255.595 ;
      LAYER met1 ;
        RECT 1360.290 1196.700 1360.610 1196.760 ;
        RECT 1363.970 1196.700 1364.290 1196.760 ;
        RECT 1360.290 1196.560 1364.290 1196.700 ;
        RECT 1360.290 1196.500 1360.610 1196.560 ;
        RECT 1363.970 1196.500 1364.290 1196.560 ;
        RECT 1360.290 1076.340 1360.610 1076.400 ;
        RECT 1360.095 1076.200 1360.610 1076.340 ;
        RECT 1360.290 1076.140 1360.610 1076.200 ;
        RECT 1360.290 1062.740 1360.610 1062.800 ;
        RECT 1360.095 1062.600 1360.610 1062.740 ;
        RECT 1360.290 1062.540 1360.610 1062.600 ;
        RECT 1359.370 966.180 1359.690 966.240 ;
        RECT 1360.290 966.180 1360.610 966.240 ;
        RECT 1359.370 966.040 1360.610 966.180 ;
        RECT 1359.370 965.980 1359.690 966.040 ;
        RECT 1360.290 965.980 1360.610 966.040 ;
        RECT 1359.370 869.620 1359.690 869.680 ;
        RECT 1360.290 869.620 1360.610 869.680 ;
        RECT 1359.370 869.480 1360.610 869.620 ;
        RECT 1359.370 869.420 1359.690 869.480 ;
        RECT 1360.290 869.420 1360.610 869.480 ;
        RECT 1359.370 772.720 1359.690 772.780 ;
        RECT 1360.290 772.720 1360.610 772.780 ;
        RECT 1359.370 772.580 1360.610 772.720 ;
        RECT 1359.370 772.520 1359.690 772.580 ;
        RECT 1360.290 772.520 1360.610 772.580 ;
        RECT 1359.370 676.160 1359.690 676.220 ;
        RECT 1360.290 676.160 1360.610 676.220 ;
        RECT 1359.370 676.020 1360.610 676.160 ;
        RECT 1359.370 675.960 1359.690 676.020 ;
        RECT 1360.290 675.960 1360.610 676.020 ;
        RECT 1359.830 572.460 1360.150 572.520 ;
        RECT 1360.290 572.460 1360.610 572.520 ;
        RECT 1359.830 572.320 1360.610 572.460 ;
        RECT 1359.830 572.260 1360.150 572.320 ;
        RECT 1360.290 572.260 1360.610 572.320 ;
        RECT 1360.290 517.380 1360.610 517.440 ;
        RECT 1360.095 517.240 1360.610 517.380 ;
        RECT 1360.290 517.180 1360.610 517.240 ;
        RECT 1360.290 469.440 1360.610 469.500 ;
        RECT 1360.095 469.300 1360.610 469.440 ;
        RECT 1360.290 469.240 1360.610 469.300 ;
        RECT 1360.290 427.620 1360.610 427.680 ;
        RECT 1360.095 427.480 1360.610 427.620 ;
        RECT 1360.290 427.420 1360.610 427.480 ;
        RECT 1360.290 379.680 1360.610 379.740 ;
        RECT 1360.095 379.540 1360.610 379.680 ;
        RECT 1360.290 379.480 1360.610 379.540 ;
        RECT 1359.385 255.580 1359.675 255.625 ;
        RECT 1360.290 255.580 1360.610 255.640 ;
        RECT 1359.385 255.440 1360.610 255.580 ;
        RECT 1359.385 255.395 1359.675 255.440 ;
        RECT 1360.290 255.380 1360.610 255.440 ;
        RECT 1359.370 241.640 1359.690 241.700 ;
        RECT 1359.175 241.500 1359.690 241.640 ;
        RECT 1359.370 241.440 1359.690 241.500 ;
        RECT 1359.830 144.740 1360.150 144.800 ;
        RECT 1360.290 144.740 1360.610 144.800 ;
        RECT 1359.830 144.600 1360.610 144.740 ;
        RECT 1359.830 144.540 1360.150 144.600 ;
        RECT 1360.290 144.540 1360.610 144.600 ;
        RECT 1197.910 17.580 1198.230 17.640 ;
        RECT 1359.830 17.580 1360.150 17.640 ;
        RECT 1197.910 17.440 1360.150 17.580 ;
        RECT 1197.910 17.380 1198.230 17.440 ;
        RECT 1359.830 17.380 1360.150 17.440 ;
      LAYER via ;
        RECT 1360.320 1196.500 1360.580 1196.760 ;
        RECT 1364.000 1196.500 1364.260 1196.760 ;
        RECT 1360.320 1076.140 1360.580 1076.400 ;
        RECT 1360.320 1062.540 1360.580 1062.800 ;
        RECT 1359.400 965.980 1359.660 966.240 ;
        RECT 1360.320 965.980 1360.580 966.240 ;
        RECT 1359.400 869.420 1359.660 869.680 ;
        RECT 1360.320 869.420 1360.580 869.680 ;
        RECT 1359.400 772.520 1359.660 772.780 ;
        RECT 1360.320 772.520 1360.580 772.780 ;
        RECT 1359.400 675.960 1359.660 676.220 ;
        RECT 1360.320 675.960 1360.580 676.220 ;
        RECT 1359.860 572.260 1360.120 572.520 ;
        RECT 1360.320 572.260 1360.580 572.520 ;
        RECT 1360.320 517.180 1360.580 517.440 ;
        RECT 1360.320 469.240 1360.580 469.500 ;
        RECT 1360.320 427.420 1360.580 427.680 ;
        RECT 1360.320 379.480 1360.580 379.740 ;
        RECT 1360.320 255.380 1360.580 255.640 ;
        RECT 1359.400 241.440 1359.660 241.700 ;
        RECT 1359.860 144.540 1360.120 144.800 ;
        RECT 1360.320 144.540 1360.580 144.800 ;
        RECT 1197.940 17.380 1198.200 17.640 ;
        RECT 1359.860 17.380 1360.120 17.640 ;
      LAYER met2 ;
        RECT 1364.930 1220.330 1365.490 1228.680 ;
        RECT 1364.060 1220.190 1365.490 1220.330 ;
        RECT 1364.060 1196.790 1364.200 1220.190 ;
        RECT 1364.930 1219.680 1365.490 1220.190 ;
        RECT 1360.320 1196.470 1360.580 1196.790 ;
        RECT 1364.000 1196.470 1364.260 1196.790 ;
        RECT 1360.380 1076.430 1360.520 1196.470 ;
        RECT 1360.320 1076.110 1360.580 1076.430 ;
        RECT 1360.320 1062.510 1360.580 1062.830 ;
        RECT 1360.380 1014.405 1360.520 1062.510 ;
        RECT 1359.390 1014.035 1359.670 1014.405 ;
        RECT 1360.310 1014.035 1360.590 1014.405 ;
        RECT 1359.460 966.270 1359.600 1014.035 ;
        RECT 1359.400 965.950 1359.660 966.270 ;
        RECT 1360.320 965.950 1360.580 966.270 ;
        RECT 1360.380 917.845 1360.520 965.950 ;
        RECT 1359.390 917.475 1359.670 917.845 ;
        RECT 1360.310 917.475 1360.590 917.845 ;
        RECT 1359.460 869.710 1359.600 917.475 ;
        RECT 1359.400 869.390 1359.660 869.710 ;
        RECT 1360.320 869.390 1360.580 869.710 ;
        RECT 1360.380 787.170 1360.520 869.390 ;
        RECT 1359.920 787.030 1360.520 787.170 ;
        RECT 1359.920 786.490 1360.060 787.030 ;
        RECT 1359.920 786.350 1360.520 786.490 ;
        RECT 1360.380 772.810 1360.520 786.350 ;
        RECT 1359.400 772.490 1359.660 772.810 ;
        RECT 1360.320 772.490 1360.580 772.810 ;
        RECT 1359.460 724.725 1359.600 772.490 ;
        RECT 1359.390 724.355 1359.670 724.725 ;
        RECT 1360.310 724.355 1360.590 724.725 ;
        RECT 1360.380 676.250 1360.520 724.355 ;
        RECT 1359.400 675.930 1359.660 676.250 ;
        RECT 1360.320 675.930 1360.580 676.250 ;
        RECT 1359.460 628.165 1359.600 675.930 ;
        RECT 1359.390 627.795 1359.670 628.165 ;
        RECT 1360.310 627.795 1360.590 628.165 ;
        RECT 1360.380 580.450 1360.520 627.795 ;
        RECT 1359.920 580.310 1360.520 580.450 ;
        RECT 1359.920 579.770 1360.060 580.310 ;
        RECT 1359.920 579.630 1360.520 579.770 ;
        RECT 1360.380 572.550 1360.520 579.630 ;
        RECT 1359.860 572.230 1360.120 572.550 ;
        RECT 1360.320 572.230 1360.580 572.550 ;
        RECT 1359.920 524.690 1360.060 572.230 ;
        RECT 1359.920 524.550 1360.520 524.690 ;
        RECT 1360.380 517.470 1360.520 524.550 ;
        RECT 1360.320 517.150 1360.580 517.470 ;
        RECT 1360.320 469.210 1360.580 469.530 ;
        RECT 1360.380 427.710 1360.520 469.210 ;
        RECT 1360.320 427.390 1360.580 427.710 ;
        RECT 1360.320 379.450 1360.580 379.770 ;
        RECT 1360.380 255.670 1360.520 379.450 ;
        RECT 1360.320 255.350 1360.580 255.670 ;
        RECT 1359.400 241.410 1359.660 241.730 ;
        RECT 1359.460 206.450 1359.600 241.410 ;
        RECT 1359.460 206.310 1360.520 206.450 ;
        RECT 1360.380 144.830 1360.520 206.310 ;
        RECT 1359.860 144.510 1360.120 144.830 ;
        RECT 1360.320 144.510 1360.580 144.830 ;
        RECT 1359.920 17.670 1360.060 144.510 ;
        RECT 1197.940 17.350 1198.200 17.670 ;
        RECT 1359.860 17.350 1360.120 17.670 ;
        RECT 1198.000 2.400 1198.140 17.350 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1359.390 1014.080 1359.670 1014.360 ;
        RECT 1360.310 1014.080 1360.590 1014.360 ;
        RECT 1359.390 917.520 1359.670 917.800 ;
        RECT 1360.310 917.520 1360.590 917.800 ;
        RECT 1359.390 724.400 1359.670 724.680 ;
        RECT 1360.310 724.400 1360.590 724.680 ;
        RECT 1359.390 627.840 1359.670 628.120 ;
        RECT 1360.310 627.840 1360.590 628.120 ;
      LAYER met3 ;
        RECT 1359.365 1014.370 1359.695 1014.385 ;
        RECT 1360.285 1014.370 1360.615 1014.385 ;
        RECT 1359.365 1014.070 1360.615 1014.370 ;
        RECT 1359.365 1014.055 1359.695 1014.070 ;
        RECT 1360.285 1014.055 1360.615 1014.070 ;
        RECT 1359.365 917.810 1359.695 917.825 ;
        RECT 1360.285 917.810 1360.615 917.825 ;
        RECT 1359.365 917.510 1360.615 917.810 ;
        RECT 1359.365 917.495 1359.695 917.510 ;
        RECT 1360.285 917.495 1360.615 917.510 ;
        RECT 1359.365 724.690 1359.695 724.705 ;
        RECT 1360.285 724.690 1360.615 724.705 ;
        RECT 1359.365 724.390 1360.615 724.690 ;
        RECT 1359.365 724.375 1359.695 724.390 ;
        RECT 1360.285 724.375 1360.615 724.390 ;
        RECT 1359.365 628.130 1359.695 628.145 ;
        RECT 1360.285 628.130 1360.615 628.145 ;
        RECT 1359.365 627.830 1360.615 628.130 ;
        RECT 1359.365 627.815 1359.695 627.830 ;
        RECT 1360.285 627.815 1360.615 627.830 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1341.965 1207.425 1342.135 1210.315 ;
      LAYER mcon ;
        RECT 1341.965 1210.145 1342.135 1210.315 ;
      LAYER met1 ;
        RECT 1220.910 1210.300 1221.230 1210.360 ;
        RECT 1341.905 1210.300 1342.195 1210.345 ;
        RECT 1220.910 1210.160 1342.195 1210.300 ;
        RECT 1220.910 1210.100 1221.230 1210.160 ;
        RECT 1341.905 1210.115 1342.195 1210.160 ;
        RECT 1341.905 1207.580 1342.195 1207.625 ;
        RECT 1374.090 1207.580 1374.410 1207.640 ;
        RECT 1341.905 1207.440 1374.410 1207.580 ;
        RECT 1341.905 1207.395 1342.195 1207.440 ;
        RECT 1374.090 1207.380 1374.410 1207.440 ;
        RECT 1215.850 18.940 1216.170 19.000 ;
        RECT 1220.910 18.940 1221.230 19.000 ;
        RECT 1215.850 18.800 1221.230 18.940 ;
        RECT 1215.850 18.740 1216.170 18.800 ;
        RECT 1220.910 18.740 1221.230 18.800 ;
      LAYER via ;
        RECT 1220.940 1210.100 1221.200 1210.360 ;
        RECT 1374.120 1207.380 1374.380 1207.640 ;
        RECT 1215.880 18.740 1216.140 19.000 ;
        RECT 1220.940 18.740 1221.200 19.000 ;
      LAYER met2 ;
        RECT 1374.130 1219.680 1374.690 1228.680 ;
        RECT 1220.940 1210.070 1221.200 1210.390 ;
        RECT 1221.000 19.030 1221.140 1210.070 ;
        RECT 1374.180 1207.670 1374.320 1219.680 ;
        RECT 1374.120 1207.350 1374.380 1207.670 ;
        RECT 1215.880 18.710 1216.140 19.030 ;
        RECT 1220.940 18.710 1221.200 19.030 ;
        RECT 1215.940 2.400 1216.080 18.710 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1341.965 18.105 1342.135 20.315 ;
      LAYER mcon ;
        RECT 1341.965 20.145 1342.135 20.315 ;
      LAYER met1 ;
        RECT 1380.070 1196.700 1380.390 1196.760 ;
        RECT 1382.370 1196.700 1382.690 1196.760 ;
        RECT 1380.070 1196.560 1382.690 1196.700 ;
        RECT 1380.070 1196.500 1380.390 1196.560 ;
        RECT 1382.370 1196.500 1382.690 1196.560 ;
        RECT 1341.905 20.300 1342.195 20.345 ;
        RECT 1380.070 20.300 1380.390 20.360 ;
        RECT 1341.905 20.160 1380.390 20.300 ;
        RECT 1341.905 20.115 1342.195 20.160 ;
        RECT 1380.070 20.100 1380.390 20.160 ;
        RECT 1233.790 18.260 1234.110 18.320 ;
        RECT 1341.905 18.260 1342.195 18.305 ;
        RECT 1233.790 18.120 1342.195 18.260 ;
        RECT 1233.790 18.060 1234.110 18.120 ;
        RECT 1341.905 18.075 1342.195 18.120 ;
      LAYER via ;
        RECT 1380.100 1196.500 1380.360 1196.760 ;
        RECT 1382.400 1196.500 1382.660 1196.760 ;
        RECT 1380.100 20.100 1380.360 20.360 ;
        RECT 1233.820 18.060 1234.080 18.320 ;
      LAYER met2 ;
        RECT 1383.330 1220.330 1383.890 1228.680 ;
        RECT 1382.460 1220.190 1383.890 1220.330 ;
        RECT 1382.460 1196.790 1382.600 1220.190 ;
        RECT 1383.330 1219.680 1383.890 1220.190 ;
        RECT 1380.100 1196.470 1380.360 1196.790 ;
        RECT 1382.400 1196.470 1382.660 1196.790 ;
        RECT 1380.160 1172.730 1380.300 1196.470 ;
        RECT 1380.160 1172.590 1380.760 1172.730 ;
        RECT 1380.620 1028.570 1380.760 1172.590 ;
        RECT 1380.160 1028.430 1380.760 1028.570 ;
        RECT 1380.160 1027.890 1380.300 1028.430 ;
        RECT 1380.160 1027.750 1380.760 1027.890 ;
        RECT 1380.620 932.010 1380.760 1027.750 ;
        RECT 1380.160 931.870 1380.760 932.010 ;
        RECT 1380.160 931.330 1380.300 931.870 ;
        RECT 1380.160 931.190 1380.760 931.330 ;
        RECT 1380.620 835.450 1380.760 931.190 ;
        RECT 1380.160 835.310 1380.760 835.450 ;
        RECT 1380.160 834.770 1380.300 835.310 ;
        RECT 1380.160 834.630 1380.760 834.770 ;
        RECT 1380.620 738.890 1380.760 834.630 ;
        RECT 1380.160 738.750 1380.760 738.890 ;
        RECT 1380.160 738.210 1380.300 738.750 ;
        RECT 1380.160 738.070 1380.760 738.210 ;
        RECT 1380.620 642.330 1380.760 738.070 ;
        RECT 1380.160 642.190 1380.760 642.330 ;
        RECT 1380.160 641.650 1380.300 642.190 ;
        RECT 1380.160 641.510 1380.760 641.650 ;
        RECT 1380.620 545.770 1380.760 641.510 ;
        RECT 1380.160 545.630 1380.760 545.770 ;
        RECT 1380.160 545.090 1380.300 545.630 ;
        RECT 1380.160 544.950 1380.760 545.090 ;
        RECT 1380.620 449.210 1380.760 544.950 ;
        RECT 1380.160 449.070 1380.760 449.210 ;
        RECT 1380.160 448.530 1380.300 449.070 ;
        RECT 1380.160 448.390 1380.760 448.530 ;
        RECT 1380.620 351.970 1380.760 448.390 ;
        RECT 1380.160 351.830 1380.760 351.970 ;
        RECT 1380.160 351.290 1380.300 351.830 ;
        RECT 1380.160 351.150 1380.760 351.290 ;
        RECT 1380.620 255.410 1380.760 351.150 ;
        RECT 1380.160 255.270 1380.760 255.410 ;
        RECT 1380.160 254.730 1380.300 255.270 ;
        RECT 1380.160 254.590 1380.760 254.730 ;
        RECT 1380.620 158.850 1380.760 254.590 ;
        RECT 1380.160 158.710 1380.760 158.850 ;
        RECT 1380.160 158.170 1380.300 158.710 ;
        RECT 1380.160 158.030 1380.760 158.170 ;
        RECT 1380.620 72.490 1380.760 158.030 ;
        RECT 1380.160 72.350 1380.760 72.490 ;
        RECT 1380.160 20.390 1380.300 72.350 ;
        RECT 1380.100 20.070 1380.360 20.390 ;
        RECT 1233.820 18.030 1234.080 18.350 ;
        RECT 1233.880 2.400 1234.020 18.030 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1371.865 1207.765 1372.035 1209.295 ;
      LAYER mcon ;
        RECT 1371.865 1209.125 1372.035 1209.295 ;
      LAYER met1 ;
        RECT 1371.805 1209.280 1372.095 1209.325 ;
        RECT 1392.490 1209.280 1392.810 1209.340 ;
        RECT 1371.805 1209.140 1392.810 1209.280 ;
        RECT 1371.805 1209.095 1372.095 1209.140 ;
        RECT 1392.490 1209.080 1392.810 1209.140 ;
        RECT 1255.410 1207.920 1255.730 1207.980 ;
        RECT 1371.805 1207.920 1372.095 1207.965 ;
        RECT 1255.410 1207.780 1372.095 1207.920 ;
        RECT 1255.410 1207.720 1255.730 1207.780 ;
        RECT 1371.805 1207.735 1372.095 1207.780 ;
        RECT 1251.730 18.940 1252.050 19.000 ;
        RECT 1255.410 18.940 1255.730 19.000 ;
        RECT 1251.730 18.800 1255.730 18.940 ;
        RECT 1251.730 18.740 1252.050 18.800 ;
        RECT 1255.410 18.740 1255.730 18.800 ;
      LAYER via ;
        RECT 1392.520 1209.080 1392.780 1209.340 ;
        RECT 1255.440 1207.720 1255.700 1207.980 ;
        RECT 1251.760 18.740 1252.020 19.000 ;
        RECT 1255.440 18.740 1255.700 19.000 ;
      LAYER met2 ;
        RECT 1392.530 1219.680 1393.090 1228.680 ;
        RECT 1392.580 1209.370 1392.720 1219.680 ;
        RECT 1392.520 1209.050 1392.780 1209.370 ;
        RECT 1255.440 1207.690 1255.700 1208.010 ;
        RECT 1255.500 19.030 1255.640 1207.690 ;
        RECT 1251.760 18.710 1252.020 19.030 ;
        RECT 1255.440 18.710 1255.700 19.030 ;
        RECT 1251.820 2.400 1251.960 18.710 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1383.825 1211.165 1383.995 1213.715 ;
      LAYER mcon ;
        RECT 1383.825 1213.545 1383.995 1213.715 ;
      LAYER met1 ;
        RECT 1383.765 1213.700 1384.055 1213.745 ;
        RECT 1401.690 1213.700 1402.010 1213.760 ;
        RECT 1383.765 1213.560 1402.010 1213.700 ;
        RECT 1383.765 1213.515 1384.055 1213.560 ;
        RECT 1401.690 1213.500 1402.010 1213.560 ;
        RECT 1273.350 1211.320 1273.670 1211.380 ;
        RECT 1383.765 1211.320 1384.055 1211.365 ;
        RECT 1273.350 1211.180 1384.055 1211.320 ;
        RECT 1273.350 1211.120 1273.670 1211.180 ;
        RECT 1383.765 1211.135 1384.055 1211.180 ;
        RECT 1269.210 16.560 1269.530 16.620 ;
        RECT 1273.350 16.560 1273.670 16.620 ;
        RECT 1269.210 16.420 1273.670 16.560 ;
        RECT 1269.210 16.360 1269.530 16.420 ;
        RECT 1273.350 16.360 1273.670 16.420 ;
      LAYER via ;
        RECT 1401.720 1213.500 1401.980 1213.760 ;
        RECT 1273.380 1211.120 1273.640 1211.380 ;
        RECT 1269.240 16.360 1269.500 16.620 ;
        RECT 1273.380 16.360 1273.640 16.620 ;
      LAYER met2 ;
        RECT 1401.730 1219.680 1402.290 1228.680 ;
        RECT 1401.780 1213.790 1401.920 1219.680 ;
        RECT 1401.720 1213.470 1401.980 1213.790 ;
        RECT 1273.380 1211.090 1273.640 1211.410 ;
        RECT 1273.440 16.650 1273.580 1211.090 ;
        RECT 1269.240 16.330 1269.500 16.650 ;
        RECT 1273.380 16.330 1273.640 16.650 ;
        RECT 1269.300 2.400 1269.440 16.330 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 1214.380 1290.230 1214.440 ;
        RECT 1289.910 1214.240 1366.500 1214.380 ;
        RECT 1289.910 1214.180 1290.230 1214.240 ;
        RECT 1366.360 1214.040 1366.500 1214.240 ;
        RECT 1410.890 1214.040 1411.210 1214.100 ;
        RECT 1366.360 1213.900 1411.210 1214.040 ;
        RECT 1410.890 1213.840 1411.210 1213.900 ;
        RECT 1287.150 16.560 1287.470 16.620 ;
        RECT 1289.910 16.560 1290.230 16.620 ;
        RECT 1287.150 16.420 1290.230 16.560 ;
        RECT 1287.150 16.360 1287.470 16.420 ;
        RECT 1289.910 16.360 1290.230 16.420 ;
      LAYER via ;
        RECT 1289.940 1214.180 1290.200 1214.440 ;
        RECT 1410.920 1213.840 1411.180 1214.100 ;
        RECT 1287.180 16.360 1287.440 16.620 ;
        RECT 1289.940 16.360 1290.200 16.620 ;
      LAYER met2 ;
        RECT 1410.930 1219.680 1411.490 1228.680 ;
        RECT 1289.940 1214.150 1290.200 1214.470 ;
        RECT 1290.000 16.650 1290.140 1214.150 ;
        RECT 1410.980 1214.130 1411.120 1219.680 ;
        RECT 1410.920 1213.810 1411.180 1214.130 ;
        RECT 1287.180 16.330 1287.440 16.650 ;
        RECT 1289.940 16.330 1290.200 16.650 ;
        RECT 1287.240 2.400 1287.380 16.330 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.030 19.280 1415.350 19.340 ;
        RECT 1306.100 19.140 1415.350 19.280 ;
        RECT 1305.090 18.940 1305.410 19.000 ;
        RECT 1306.100 18.940 1306.240 19.140 ;
        RECT 1415.030 19.080 1415.350 19.140 ;
        RECT 1305.090 18.800 1306.240 18.940 ;
        RECT 1305.090 18.740 1305.410 18.800 ;
      LAYER via ;
        RECT 1305.120 18.740 1305.380 19.000 ;
        RECT 1415.060 19.080 1415.320 19.340 ;
      LAYER met2 ;
        RECT 1420.130 1221.010 1420.690 1228.680 ;
        RECT 1417.880 1220.870 1420.690 1221.010 ;
        RECT 1417.880 1206.730 1418.020 1220.870 ;
        RECT 1420.130 1219.680 1420.690 1220.870 ;
        RECT 1415.120 1206.590 1418.020 1206.730 ;
        RECT 1415.120 19.370 1415.260 1206.590 ;
        RECT 1415.060 19.050 1415.320 19.370 ;
        RECT 1305.120 18.710 1305.380 19.030 ;
        RECT 1305.180 2.400 1305.320 18.710 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1323.030 19.960 1323.350 20.020 ;
        RECT 1428.830 19.960 1429.150 20.020 ;
        RECT 1323.030 19.820 1429.150 19.960 ;
        RECT 1323.030 19.760 1323.350 19.820 ;
        RECT 1428.830 19.760 1429.150 19.820 ;
      LAYER via ;
        RECT 1323.060 19.760 1323.320 20.020 ;
        RECT 1428.860 19.760 1429.120 20.020 ;
      LAYER met2 ;
        RECT 1429.330 1220.330 1429.890 1228.680 ;
        RECT 1428.920 1220.190 1429.890 1220.330 ;
        RECT 1428.920 20.050 1429.060 1220.190 ;
        RECT 1429.330 1219.680 1429.890 1220.190 ;
        RECT 1323.060 19.730 1323.320 20.050 ;
        RECT 1428.860 19.730 1429.120 20.050 ;
        RECT 1323.120 2.400 1323.260 19.730 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 1209.960 1345.430 1210.020 ;
        RECT 1438.490 1209.960 1438.810 1210.020 ;
        RECT 1345.110 1209.820 1438.810 1209.960 ;
        RECT 1345.110 1209.760 1345.430 1209.820 ;
        RECT 1438.490 1209.760 1438.810 1209.820 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1345.110 20.640 1345.430 20.700 ;
        RECT 1340.510 20.500 1345.430 20.640 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
        RECT 1345.110 20.440 1345.430 20.500 ;
      LAYER via ;
        RECT 1345.140 1209.760 1345.400 1210.020 ;
        RECT 1438.520 1209.760 1438.780 1210.020 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
        RECT 1345.140 20.440 1345.400 20.700 ;
      LAYER met2 ;
        RECT 1438.530 1219.680 1439.090 1228.680 ;
        RECT 1438.580 1210.050 1438.720 1219.680 ;
        RECT 1345.140 1209.730 1345.400 1210.050 ;
        RECT 1438.520 1209.730 1438.780 1210.050 ;
        RECT 1345.200 20.730 1345.340 1209.730 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1345.140 20.410 1345.400 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1104.070 1196.700 1104.390 1196.760 ;
        RECT 1106.830 1196.700 1107.150 1196.760 ;
        RECT 1104.070 1196.560 1107.150 1196.700 ;
        RECT 1104.070 1196.500 1104.390 1196.560 ;
        RECT 1106.830 1196.500 1107.150 1196.560 ;
        RECT 698.350 29.480 698.670 29.540 ;
        RECT 1104.070 29.480 1104.390 29.540 ;
        RECT 698.350 29.340 1104.390 29.480 ;
        RECT 698.350 29.280 698.670 29.340 ;
        RECT 1104.070 29.280 1104.390 29.340 ;
      LAYER via ;
        RECT 1104.100 1196.500 1104.360 1196.760 ;
        RECT 1106.860 1196.500 1107.120 1196.760 ;
        RECT 698.380 29.280 698.640 29.540 ;
        RECT 1104.100 29.280 1104.360 29.540 ;
      LAYER met2 ;
        RECT 1108.710 1220.330 1109.270 1228.680 ;
        RECT 1106.920 1220.190 1109.270 1220.330 ;
        RECT 1106.920 1196.790 1107.060 1220.190 ;
        RECT 1108.710 1219.680 1109.270 1220.190 ;
        RECT 1104.100 1196.470 1104.360 1196.790 ;
        RECT 1106.860 1196.470 1107.120 1196.790 ;
        RECT 1104.160 29.570 1104.300 1196.470 ;
        RECT 698.380 29.250 698.640 29.570 ;
        RECT 1104.100 29.250 1104.360 29.570 ;
        RECT 698.440 2.400 698.580 29.250 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.910 1209.620 1359.230 1209.680 ;
        RECT 1447.690 1209.620 1448.010 1209.680 ;
        RECT 1358.910 1209.480 1448.010 1209.620 ;
        RECT 1358.910 1209.420 1359.230 1209.480 ;
        RECT 1447.690 1209.420 1448.010 1209.480 ;
      LAYER via ;
        RECT 1358.940 1209.420 1359.200 1209.680 ;
        RECT 1447.720 1209.420 1447.980 1209.680 ;
      LAYER met2 ;
        RECT 1447.730 1219.680 1448.290 1228.680 ;
        RECT 1447.780 1209.710 1447.920 1219.680 ;
        RECT 1358.940 1209.390 1359.200 1209.710 ;
        RECT 1447.720 1209.390 1447.980 1209.710 ;
        RECT 1359.000 3.130 1359.140 1209.390 ;
        RECT 1358.540 2.990 1359.140 3.130 ;
        RECT 1358.540 2.400 1358.680 2.990 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.610 1210.300 1379.930 1210.360 ;
        RECT 1456.890 1210.300 1457.210 1210.360 ;
        RECT 1379.610 1210.160 1457.210 1210.300 ;
        RECT 1379.610 1210.100 1379.930 1210.160 ;
        RECT 1456.890 1210.100 1457.210 1210.160 ;
        RECT 1376.390 15.200 1376.710 15.260 ;
        RECT 1379.610 15.200 1379.930 15.260 ;
        RECT 1376.390 15.060 1379.930 15.200 ;
        RECT 1376.390 15.000 1376.710 15.060 ;
        RECT 1379.610 15.000 1379.930 15.060 ;
      LAYER via ;
        RECT 1379.640 1210.100 1379.900 1210.360 ;
        RECT 1456.920 1210.100 1457.180 1210.360 ;
        RECT 1376.420 15.000 1376.680 15.260 ;
        RECT 1379.640 15.000 1379.900 15.260 ;
      LAYER met2 ;
        RECT 1456.930 1219.680 1457.490 1228.680 ;
        RECT 1456.980 1210.390 1457.120 1219.680 ;
        RECT 1379.640 1210.070 1379.900 1210.390 ;
        RECT 1456.920 1210.070 1457.180 1210.390 ;
        RECT 1379.700 15.290 1379.840 1210.070 ;
        RECT 1376.420 14.970 1376.680 15.290 ;
        RECT 1379.640 14.970 1379.900 15.290 ;
        RECT 1376.480 2.400 1376.620 14.970 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1459.190 1207.580 1459.510 1207.640 ;
        RECT 1466.090 1207.580 1466.410 1207.640 ;
        RECT 1459.190 1207.440 1466.410 1207.580 ;
        RECT 1459.190 1207.380 1459.510 1207.440 ;
        RECT 1466.090 1207.380 1466.410 1207.440 ;
        RECT 1394.330 17.240 1394.650 17.300 ;
        RECT 1394.330 17.100 1436.880 17.240 ;
        RECT 1394.330 17.040 1394.650 17.100 ;
        RECT 1436.740 16.900 1436.880 17.100 ;
        RECT 1459.190 16.900 1459.510 16.960 ;
        RECT 1436.740 16.760 1459.510 16.900 ;
        RECT 1459.190 16.700 1459.510 16.760 ;
      LAYER via ;
        RECT 1459.220 1207.380 1459.480 1207.640 ;
        RECT 1466.120 1207.380 1466.380 1207.640 ;
        RECT 1394.360 17.040 1394.620 17.300 ;
        RECT 1459.220 16.700 1459.480 16.960 ;
      LAYER met2 ;
        RECT 1466.130 1219.680 1466.690 1228.680 ;
        RECT 1466.180 1207.670 1466.320 1219.680 ;
        RECT 1459.220 1207.350 1459.480 1207.670 ;
        RECT 1466.120 1207.350 1466.380 1207.670 ;
        RECT 1394.360 17.010 1394.620 17.330 ;
        RECT 1394.420 2.400 1394.560 17.010 ;
        RECT 1459.280 16.990 1459.420 1207.350 ;
        RECT 1459.220 16.670 1459.480 16.990 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1412.270 18.260 1412.590 18.320 ;
        RECT 1470.690 18.260 1471.010 18.320 ;
        RECT 1412.270 18.120 1471.010 18.260 ;
        RECT 1412.270 18.060 1412.590 18.120 ;
        RECT 1470.690 18.060 1471.010 18.120 ;
      LAYER via ;
        RECT 1412.300 18.060 1412.560 18.320 ;
        RECT 1470.720 18.060 1470.980 18.320 ;
      LAYER met2 ;
        RECT 1475.330 1220.330 1475.890 1228.680 ;
        RECT 1473.080 1220.190 1475.890 1220.330 ;
        RECT 1473.080 1206.730 1473.220 1220.190 ;
        RECT 1475.330 1219.680 1475.890 1220.190 ;
        RECT 1470.780 1206.590 1473.220 1206.730 ;
        RECT 1470.780 18.350 1470.920 1206.590 ;
        RECT 1412.300 18.030 1412.560 18.350 ;
        RECT 1470.720 18.030 1470.980 18.350 ;
        RECT 1412.360 2.400 1412.500 18.030 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1473.910 1213.700 1474.230 1213.760 ;
        RECT 1484.030 1213.700 1484.350 1213.760 ;
        RECT 1473.910 1213.560 1484.350 1213.700 ;
        RECT 1473.910 1213.500 1474.230 1213.560 ;
        RECT 1484.030 1213.500 1484.350 1213.560 ;
        RECT 1429.750 18.600 1430.070 18.660 ;
        RECT 1472.990 18.600 1473.310 18.660 ;
        RECT 1429.750 18.460 1473.310 18.600 ;
        RECT 1429.750 18.400 1430.070 18.460 ;
        RECT 1472.990 18.400 1473.310 18.460 ;
      LAYER via ;
        RECT 1473.940 1213.500 1474.200 1213.760 ;
        RECT 1484.060 1213.500 1484.320 1213.760 ;
        RECT 1429.780 18.400 1430.040 18.660 ;
        RECT 1473.020 18.400 1473.280 18.660 ;
      LAYER met2 ;
        RECT 1484.070 1219.680 1484.630 1228.680 ;
        RECT 1484.120 1213.790 1484.260 1219.680 ;
        RECT 1473.940 1213.470 1474.200 1213.790 ;
        RECT 1484.060 1213.470 1484.320 1213.790 ;
        RECT 1474.000 1193.810 1474.140 1213.470 ;
        RECT 1473.080 1193.670 1474.140 1193.810 ;
        RECT 1473.080 18.690 1473.220 1193.670 ;
        RECT 1429.780 18.370 1430.040 18.690 ;
        RECT 1473.020 18.370 1473.280 18.690 ;
        RECT 1429.840 2.400 1429.980 18.370 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1486.790 1207.580 1487.110 1207.640 ;
        RECT 1493.230 1207.580 1493.550 1207.640 ;
        RECT 1486.790 1207.440 1493.550 1207.580 ;
        RECT 1486.790 1207.380 1487.110 1207.440 ;
        RECT 1493.230 1207.380 1493.550 1207.440 ;
        RECT 1447.690 17.240 1448.010 17.300 ;
        RECT 1486.790 17.240 1487.110 17.300 ;
        RECT 1447.690 17.100 1487.110 17.240 ;
        RECT 1447.690 17.040 1448.010 17.100 ;
        RECT 1486.790 17.040 1487.110 17.100 ;
      LAYER via ;
        RECT 1486.820 1207.380 1487.080 1207.640 ;
        RECT 1493.260 1207.380 1493.520 1207.640 ;
        RECT 1447.720 17.040 1447.980 17.300 ;
        RECT 1486.820 17.040 1487.080 17.300 ;
      LAYER met2 ;
        RECT 1493.270 1219.680 1493.830 1228.680 ;
        RECT 1493.320 1207.670 1493.460 1219.680 ;
        RECT 1486.820 1207.350 1487.080 1207.670 ;
        RECT 1493.260 1207.350 1493.520 1207.670 ;
        RECT 1486.880 17.330 1487.020 1207.350 ;
        RECT 1447.720 17.010 1447.980 17.330 ;
        RECT 1486.820 17.010 1487.080 17.330 ;
        RECT 1447.780 2.400 1447.920 17.010 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1494.150 1207.580 1494.470 1207.640 ;
        RECT 1502.430 1207.580 1502.750 1207.640 ;
        RECT 1494.150 1207.440 1502.750 1207.580 ;
        RECT 1494.150 1207.380 1494.470 1207.440 ;
        RECT 1502.430 1207.380 1502.750 1207.440 ;
        RECT 1465.630 15.200 1465.950 15.260 ;
        RECT 1494.150 15.200 1494.470 15.260 ;
        RECT 1465.630 15.060 1494.470 15.200 ;
        RECT 1465.630 15.000 1465.950 15.060 ;
        RECT 1494.150 15.000 1494.470 15.060 ;
      LAYER via ;
        RECT 1494.180 1207.380 1494.440 1207.640 ;
        RECT 1502.460 1207.380 1502.720 1207.640 ;
        RECT 1465.660 15.000 1465.920 15.260 ;
        RECT 1494.180 15.000 1494.440 15.260 ;
      LAYER met2 ;
        RECT 1502.470 1219.680 1503.030 1228.680 ;
        RECT 1502.520 1207.670 1502.660 1219.680 ;
        RECT 1494.180 1207.350 1494.440 1207.670 ;
        RECT 1502.460 1207.350 1502.720 1207.670 ;
        RECT 1494.240 15.290 1494.380 1207.350 ;
        RECT 1465.660 14.970 1465.920 15.290 ;
        RECT 1494.180 14.970 1494.440 15.290 ;
        RECT 1465.720 2.400 1465.860 14.970 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.570 14.520 1483.890 14.580 ;
        RECT 1512.090 14.520 1512.410 14.580 ;
        RECT 1483.570 14.380 1512.410 14.520 ;
        RECT 1483.570 14.320 1483.890 14.380 ;
        RECT 1512.090 14.320 1512.410 14.380 ;
      LAYER via ;
        RECT 1483.600 14.320 1483.860 14.580 ;
        RECT 1512.120 14.320 1512.380 14.580 ;
      LAYER met2 ;
        RECT 1511.670 1220.330 1512.230 1228.680 ;
        RECT 1511.670 1219.680 1512.320 1220.330 ;
        RECT 1512.180 14.610 1512.320 1219.680 ;
        RECT 1483.600 14.290 1483.860 14.610 ;
        RECT 1512.120 14.290 1512.380 14.610 ;
        RECT 1483.660 2.400 1483.800 14.290 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1519.065 1159.145 1519.235 1207.255 ;
        RECT 1519.525 350.965 1519.695 386.155 ;
      LAYER mcon ;
        RECT 1519.065 1207.085 1519.235 1207.255 ;
        RECT 1519.525 385.985 1519.695 386.155 ;
      LAYER met1 ;
        RECT 1518.990 1207.240 1519.310 1207.300 ;
        RECT 1518.795 1207.100 1519.310 1207.240 ;
        RECT 1518.990 1207.040 1519.310 1207.100 ;
        RECT 1519.005 1159.300 1519.295 1159.345 ;
        RECT 1519.450 1159.300 1519.770 1159.360 ;
        RECT 1519.005 1159.160 1519.770 1159.300 ;
        RECT 1519.005 1159.115 1519.295 1159.160 ;
        RECT 1519.450 1159.100 1519.770 1159.160 ;
        RECT 1519.450 724.440 1519.770 724.500 ;
        RECT 1519.910 724.440 1520.230 724.500 ;
        RECT 1519.450 724.300 1520.230 724.440 ;
        RECT 1519.450 724.240 1519.770 724.300 ;
        RECT 1519.910 724.240 1520.230 724.300 ;
        RECT 1519.450 627.880 1519.770 627.940 ;
        RECT 1519.910 627.880 1520.230 627.940 ;
        RECT 1519.450 627.740 1520.230 627.880 ;
        RECT 1519.450 627.680 1519.770 627.740 ;
        RECT 1519.910 627.680 1520.230 627.740 ;
        RECT 1518.070 483.040 1518.390 483.100 ;
        RECT 1518.530 483.040 1518.850 483.100 ;
        RECT 1518.070 482.900 1518.850 483.040 ;
        RECT 1518.070 482.840 1518.390 482.900 ;
        RECT 1518.530 482.840 1518.850 482.900 ;
        RECT 1519.450 386.140 1519.770 386.200 ;
        RECT 1519.255 386.000 1519.770 386.140 ;
        RECT 1519.450 385.940 1519.770 386.000 ;
        RECT 1519.450 351.120 1519.770 351.180 ;
        RECT 1519.255 350.980 1519.770 351.120 ;
        RECT 1519.450 350.920 1519.770 350.980 ;
        RECT 1518.070 289.920 1518.390 289.980 ;
        RECT 1519.450 289.920 1519.770 289.980 ;
        RECT 1518.070 289.780 1519.770 289.920 ;
        RECT 1518.070 289.720 1518.390 289.780 ;
        RECT 1519.450 289.720 1519.770 289.780 ;
        RECT 1501.510 18.260 1501.830 18.320 ;
        RECT 1518.070 18.260 1518.390 18.320 ;
        RECT 1501.510 18.120 1518.390 18.260 ;
        RECT 1501.510 18.060 1501.830 18.120 ;
        RECT 1518.070 18.060 1518.390 18.120 ;
      LAYER via ;
        RECT 1519.020 1207.040 1519.280 1207.300 ;
        RECT 1519.480 1159.100 1519.740 1159.360 ;
        RECT 1519.480 724.240 1519.740 724.500 ;
        RECT 1519.940 724.240 1520.200 724.500 ;
        RECT 1519.480 627.680 1519.740 627.940 ;
        RECT 1519.940 627.680 1520.200 627.940 ;
        RECT 1518.100 482.840 1518.360 483.100 ;
        RECT 1518.560 482.840 1518.820 483.100 ;
        RECT 1519.480 385.940 1519.740 386.200 ;
        RECT 1519.480 350.920 1519.740 351.180 ;
        RECT 1518.100 289.720 1518.360 289.980 ;
        RECT 1519.480 289.720 1519.740 289.980 ;
        RECT 1501.540 18.060 1501.800 18.320 ;
        RECT 1518.100 18.060 1518.360 18.320 ;
      LAYER met2 ;
        RECT 1520.870 1221.010 1521.430 1228.680 ;
        RECT 1519.080 1220.870 1521.430 1221.010 ;
        RECT 1519.080 1207.330 1519.220 1220.870 ;
        RECT 1520.870 1219.680 1521.430 1220.870 ;
        RECT 1519.020 1207.010 1519.280 1207.330 ;
        RECT 1519.480 1159.070 1519.740 1159.390 ;
        RECT 1519.540 724.530 1519.680 1159.070 ;
        RECT 1519.480 724.210 1519.740 724.530 ;
        RECT 1519.940 724.210 1520.200 724.530 ;
        RECT 1520.000 689.930 1520.140 724.210 ;
        RECT 1519.540 689.790 1520.140 689.930 ;
        RECT 1519.540 627.970 1519.680 689.790 ;
        RECT 1519.480 627.650 1519.740 627.970 ;
        RECT 1519.940 627.650 1520.200 627.970 ;
        RECT 1520.000 593.370 1520.140 627.650 ;
        RECT 1519.540 593.230 1520.140 593.370 ;
        RECT 1519.540 531.490 1519.680 593.230 ;
        RECT 1519.540 531.350 1520.140 531.490 ;
        RECT 1520.000 483.325 1520.140 531.350 ;
        RECT 1518.090 482.955 1518.370 483.325 ;
        RECT 1518.100 482.810 1518.360 482.955 ;
        RECT 1518.560 482.810 1518.820 483.130 ;
        RECT 1519.930 482.955 1520.210 483.325 ;
        RECT 1518.620 434.930 1518.760 482.810 ;
        RECT 1518.620 434.790 1519.220 434.930 ;
        RECT 1519.080 386.650 1519.220 434.790 ;
        RECT 1519.080 386.510 1519.680 386.650 ;
        RECT 1519.540 386.230 1519.680 386.510 ;
        RECT 1519.480 385.910 1519.740 386.230 ;
        RECT 1519.480 350.890 1519.740 351.210 ;
        RECT 1519.540 290.010 1519.680 350.890 ;
        RECT 1518.100 289.690 1518.360 290.010 ;
        RECT 1519.480 289.690 1519.740 290.010 ;
        RECT 1518.160 18.350 1518.300 289.690 ;
        RECT 1501.540 18.030 1501.800 18.350 ;
        RECT 1518.100 18.030 1518.360 18.350 ;
        RECT 1501.600 2.400 1501.740 18.030 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
      LAYER via2 ;
        RECT 1518.090 483.000 1518.370 483.280 ;
        RECT 1519.930 483.000 1520.210 483.280 ;
      LAYER met3 ;
        RECT 1518.065 483.290 1518.395 483.305 ;
        RECT 1519.905 483.290 1520.235 483.305 ;
        RECT 1518.065 482.990 1520.235 483.290 ;
        RECT 1518.065 482.975 1518.395 482.990 ;
        RECT 1519.905 482.975 1520.235 482.990 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 1207.580 1524.830 1207.640 ;
        RECT 1530.030 1207.580 1530.350 1207.640 ;
        RECT 1524.510 1207.440 1530.350 1207.580 ;
        RECT 1524.510 1207.380 1524.830 1207.440 ;
        RECT 1530.030 1207.380 1530.350 1207.440 ;
        RECT 1518.990 20.640 1519.310 20.700 ;
        RECT 1524.510 20.640 1524.830 20.700 ;
        RECT 1518.990 20.500 1524.830 20.640 ;
        RECT 1518.990 20.440 1519.310 20.500 ;
        RECT 1524.510 20.440 1524.830 20.500 ;
      LAYER via ;
        RECT 1524.540 1207.380 1524.800 1207.640 ;
        RECT 1530.060 1207.380 1530.320 1207.640 ;
        RECT 1519.020 20.440 1519.280 20.700 ;
        RECT 1524.540 20.440 1524.800 20.700 ;
      LAYER met2 ;
        RECT 1530.070 1219.680 1530.630 1228.680 ;
        RECT 1530.120 1207.670 1530.260 1219.680 ;
        RECT 1524.540 1207.350 1524.800 1207.670 ;
        RECT 1530.060 1207.350 1530.320 1207.670 ;
        RECT 1524.600 20.730 1524.740 1207.350 ;
        RECT 1519.020 20.410 1519.280 20.730 ;
        RECT 1524.540 20.410 1524.800 20.730 ;
        RECT 1519.080 2.400 1519.220 20.410 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 1196.700 1111.290 1196.760 ;
        RECT 1116.030 1196.700 1116.350 1196.760 ;
        RECT 1110.970 1196.560 1116.350 1196.700 ;
        RECT 1110.970 1196.500 1111.290 1196.560 ;
        RECT 1116.030 1196.500 1116.350 1196.560 ;
        RECT 716.290 29.140 716.610 29.200 ;
        RECT 1110.970 29.140 1111.290 29.200 ;
        RECT 716.290 29.000 1111.290 29.140 ;
        RECT 716.290 28.940 716.610 29.000 ;
        RECT 1110.970 28.940 1111.290 29.000 ;
      LAYER via ;
        RECT 1111.000 1196.500 1111.260 1196.760 ;
        RECT 1116.060 1196.500 1116.320 1196.760 ;
        RECT 716.320 28.940 716.580 29.200 ;
        RECT 1111.000 28.940 1111.260 29.200 ;
      LAYER met2 ;
        RECT 1117.450 1220.330 1118.010 1228.680 ;
        RECT 1116.120 1220.190 1118.010 1220.330 ;
        RECT 1116.120 1196.790 1116.260 1220.190 ;
        RECT 1117.450 1219.680 1118.010 1220.190 ;
        RECT 1111.000 1196.470 1111.260 1196.790 ;
        RECT 1116.060 1196.470 1116.320 1196.790 ;
        RECT 1111.060 29.230 1111.200 1196.470 ;
        RECT 716.320 28.910 716.580 29.230 ;
        RECT 1111.000 28.910 1111.260 29.230 ;
        RECT 716.380 2.400 716.520 28.910 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1539.270 1220.330 1539.830 1228.680 ;
        RECT 1538.860 1220.190 1539.830 1220.330 ;
        RECT 1538.860 20.130 1539.000 1220.190 ;
        RECT 1539.270 1219.680 1539.830 1220.190 ;
        RECT 1537.020 19.990 1539.000 20.130 ;
        RECT 1537.020 2.400 1537.160 19.990 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1548.430 1207.580 1548.750 1207.640 ;
        RECT 1552.110 1207.580 1552.430 1207.640 ;
        RECT 1548.430 1207.440 1552.430 1207.580 ;
        RECT 1548.430 1207.380 1548.750 1207.440 ;
        RECT 1552.110 1207.380 1552.430 1207.440 ;
        RECT 1552.110 20.640 1552.430 20.700 ;
        RECT 1554.870 20.640 1555.190 20.700 ;
        RECT 1552.110 20.500 1555.190 20.640 ;
        RECT 1552.110 20.440 1552.430 20.500 ;
        RECT 1554.870 20.440 1555.190 20.500 ;
      LAYER via ;
        RECT 1548.460 1207.380 1548.720 1207.640 ;
        RECT 1552.140 1207.380 1552.400 1207.640 ;
        RECT 1552.140 20.440 1552.400 20.700 ;
        RECT 1554.900 20.440 1555.160 20.700 ;
      LAYER met2 ;
        RECT 1548.470 1219.680 1549.030 1228.680 ;
        RECT 1548.520 1207.670 1548.660 1219.680 ;
        RECT 1548.460 1207.350 1548.720 1207.670 ;
        RECT 1552.140 1207.350 1552.400 1207.670 ;
        RECT 1552.200 20.730 1552.340 1207.350 ;
        RECT 1552.140 20.410 1552.400 20.730 ;
        RECT 1554.900 20.410 1555.160 20.730 ;
        RECT 1554.960 2.400 1555.100 20.410 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 17.240 1559.330 17.300 ;
        RECT 1572.810 17.240 1573.130 17.300 ;
        RECT 1559.010 17.100 1573.130 17.240 ;
        RECT 1559.010 17.040 1559.330 17.100 ;
        RECT 1572.810 17.040 1573.130 17.100 ;
      LAYER via ;
        RECT 1559.040 17.040 1559.300 17.300 ;
        RECT 1572.840 17.040 1573.100 17.300 ;
      LAYER met2 ;
        RECT 1557.670 1220.330 1558.230 1228.680 ;
        RECT 1557.670 1220.190 1559.240 1220.330 ;
        RECT 1557.670 1219.680 1558.230 1220.190 ;
        RECT 1559.100 17.330 1559.240 1220.190 ;
        RECT 1559.040 17.010 1559.300 17.330 ;
        RECT 1572.840 17.010 1573.100 17.330 ;
        RECT 1572.900 2.400 1573.040 17.010 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1566.830 1213.020 1567.150 1213.080 ;
        RECT 1583.390 1213.020 1583.710 1213.080 ;
        RECT 1566.830 1212.880 1583.710 1213.020 ;
        RECT 1566.830 1212.820 1567.150 1212.880 ;
        RECT 1583.390 1212.820 1583.710 1212.880 ;
        RECT 1583.390 17.920 1583.710 17.980 ;
        RECT 1590.290 17.920 1590.610 17.980 ;
        RECT 1583.390 17.780 1590.610 17.920 ;
        RECT 1583.390 17.720 1583.710 17.780 ;
        RECT 1590.290 17.720 1590.610 17.780 ;
      LAYER via ;
        RECT 1566.860 1212.820 1567.120 1213.080 ;
        RECT 1583.420 1212.820 1583.680 1213.080 ;
        RECT 1583.420 17.720 1583.680 17.980 ;
        RECT 1590.320 17.720 1590.580 17.980 ;
      LAYER met2 ;
        RECT 1566.870 1219.680 1567.430 1228.680 ;
        RECT 1566.920 1213.110 1567.060 1219.680 ;
        RECT 1566.860 1212.790 1567.120 1213.110 ;
        RECT 1583.420 1212.790 1583.680 1213.110 ;
        RECT 1583.480 18.010 1583.620 1212.790 ;
        RECT 1583.420 17.690 1583.680 18.010 ;
        RECT 1590.320 17.690 1590.580 18.010 ;
        RECT 1590.380 2.400 1590.520 17.690 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.030 1211.660 1576.350 1211.720 ;
        RECT 1608.230 1211.660 1608.550 1211.720 ;
        RECT 1576.030 1211.520 1608.550 1211.660 ;
        RECT 1576.030 1211.460 1576.350 1211.520 ;
        RECT 1608.230 1211.460 1608.550 1211.520 ;
      LAYER via ;
        RECT 1576.060 1211.460 1576.320 1211.720 ;
        RECT 1608.260 1211.460 1608.520 1211.720 ;
      LAYER met2 ;
        RECT 1576.070 1219.680 1576.630 1228.680 ;
        RECT 1576.120 1211.750 1576.260 1219.680 ;
        RECT 1576.060 1211.430 1576.320 1211.750 ;
        RECT 1608.260 1211.430 1608.520 1211.750 ;
        RECT 1608.320 2.400 1608.460 1211.430 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1585.230 1208.260 1585.550 1208.320 ;
        RECT 1610.990 1208.260 1611.310 1208.320 ;
        RECT 1585.230 1208.120 1611.310 1208.260 ;
        RECT 1585.230 1208.060 1585.550 1208.120 ;
        RECT 1610.990 1208.060 1611.310 1208.120 ;
        RECT 1610.990 17.580 1611.310 17.640 ;
        RECT 1626.170 17.580 1626.490 17.640 ;
        RECT 1610.990 17.440 1626.490 17.580 ;
        RECT 1610.990 17.380 1611.310 17.440 ;
        RECT 1626.170 17.380 1626.490 17.440 ;
      LAYER via ;
        RECT 1585.260 1208.060 1585.520 1208.320 ;
        RECT 1611.020 1208.060 1611.280 1208.320 ;
        RECT 1611.020 17.380 1611.280 17.640 ;
        RECT 1626.200 17.380 1626.460 17.640 ;
      LAYER met2 ;
        RECT 1585.270 1219.680 1585.830 1228.680 ;
        RECT 1585.320 1208.350 1585.460 1219.680 ;
        RECT 1585.260 1208.030 1585.520 1208.350 ;
        RECT 1611.020 1208.030 1611.280 1208.350 ;
        RECT 1611.080 17.670 1611.220 1208.030 ;
        RECT 1611.020 17.350 1611.280 17.670 ;
        RECT 1626.200 17.350 1626.460 17.670 ;
        RECT 1626.260 2.400 1626.400 17.350 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1594.430 1208.600 1594.750 1208.660 ;
        RECT 1617.890 1208.600 1618.210 1208.660 ;
        RECT 1594.430 1208.460 1618.210 1208.600 ;
        RECT 1594.430 1208.400 1594.750 1208.460 ;
        RECT 1617.890 1208.400 1618.210 1208.460 ;
        RECT 1617.890 16.560 1618.210 16.620 ;
        RECT 1644.110 16.560 1644.430 16.620 ;
        RECT 1617.890 16.420 1644.430 16.560 ;
        RECT 1617.890 16.360 1618.210 16.420 ;
        RECT 1644.110 16.360 1644.430 16.420 ;
      LAYER via ;
        RECT 1594.460 1208.400 1594.720 1208.660 ;
        RECT 1617.920 1208.400 1618.180 1208.660 ;
        RECT 1617.920 16.360 1618.180 16.620 ;
        RECT 1644.140 16.360 1644.400 16.620 ;
      LAYER met2 ;
        RECT 1594.470 1219.680 1595.030 1228.680 ;
        RECT 1594.520 1208.690 1594.660 1219.680 ;
        RECT 1594.460 1208.370 1594.720 1208.690 ;
        RECT 1617.920 1208.370 1618.180 1208.690 ;
        RECT 1617.980 16.650 1618.120 1208.370 ;
        RECT 1617.920 16.330 1618.180 16.650 ;
        RECT 1644.140 16.330 1644.400 16.650 ;
        RECT 1644.200 2.400 1644.340 16.330 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1603.170 1207.580 1603.490 1207.640 ;
        RECT 1607.310 1207.580 1607.630 1207.640 ;
        RECT 1603.170 1207.440 1607.630 1207.580 ;
        RECT 1603.170 1207.380 1603.490 1207.440 ;
        RECT 1607.310 1207.380 1607.630 1207.440 ;
        RECT 1607.310 20.300 1607.630 20.360 ;
        RECT 1662.050 20.300 1662.370 20.360 ;
        RECT 1607.310 20.160 1662.370 20.300 ;
        RECT 1607.310 20.100 1607.630 20.160 ;
        RECT 1662.050 20.100 1662.370 20.160 ;
      LAYER via ;
        RECT 1603.200 1207.380 1603.460 1207.640 ;
        RECT 1607.340 1207.380 1607.600 1207.640 ;
        RECT 1607.340 20.100 1607.600 20.360 ;
        RECT 1662.080 20.100 1662.340 20.360 ;
      LAYER met2 ;
        RECT 1603.210 1219.680 1603.770 1228.680 ;
        RECT 1603.260 1207.670 1603.400 1219.680 ;
        RECT 1603.200 1207.350 1603.460 1207.670 ;
        RECT 1607.340 1207.350 1607.600 1207.670 ;
        RECT 1607.400 20.390 1607.540 1207.350 ;
        RECT 1607.340 20.070 1607.600 20.390 ;
        RECT 1662.080 20.070 1662.340 20.390 ;
        RECT 1662.140 2.400 1662.280 20.070 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.750 18.260 1614.070 18.320 ;
        RECT 1679.530 18.260 1679.850 18.320 ;
        RECT 1613.750 18.120 1679.850 18.260 ;
        RECT 1613.750 18.060 1614.070 18.120 ;
        RECT 1679.530 18.060 1679.850 18.120 ;
      LAYER via ;
        RECT 1613.780 18.060 1614.040 18.320 ;
        RECT 1679.560 18.060 1679.820 18.320 ;
      LAYER met2 ;
        RECT 1612.410 1220.330 1612.970 1228.680 ;
        RECT 1612.410 1220.190 1613.980 1220.330 ;
        RECT 1612.410 1219.680 1612.970 1220.190 ;
        RECT 1613.840 18.350 1613.980 1220.190 ;
        RECT 1613.780 18.030 1614.040 18.350 ;
        RECT 1679.560 18.030 1679.820 18.350 ;
        RECT 1679.620 2.400 1679.760 18.030 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1621.570 1207.580 1621.890 1207.640 ;
        RECT 1628.010 1207.580 1628.330 1207.640 ;
        RECT 1621.570 1207.440 1628.330 1207.580 ;
        RECT 1621.570 1207.380 1621.890 1207.440 ;
        RECT 1628.010 1207.380 1628.330 1207.440 ;
        RECT 1628.010 17.580 1628.330 17.640 ;
        RECT 1697.470 17.580 1697.790 17.640 ;
        RECT 1628.010 17.440 1697.790 17.580 ;
        RECT 1628.010 17.380 1628.330 17.440 ;
        RECT 1697.470 17.380 1697.790 17.440 ;
      LAYER via ;
        RECT 1621.600 1207.380 1621.860 1207.640 ;
        RECT 1628.040 1207.380 1628.300 1207.640 ;
        RECT 1628.040 17.380 1628.300 17.640 ;
        RECT 1697.500 17.380 1697.760 17.640 ;
      LAYER met2 ;
        RECT 1621.610 1219.680 1622.170 1228.680 ;
        RECT 1621.660 1207.670 1621.800 1219.680 ;
        RECT 1621.600 1207.350 1621.860 1207.670 ;
        RECT 1628.040 1207.350 1628.300 1207.670 ;
        RECT 1628.100 17.670 1628.240 1207.350 ;
        RECT 1628.040 17.350 1628.300 17.670 ;
        RECT 1697.500 17.350 1697.760 17.670 ;
        RECT 1697.560 2.400 1697.700 17.350 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 734.230 28.800 734.550 28.860 ;
        RECT 1124.770 28.800 1125.090 28.860 ;
        RECT 734.230 28.660 1125.090 28.800 ;
        RECT 734.230 28.600 734.550 28.660 ;
        RECT 1124.770 28.600 1125.090 28.660 ;
      LAYER via ;
        RECT 734.260 28.600 734.520 28.860 ;
        RECT 1124.800 28.600 1125.060 28.860 ;
      LAYER met2 ;
        RECT 1126.650 1220.330 1127.210 1228.680 ;
        RECT 1124.860 1220.190 1127.210 1220.330 ;
        RECT 1124.860 28.890 1125.000 1220.190 ;
        RECT 1126.650 1219.680 1127.210 1220.190 ;
        RECT 734.260 28.570 734.520 28.890 ;
        RECT 1124.800 28.570 1125.060 28.890 ;
        RECT 734.320 2.400 734.460 28.570 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1630.770 1207.580 1631.090 1207.640 ;
        RECT 1634.910 1207.580 1635.230 1207.640 ;
        RECT 1630.770 1207.440 1635.230 1207.580 ;
        RECT 1630.770 1207.380 1631.090 1207.440 ;
        RECT 1634.910 1207.380 1635.230 1207.440 ;
        RECT 1634.910 17.240 1635.230 17.300 ;
        RECT 1715.410 17.240 1715.730 17.300 ;
        RECT 1634.910 17.100 1715.730 17.240 ;
        RECT 1634.910 17.040 1635.230 17.100 ;
        RECT 1715.410 17.040 1715.730 17.100 ;
      LAYER via ;
        RECT 1630.800 1207.380 1631.060 1207.640 ;
        RECT 1634.940 1207.380 1635.200 1207.640 ;
        RECT 1634.940 17.040 1635.200 17.300 ;
        RECT 1715.440 17.040 1715.700 17.300 ;
      LAYER met2 ;
        RECT 1630.810 1219.680 1631.370 1228.680 ;
        RECT 1630.860 1207.670 1631.000 1219.680 ;
        RECT 1630.800 1207.350 1631.060 1207.670 ;
        RECT 1634.940 1207.350 1635.200 1207.670 ;
        RECT 1635.000 17.330 1635.140 1207.350 ;
        RECT 1634.940 17.010 1635.200 17.330 ;
        RECT 1715.440 17.010 1715.700 17.330 ;
        RECT 1715.500 2.400 1715.640 17.010 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1641.350 19.620 1641.670 19.680 ;
        RECT 1733.350 19.620 1733.670 19.680 ;
        RECT 1641.350 19.480 1733.670 19.620 ;
        RECT 1641.350 19.420 1641.670 19.480 ;
        RECT 1733.350 19.420 1733.670 19.480 ;
      LAYER via ;
        RECT 1641.380 19.420 1641.640 19.680 ;
        RECT 1733.380 19.420 1733.640 19.680 ;
      LAYER met2 ;
        RECT 1640.010 1220.330 1640.570 1228.680 ;
        RECT 1640.010 1220.190 1641.580 1220.330 ;
        RECT 1640.010 1219.680 1640.570 1220.190 ;
        RECT 1641.440 19.710 1641.580 1220.190 ;
        RECT 1641.380 19.390 1641.640 19.710 ;
        RECT 1733.380 19.390 1733.640 19.710 ;
        RECT 1733.440 2.400 1733.580 19.390 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1649.170 1213.700 1649.490 1213.760 ;
        RECT 1700.690 1213.700 1701.010 1213.760 ;
        RECT 1649.170 1213.560 1701.010 1213.700 ;
        RECT 1649.170 1213.500 1649.490 1213.560 ;
        RECT 1700.690 1213.500 1701.010 1213.560 ;
        RECT 1700.690 16.900 1701.010 16.960 ;
        RECT 1700.690 16.760 1704.140 16.900 ;
        RECT 1700.690 16.700 1701.010 16.760 ;
        RECT 1704.000 16.560 1704.140 16.760 ;
        RECT 1751.290 16.560 1751.610 16.620 ;
        RECT 1704.000 16.420 1751.610 16.560 ;
        RECT 1751.290 16.360 1751.610 16.420 ;
      LAYER via ;
        RECT 1649.200 1213.500 1649.460 1213.760 ;
        RECT 1700.720 1213.500 1700.980 1213.760 ;
        RECT 1700.720 16.700 1700.980 16.960 ;
        RECT 1751.320 16.360 1751.580 16.620 ;
      LAYER met2 ;
        RECT 1649.210 1219.680 1649.770 1228.680 ;
        RECT 1649.260 1213.790 1649.400 1219.680 ;
        RECT 1649.200 1213.470 1649.460 1213.790 ;
        RECT 1700.720 1213.470 1700.980 1213.790 ;
        RECT 1700.780 16.990 1700.920 1213.470 ;
        RECT 1700.720 16.670 1700.980 16.990 ;
        RECT 1751.320 16.330 1751.580 16.650 ;
        RECT 1751.380 2.400 1751.520 16.330 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1658.370 1214.040 1658.690 1214.100 ;
        RECT 1707.590 1214.040 1707.910 1214.100 ;
        RECT 1658.370 1213.900 1707.910 1214.040 ;
        RECT 1658.370 1213.840 1658.690 1213.900 ;
        RECT 1707.590 1213.840 1707.910 1213.900 ;
        RECT 1768.770 16.900 1769.090 16.960 ;
        RECT 1751.840 16.760 1769.090 16.900 ;
        RECT 1707.590 15.880 1707.910 15.940 ;
        RECT 1751.840 15.880 1751.980 16.760 ;
        RECT 1768.770 16.700 1769.090 16.760 ;
        RECT 1707.590 15.740 1751.980 15.880 ;
        RECT 1707.590 15.680 1707.910 15.740 ;
      LAYER via ;
        RECT 1658.400 1213.840 1658.660 1214.100 ;
        RECT 1707.620 1213.840 1707.880 1214.100 ;
        RECT 1707.620 15.680 1707.880 15.940 ;
        RECT 1768.800 16.700 1769.060 16.960 ;
      LAYER met2 ;
        RECT 1658.410 1219.680 1658.970 1228.680 ;
        RECT 1658.460 1214.130 1658.600 1219.680 ;
        RECT 1658.400 1213.810 1658.660 1214.130 ;
        RECT 1707.620 1213.810 1707.880 1214.130 ;
        RECT 1707.680 15.970 1707.820 1213.810 ;
        RECT 1768.800 16.670 1769.060 16.990 ;
        RECT 1707.620 15.650 1707.880 15.970 ;
        RECT 1768.860 2.400 1769.000 16.670 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1714.565 1212.525 1714.735 1214.735 ;
        RECT 1738.485 1212.865 1738.655 1214.735 ;
        RECT 1752.745 1213.205 1753.835 1213.375 ;
        RECT 1753.665 1209.635 1753.835 1213.205 ;
        RECT 1753.665 1209.465 1754.755 1209.635 ;
        RECT 1775.745 1207.085 1775.915 1209.635 ;
      LAYER mcon ;
        RECT 1714.565 1214.565 1714.735 1214.735 ;
        RECT 1738.485 1214.565 1738.655 1214.735 ;
        RECT 1754.585 1209.465 1754.755 1209.635 ;
        RECT 1775.745 1209.465 1775.915 1209.635 ;
      LAYER met1 ;
        RECT 1714.505 1214.720 1714.795 1214.765 ;
        RECT 1738.425 1214.720 1738.715 1214.765 ;
        RECT 1714.505 1214.580 1738.715 1214.720 ;
        RECT 1714.505 1214.535 1714.795 1214.580 ;
        RECT 1738.425 1214.535 1738.715 1214.580 ;
        RECT 1752.685 1213.175 1752.975 1213.405 ;
        RECT 1738.425 1213.020 1738.715 1213.065 ;
        RECT 1752.760 1213.020 1752.900 1213.175 ;
        RECT 1738.425 1212.880 1752.900 1213.020 ;
        RECT 1738.425 1212.835 1738.715 1212.880 ;
        RECT 1667.570 1212.680 1667.890 1212.740 ;
        RECT 1714.505 1212.680 1714.795 1212.725 ;
        RECT 1667.570 1212.540 1714.795 1212.680 ;
        RECT 1667.570 1212.480 1667.890 1212.540 ;
        RECT 1714.505 1212.495 1714.795 1212.540 ;
        RECT 1754.525 1209.620 1754.815 1209.665 ;
        RECT 1775.685 1209.620 1775.975 1209.665 ;
        RECT 1754.525 1209.480 1775.975 1209.620 ;
        RECT 1754.525 1209.435 1754.815 1209.480 ;
        RECT 1775.685 1209.435 1775.975 1209.480 ;
        RECT 1775.685 1207.240 1775.975 1207.285 ;
        RECT 1781.650 1207.240 1781.970 1207.300 ;
        RECT 1775.685 1207.100 1781.970 1207.240 ;
        RECT 1775.685 1207.055 1775.975 1207.100 ;
        RECT 1781.650 1207.040 1781.970 1207.100 ;
        RECT 1781.650 61.920 1781.970 62.180 ;
        RECT 1781.740 61.780 1781.880 61.920 ;
        RECT 1786.710 61.780 1787.030 61.840 ;
        RECT 1781.740 61.640 1787.030 61.780 ;
        RECT 1786.710 61.580 1787.030 61.640 ;
      LAYER via ;
        RECT 1667.600 1212.480 1667.860 1212.740 ;
        RECT 1781.680 1207.040 1781.940 1207.300 ;
        RECT 1781.680 61.920 1781.940 62.180 ;
        RECT 1786.740 61.580 1787.000 61.840 ;
      LAYER met2 ;
        RECT 1667.610 1219.680 1668.170 1228.680 ;
        RECT 1667.660 1212.770 1667.800 1219.680 ;
        RECT 1667.600 1212.450 1667.860 1212.770 ;
        RECT 1781.680 1207.010 1781.940 1207.330 ;
        RECT 1781.740 62.210 1781.880 1207.010 ;
        RECT 1781.680 61.890 1781.940 62.210 ;
        RECT 1786.740 61.550 1787.000 61.870 ;
        RECT 1786.800 2.400 1786.940 61.550 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1720.085 1208.275 1720.255 1209.635 ;
        RECT 1721.005 1208.275 1721.175 1208.615 ;
        RECT 1720.085 1208.105 1721.175 1208.275 ;
      LAYER mcon ;
        RECT 1720.085 1209.465 1720.255 1209.635 ;
        RECT 1721.005 1208.445 1721.175 1208.615 ;
      LAYER met1 ;
        RECT 1676.770 1209.620 1677.090 1209.680 ;
        RECT 1720.025 1209.620 1720.315 1209.665 ;
        RECT 1676.770 1209.480 1720.315 1209.620 ;
        RECT 1676.770 1209.420 1677.090 1209.480 ;
        RECT 1720.025 1209.435 1720.315 1209.480 ;
        RECT 1720.945 1208.600 1721.235 1208.645 ;
        RECT 1728.290 1208.600 1728.610 1208.660 ;
        RECT 1720.945 1208.460 1728.610 1208.600 ;
        RECT 1720.945 1208.415 1721.235 1208.460 ;
        RECT 1728.290 1208.400 1728.610 1208.460 ;
        RECT 1728.290 20.640 1728.610 20.700 ;
        RECT 1804.650 20.640 1804.970 20.700 ;
        RECT 1728.290 20.500 1804.970 20.640 ;
        RECT 1728.290 20.440 1728.610 20.500 ;
        RECT 1804.650 20.440 1804.970 20.500 ;
      LAYER via ;
        RECT 1676.800 1209.420 1677.060 1209.680 ;
        RECT 1728.320 1208.400 1728.580 1208.660 ;
        RECT 1728.320 20.440 1728.580 20.700 ;
        RECT 1804.680 20.440 1804.940 20.700 ;
      LAYER met2 ;
        RECT 1676.810 1219.680 1677.370 1228.680 ;
        RECT 1676.860 1209.710 1677.000 1219.680 ;
        RECT 1676.800 1209.390 1677.060 1209.710 ;
        RECT 1728.320 1208.370 1728.580 1208.690 ;
        RECT 1728.380 20.730 1728.520 1208.370 ;
        RECT 1728.320 20.410 1728.580 20.730 ;
        RECT 1804.680 20.410 1804.940 20.730 ;
        RECT 1804.740 2.400 1804.880 20.410 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.970 1208.260 1686.290 1208.320 ;
        RECT 1685.970 1208.120 1694.940 1208.260 ;
        RECT 1685.970 1208.060 1686.290 1208.120 ;
        RECT 1694.800 1207.920 1694.940 1208.120 ;
        RECT 1783.490 1207.920 1783.810 1207.980 ;
        RECT 1694.800 1207.780 1783.810 1207.920 ;
        RECT 1783.490 1207.720 1783.810 1207.780 ;
        RECT 1783.490 18.940 1783.810 19.000 ;
        RECT 1822.590 18.940 1822.910 19.000 ;
        RECT 1783.490 18.800 1822.910 18.940 ;
        RECT 1783.490 18.740 1783.810 18.800 ;
        RECT 1822.590 18.740 1822.910 18.800 ;
      LAYER via ;
        RECT 1686.000 1208.060 1686.260 1208.320 ;
        RECT 1783.520 1207.720 1783.780 1207.980 ;
        RECT 1783.520 18.740 1783.780 19.000 ;
        RECT 1822.620 18.740 1822.880 19.000 ;
      LAYER met2 ;
        RECT 1686.010 1219.680 1686.570 1228.680 ;
        RECT 1686.060 1208.350 1686.200 1219.680 ;
        RECT 1686.000 1208.030 1686.260 1208.350 ;
        RECT 1783.520 1207.690 1783.780 1208.010 ;
        RECT 1783.580 19.030 1783.720 1207.690 ;
        RECT 1783.520 18.710 1783.780 19.030 ;
        RECT 1822.620 18.710 1822.880 19.030 ;
        RECT 1822.680 2.400 1822.820 18.710 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1695.170 1208.260 1695.490 1208.320 ;
        RECT 1790.390 1208.260 1790.710 1208.320 ;
        RECT 1695.170 1208.120 1790.710 1208.260 ;
        RECT 1695.170 1208.060 1695.490 1208.120 ;
        RECT 1790.390 1208.060 1790.710 1208.120 ;
        RECT 1790.390 16.560 1790.710 16.620 ;
        RECT 1840.070 16.560 1840.390 16.620 ;
        RECT 1790.390 16.420 1840.390 16.560 ;
        RECT 1790.390 16.360 1790.710 16.420 ;
        RECT 1840.070 16.360 1840.390 16.420 ;
      LAYER via ;
        RECT 1695.200 1208.060 1695.460 1208.320 ;
        RECT 1790.420 1208.060 1790.680 1208.320 ;
        RECT 1790.420 16.360 1790.680 16.620 ;
        RECT 1840.100 16.360 1840.360 16.620 ;
      LAYER met2 ;
        RECT 1695.210 1219.680 1695.770 1228.680 ;
        RECT 1695.260 1208.350 1695.400 1219.680 ;
        RECT 1695.200 1208.030 1695.460 1208.350 ;
        RECT 1790.420 1208.030 1790.680 1208.350 ;
        RECT 1790.480 16.650 1790.620 1208.030 ;
        RECT 1790.420 16.330 1790.680 16.650 ;
        RECT 1840.100 16.330 1840.360 16.650 ;
        RECT 1840.160 2.400 1840.300 16.330 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1753.205 1207.595 1753.375 1212.695 ;
        RECT 1752.745 1207.425 1753.375 1207.595 ;
      LAYER mcon ;
        RECT 1753.205 1212.525 1753.375 1212.695 ;
      LAYER met1 ;
        RECT 1753.145 1212.680 1753.435 1212.725 ;
        RECT 1753.145 1212.540 1776.820 1212.680 ;
        RECT 1753.145 1212.495 1753.435 1212.540 ;
        RECT 1776.680 1212.340 1776.820 1212.540 ;
        RECT 1797.290 1212.340 1797.610 1212.400 ;
        RECT 1776.680 1212.200 1797.610 1212.340 ;
        RECT 1797.290 1212.140 1797.610 1212.200 ;
        RECT 1704.370 1207.580 1704.690 1207.640 ;
        RECT 1752.685 1207.580 1752.975 1207.625 ;
        RECT 1704.370 1207.440 1740.480 1207.580 ;
        RECT 1704.370 1207.380 1704.690 1207.440 ;
        RECT 1740.340 1207.240 1740.480 1207.440 ;
        RECT 1745.860 1207.440 1752.975 1207.580 ;
        RECT 1745.860 1207.240 1746.000 1207.440 ;
        RECT 1752.685 1207.395 1752.975 1207.440 ;
        RECT 1740.340 1207.100 1746.000 1207.240 ;
        RECT 1797.290 16.900 1797.610 16.960 ;
        RECT 1858.010 16.900 1858.330 16.960 ;
        RECT 1797.290 16.760 1858.330 16.900 ;
        RECT 1797.290 16.700 1797.610 16.760 ;
        RECT 1858.010 16.700 1858.330 16.760 ;
      LAYER via ;
        RECT 1797.320 1212.140 1797.580 1212.400 ;
        RECT 1704.400 1207.380 1704.660 1207.640 ;
        RECT 1797.320 16.700 1797.580 16.960 ;
        RECT 1858.040 16.700 1858.300 16.960 ;
      LAYER met2 ;
        RECT 1704.410 1219.680 1704.970 1228.680 ;
        RECT 1704.460 1207.670 1704.600 1219.680 ;
        RECT 1797.320 1212.110 1797.580 1212.430 ;
        RECT 1704.400 1207.350 1704.660 1207.670 ;
        RECT 1797.380 16.990 1797.520 1212.110 ;
        RECT 1797.320 16.670 1797.580 16.990 ;
        RECT 1858.040 16.670 1858.300 16.990 ;
        RECT 1858.100 2.400 1858.240 16.670 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1713.570 1210.300 1713.890 1210.360 ;
        RECT 1870.430 1210.300 1870.750 1210.360 ;
        RECT 1713.570 1210.160 1870.750 1210.300 ;
        RECT 1713.570 1210.100 1713.890 1210.160 ;
        RECT 1870.430 1210.100 1870.750 1210.160 ;
        RECT 1870.430 7.720 1870.750 7.780 ;
        RECT 1875.950 7.720 1876.270 7.780 ;
        RECT 1870.430 7.580 1876.270 7.720 ;
        RECT 1870.430 7.520 1870.750 7.580 ;
        RECT 1875.950 7.520 1876.270 7.580 ;
      LAYER via ;
        RECT 1713.600 1210.100 1713.860 1210.360 ;
        RECT 1870.460 1210.100 1870.720 1210.360 ;
        RECT 1870.460 7.520 1870.720 7.780 ;
        RECT 1875.980 7.520 1876.240 7.780 ;
      LAYER met2 ;
        RECT 1713.610 1219.680 1714.170 1228.680 ;
        RECT 1713.660 1210.390 1713.800 1219.680 ;
        RECT 1713.600 1210.070 1713.860 1210.390 ;
        RECT 1870.460 1210.070 1870.720 1210.390 ;
        RECT 1870.520 7.810 1870.660 1210.070 ;
        RECT 1870.460 7.490 1870.720 7.810 ;
        RECT 1875.980 7.490 1876.240 7.810 ;
        RECT 1876.040 2.400 1876.180 7.490 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1133.125 462.485 1133.295 469.115 ;
        RECT 1132.665 276.165 1132.835 414.035 ;
      LAYER mcon ;
        RECT 1133.125 468.945 1133.295 469.115 ;
        RECT 1132.665 413.865 1132.835 414.035 ;
      LAYER met1 ;
        RECT 1133.050 1159.300 1133.370 1159.360 ;
        RECT 1133.970 1159.300 1134.290 1159.360 ;
        RECT 1133.050 1159.160 1134.290 1159.300 ;
        RECT 1133.050 1159.100 1133.370 1159.160 ;
        RECT 1133.970 1159.100 1134.290 1159.160 ;
        RECT 1132.590 1014.460 1132.910 1014.520 ;
        RECT 1133.050 1014.460 1133.370 1014.520 ;
        RECT 1132.590 1014.320 1133.370 1014.460 ;
        RECT 1132.590 1014.260 1132.910 1014.320 ;
        RECT 1133.050 1014.260 1133.370 1014.320 ;
        RECT 1133.050 1007.320 1133.370 1007.380 ;
        RECT 1133.970 1007.320 1134.290 1007.380 ;
        RECT 1133.050 1007.180 1134.290 1007.320 ;
        RECT 1133.050 1007.120 1133.370 1007.180 ;
        RECT 1133.970 1007.120 1134.290 1007.180 ;
        RECT 1133.510 1000.520 1133.830 1000.580 ;
        RECT 1133.970 1000.520 1134.290 1000.580 ;
        RECT 1133.510 1000.380 1134.290 1000.520 ;
        RECT 1133.510 1000.320 1133.830 1000.380 ;
        RECT 1133.970 1000.320 1134.290 1000.380 ;
        RECT 1132.130 952.240 1132.450 952.300 ;
        RECT 1133.970 952.240 1134.290 952.300 ;
        RECT 1132.130 952.100 1134.290 952.240 ;
        RECT 1132.130 952.040 1132.450 952.100 ;
        RECT 1133.970 952.040 1134.290 952.100 ;
        RECT 1133.050 869.960 1133.370 870.020 ;
        RECT 1132.680 869.820 1133.370 869.960 ;
        RECT 1132.680 869.340 1132.820 869.820 ;
        RECT 1133.050 869.760 1133.370 869.820 ;
        RECT 1132.590 869.080 1132.910 869.340 ;
        RECT 1132.590 772.720 1132.910 772.780 ;
        RECT 1133.050 772.720 1133.370 772.780 ;
        RECT 1132.590 772.580 1133.370 772.720 ;
        RECT 1132.590 772.520 1132.910 772.580 ;
        RECT 1133.050 772.520 1133.370 772.580 ;
        RECT 1133.050 469.100 1133.370 469.160 ;
        RECT 1132.855 468.960 1133.370 469.100 ;
        RECT 1133.050 468.900 1133.370 468.960 ;
        RECT 1133.050 462.640 1133.370 462.700 ;
        RECT 1132.855 462.500 1133.370 462.640 ;
        RECT 1133.050 462.440 1133.370 462.500 ;
        RECT 1132.605 414.020 1132.895 414.065 ;
        RECT 1133.050 414.020 1133.370 414.080 ;
        RECT 1132.605 413.880 1133.370 414.020 ;
        RECT 1132.605 413.835 1132.895 413.880 ;
        RECT 1133.050 413.820 1133.370 413.880 ;
        RECT 1132.605 276.320 1132.895 276.365 ;
        RECT 1133.510 276.320 1133.830 276.380 ;
        RECT 1132.605 276.180 1133.830 276.320 ;
        RECT 1132.605 276.135 1132.895 276.180 ;
        RECT 1133.510 276.120 1133.830 276.180 ;
        RECT 752.170 28.460 752.490 28.520 ;
        RECT 1132.590 28.460 1132.910 28.520 ;
        RECT 752.170 28.320 1132.910 28.460 ;
        RECT 752.170 28.260 752.490 28.320 ;
        RECT 1132.590 28.260 1132.910 28.320 ;
      LAYER via ;
        RECT 1133.080 1159.100 1133.340 1159.360 ;
        RECT 1134.000 1159.100 1134.260 1159.360 ;
        RECT 1132.620 1014.260 1132.880 1014.520 ;
        RECT 1133.080 1014.260 1133.340 1014.520 ;
        RECT 1133.080 1007.120 1133.340 1007.380 ;
        RECT 1134.000 1007.120 1134.260 1007.380 ;
        RECT 1133.540 1000.320 1133.800 1000.580 ;
        RECT 1134.000 1000.320 1134.260 1000.580 ;
        RECT 1132.160 952.040 1132.420 952.300 ;
        RECT 1134.000 952.040 1134.260 952.300 ;
        RECT 1133.080 869.760 1133.340 870.020 ;
        RECT 1132.620 869.080 1132.880 869.340 ;
        RECT 1132.620 772.520 1132.880 772.780 ;
        RECT 1133.080 772.520 1133.340 772.780 ;
        RECT 1133.080 468.900 1133.340 469.160 ;
        RECT 1133.080 462.440 1133.340 462.700 ;
        RECT 1133.080 413.820 1133.340 414.080 ;
        RECT 1133.540 276.120 1133.800 276.380 ;
        RECT 752.200 28.260 752.460 28.520 ;
        RECT 1132.620 28.260 1132.880 28.520 ;
      LAYER met2 ;
        RECT 1135.850 1221.010 1136.410 1228.680 ;
        RECT 1134.060 1220.870 1136.410 1221.010 ;
        RECT 1134.060 1159.390 1134.200 1220.870 ;
        RECT 1135.850 1219.680 1136.410 1220.870 ;
        RECT 1133.080 1159.070 1133.340 1159.390 ;
        RECT 1134.000 1159.070 1134.260 1159.390 ;
        RECT 1133.140 1076.850 1133.280 1159.070 ;
        RECT 1132.680 1076.710 1133.280 1076.850 ;
        RECT 1132.680 1014.550 1132.820 1076.710 ;
        RECT 1132.620 1014.230 1132.880 1014.550 ;
        RECT 1133.080 1014.230 1133.340 1014.550 ;
        RECT 1133.140 1007.410 1133.280 1014.230 ;
        RECT 1133.080 1007.090 1133.340 1007.410 ;
        RECT 1134.000 1007.090 1134.260 1007.410 ;
        RECT 1134.060 1000.610 1134.200 1007.090 ;
        RECT 1133.540 1000.290 1133.800 1000.610 ;
        RECT 1134.000 1000.290 1134.260 1000.610 ;
        RECT 1133.600 953.205 1133.740 1000.290 ;
        RECT 1133.530 952.835 1133.810 953.205 ;
        RECT 1132.150 952.155 1132.430 952.525 ;
        RECT 1132.160 952.010 1132.420 952.155 ;
        RECT 1134.000 952.010 1134.260 952.330 ;
        RECT 1134.060 904.245 1134.200 952.010 ;
        RECT 1133.070 903.875 1133.350 904.245 ;
        RECT 1133.990 903.875 1134.270 904.245 ;
        RECT 1133.140 870.050 1133.280 903.875 ;
        RECT 1133.080 869.730 1133.340 870.050 ;
        RECT 1132.620 869.050 1132.880 869.370 ;
        RECT 1132.680 773.685 1132.820 869.050 ;
        RECT 1132.610 773.315 1132.890 773.685 ;
        RECT 1132.610 772.635 1132.890 773.005 ;
        RECT 1132.620 772.490 1132.880 772.635 ;
        RECT 1133.080 772.490 1133.340 772.810 ;
        RECT 1133.140 724.610 1133.280 772.490 ;
        RECT 1133.140 724.470 1133.740 724.610 ;
        RECT 1133.600 676.445 1133.740 724.470 ;
        RECT 1132.610 676.075 1132.890 676.445 ;
        RECT 1133.530 676.075 1133.810 676.445 ;
        RECT 1132.680 628.050 1132.820 676.075 ;
        RECT 1132.680 627.910 1133.280 628.050 ;
        RECT 1133.140 469.190 1133.280 627.910 ;
        RECT 1133.080 468.870 1133.340 469.190 ;
        RECT 1133.080 462.410 1133.340 462.730 ;
        RECT 1133.140 414.110 1133.280 462.410 ;
        RECT 1133.080 413.790 1133.340 414.110 ;
        RECT 1133.540 276.090 1133.800 276.410 ;
        RECT 1133.600 193.530 1133.740 276.090 ;
        RECT 1133.140 193.390 1133.740 193.530 ;
        RECT 1133.140 193.020 1133.280 193.390 ;
        RECT 1132.680 192.880 1133.280 193.020 ;
        RECT 1132.680 137.770 1132.820 192.880 ;
        RECT 1132.680 137.630 1133.280 137.770 ;
        RECT 1133.140 90.170 1133.280 137.630 ;
        RECT 1132.680 90.030 1133.280 90.170 ;
        RECT 1132.680 28.550 1132.820 90.030 ;
        RECT 752.200 28.230 752.460 28.550 ;
        RECT 1132.620 28.230 1132.880 28.550 ;
        RECT 752.260 2.400 752.400 28.230 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 1133.530 952.880 1133.810 953.160 ;
        RECT 1132.150 952.200 1132.430 952.480 ;
        RECT 1133.070 903.920 1133.350 904.200 ;
        RECT 1133.990 903.920 1134.270 904.200 ;
        RECT 1132.610 773.360 1132.890 773.640 ;
        RECT 1132.610 772.680 1132.890 772.960 ;
        RECT 1132.610 676.120 1132.890 676.400 ;
        RECT 1133.530 676.120 1133.810 676.400 ;
      LAYER met3 ;
        RECT 1133.505 953.170 1133.835 953.185 ;
        RECT 1131.910 952.870 1133.835 953.170 ;
        RECT 1131.910 952.505 1132.210 952.870 ;
        RECT 1133.505 952.855 1133.835 952.870 ;
        RECT 1131.910 952.190 1132.455 952.505 ;
        RECT 1132.125 952.175 1132.455 952.190 ;
        RECT 1133.045 904.210 1133.375 904.225 ;
        RECT 1133.965 904.210 1134.295 904.225 ;
        RECT 1133.045 903.910 1134.295 904.210 ;
        RECT 1133.045 903.895 1133.375 903.910 ;
        RECT 1133.965 903.895 1134.295 903.910 ;
        RECT 1132.585 773.650 1132.915 773.665 ;
        RECT 1132.585 773.335 1133.130 773.650 ;
        RECT 1132.830 772.985 1133.130 773.335 ;
        RECT 1132.585 772.670 1133.130 772.985 ;
        RECT 1132.585 772.655 1132.915 772.670 ;
        RECT 1132.585 676.410 1132.915 676.425 ;
        RECT 1133.505 676.410 1133.835 676.425 ;
        RECT 1132.585 676.110 1133.835 676.410 ;
        RECT 1132.585 676.095 1132.915 676.110 ;
        RECT 1133.505 676.095 1133.835 676.110 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.610 17.240 1724.930 17.300 ;
        RECT 1893.890 17.240 1894.210 17.300 ;
        RECT 1724.610 17.100 1894.210 17.240 ;
        RECT 1724.610 17.040 1724.930 17.100 ;
        RECT 1893.890 17.040 1894.210 17.100 ;
      LAYER via ;
        RECT 1724.640 17.040 1724.900 17.300 ;
        RECT 1893.920 17.040 1894.180 17.300 ;
      LAYER met2 ;
        RECT 1722.810 1220.330 1723.370 1228.680 ;
        RECT 1722.810 1220.190 1724.840 1220.330 ;
        RECT 1722.810 1219.680 1723.370 1220.190 ;
        RECT 1724.700 17.330 1724.840 1220.190 ;
        RECT 1724.640 17.010 1724.900 17.330 ;
        RECT 1893.920 17.010 1894.180 17.330 ;
        RECT 1893.980 2.400 1894.120 17.010 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1750.905 1214.225 1751.995 1214.395 ;
      LAYER mcon ;
        RECT 1751.825 1214.225 1751.995 1214.395 ;
      LAYER met1 ;
        RECT 1731.510 1214.380 1731.830 1214.440 ;
        RECT 1750.845 1214.380 1751.135 1214.425 ;
        RECT 1731.510 1214.240 1751.135 1214.380 ;
        RECT 1731.510 1214.180 1731.830 1214.240 ;
        RECT 1750.845 1214.195 1751.135 1214.240 ;
        RECT 1751.765 1214.380 1752.055 1214.425 ;
        RECT 1886.990 1214.380 1887.310 1214.440 ;
        RECT 1751.765 1214.240 1887.310 1214.380 ;
        RECT 1751.765 1214.195 1752.055 1214.240 ;
        RECT 1886.990 1214.180 1887.310 1214.240 ;
        RECT 1886.990 15.540 1887.310 15.600 ;
        RECT 1911.830 15.540 1912.150 15.600 ;
        RECT 1886.990 15.400 1912.150 15.540 ;
        RECT 1886.990 15.340 1887.310 15.400 ;
        RECT 1911.830 15.340 1912.150 15.400 ;
      LAYER via ;
        RECT 1731.540 1214.180 1731.800 1214.440 ;
        RECT 1887.020 1214.180 1887.280 1214.440 ;
        RECT 1887.020 15.340 1887.280 15.600 ;
        RECT 1911.860 15.340 1912.120 15.600 ;
      LAYER met2 ;
        RECT 1731.550 1219.680 1732.110 1228.680 ;
        RECT 1731.600 1214.470 1731.740 1219.680 ;
        RECT 1731.540 1214.150 1731.800 1214.470 ;
        RECT 1887.020 1214.150 1887.280 1214.470 ;
        RECT 1887.080 15.630 1887.220 1214.150 ;
        RECT 1887.020 15.310 1887.280 15.630 ;
        RECT 1911.860 15.310 1912.120 15.630 ;
        RECT 1911.920 2.400 1912.060 15.310 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1740.710 1207.580 1741.030 1207.640 ;
        RECT 1745.310 1207.580 1745.630 1207.640 ;
        RECT 1740.710 1207.440 1745.630 1207.580 ;
        RECT 1740.710 1207.380 1741.030 1207.440 ;
        RECT 1745.310 1207.380 1745.630 1207.440 ;
        RECT 1745.310 20.300 1745.630 20.360 ;
        RECT 1929.310 20.300 1929.630 20.360 ;
        RECT 1745.310 20.160 1929.630 20.300 ;
        RECT 1745.310 20.100 1745.630 20.160 ;
        RECT 1929.310 20.100 1929.630 20.160 ;
      LAYER via ;
        RECT 1740.740 1207.380 1741.000 1207.640 ;
        RECT 1745.340 1207.380 1745.600 1207.640 ;
        RECT 1745.340 20.100 1745.600 20.360 ;
        RECT 1929.340 20.100 1929.600 20.360 ;
      LAYER met2 ;
        RECT 1740.750 1219.680 1741.310 1228.680 ;
        RECT 1740.800 1207.670 1740.940 1219.680 ;
        RECT 1740.740 1207.350 1741.000 1207.670 ;
        RECT 1745.340 1207.350 1745.600 1207.670 ;
        RECT 1745.400 20.390 1745.540 1207.350 ;
        RECT 1745.340 20.070 1745.600 20.390 ;
        RECT 1929.340 20.070 1929.600 20.390 ;
        RECT 1929.400 2.400 1929.540 20.070 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1776.205 1209.465 1776.375 1212.355 ;
      LAYER mcon ;
        RECT 1776.205 1212.185 1776.375 1212.355 ;
      LAYER met1 ;
        RECT 1749.910 1212.340 1750.230 1212.400 ;
        RECT 1776.145 1212.340 1776.435 1212.385 ;
        RECT 1749.910 1212.200 1776.435 1212.340 ;
        RECT 1749.910 1212.140 1750.230 1212.200 ;
        RECT 1776.145 1212.155 1776.435 1212.200 ;
        RECT 1776.145 1209.620 1776.435 1209.665 ;
        RECT 1900.790 1209.620 1901.110 1209.680 ;
        RECT 1776.145 1209.480 1901.110 1209.620 ;
        RECT 1776.145 1209.435 1776.435 1209.480 ;
        RECT 1900.790 1209.420 1901.110 1209.480 ;
        RECT 1900.790 16.560 1901.110 16.620 ;
        RECT 1947.250 16.560 1947.570 16.620 ;
        RECT 1900.790 16.420 1947.570 16.560 ;
        RECT 1900.790 16.360 1901.110 16.420 ;
        RECT 1947.250 16.360 1947.570 16.420 ;
      LAYER via ;
        RECT 1749.940 1212.140 1750.200 1212.400 ;
        RECT 1900.820 1209.420 1901.080 1209.680 ;
        RECT 1900.820 16.360 1901.080 16.620 ;
        RECT 1947.280 16.360 1947.540 16.620 ;
      LAYER met2 ;
        RECT 1749.950 1219.680 1750.510 1228.680 ;
        RECT 1750.000 1212.430 1750.140 1219.680 ;
        RECT 1749.940 1212.110 1750.200 1212.430 ;
        RECT 1900.820 1209.390 1901.080 1209.710 ;
        RECT 1900.880 16.650 1901.020 1209.390 ;
        RECT 1900.820 16.330 1901.080 16.650 ;
        RECT 1947.280 16.330 1947.540 16.650 ;
        RECT 1947.340 2.400 1947.480 16.330 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 1213.360 1759.430 1213.420 ;
        RECT 1835.470 1213.360 1835.790 1213.420 ;
        RECT 1759.110 1213.220 1835.790 1213.360 ;
        RECT 1759.110 1213.160 1759.430 1213.220 ;
        RECT 1835.470 1213.160 1835.790 1213.220 ;
        RECT 1871.350 1210.640 1871.670 1210.700 ;
        RECT 1921.490 1210.640 1921.810 1210.700 ;
        RECT 1871.350 1210.500 1921.810 1210.640 ;
        RECT 1871.350 1210.440 1871.670 1210.500 ;
        RECT 1921.490 1210.440 1921.810 1210.500 ;
        RECT 1921.490 15.880 1921.810 15.940 ;
        RECT 1965.190 15.880 1965.510 15.940 ;
        RECT 1921.490 15.740 1965.510 15.880 ;
        RECT 1921.490 15.680 1921.810 15.740 ;
        RECT 1965.190 15.680 1965.510 15.740 ;
      LAYER via ;
        RECT 1759.140 1213.160 1759.400 1213.420 ;
        RECT 1835.500 1213.160 1835.760 1213.420 ;
        RECT 1871.380 1210.440 1871.640 1210.700 ;
        RECT 1921.520 1210.440 1921.780 1210.700 ;
        RECT 1921.520 15.680 1921.780 15.940 ;
        RECT 1965.220 15.680 1965.480 15.940 ;
      LAYER met2 ;
        RECT 1759.150 1219.680 1759.710 1228.680 ;
        RECT 1759.200 1213.450 1759.340 1219.680 ;
        RECT 1759.140 1213.130 1759.400 1213.450 ;
        RECT 1835.490 1213.275 1835.770 1213.645 ;
        RECT 1871.370 1213.275 1871.650 1213.645 ;
        RECT 1835.500 1213.130 1835.760 1213.275 ;
        RECT 1871.440 1210.730 1871.580 1213.275 ;
        RECT 1871.380 1210.410 1871.640 1210.730 ;
        RECT 1921.520 1210.410 1921.780 1210.730 ;
        RECT 1921.580 15.970 1921.720 1210.410 ;
        RECT 1921.520 15.650 1921.780 15.970 ;
        RECT 1965.220 15.650 1965.480 15.970 ;
        RECT 1965.280 2.400 1965.420 15.650 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 1835.490 1213.320 1835.770 1213.600 ;
        RECT 1871.370 1213.320 1871.650 1213.600 ;
      LAYER met3 ;
        RECT 1835.465 1213.610 1835.795 1213.625 ;
        RECT 1871.345 1213.610 1871.675 1213.625 ;
        RECT 1835.465 1213.310 1871.675 1213.610 ;
        RECT 1835.465 1213.295 1835.795 1213.310 ;
        RECT 1871.345 1213.295 1871.675 1213.310 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1942.190 15.200 1942.510 15.260 ;
        RECT 1983.130 15.200 1983.450 15.260 ;
        RECT 1942.190 15.060 1983.450 15.200 ;
        RECT 1942.190 15.000 1942.510 15.060 ;
        RECT 1983.130 15.000 1983.450 15.060 ;
      LAYER via ;
        RECT 1942.220 15.000 1942.480 15.260 ;
        RECT 1983.160 15.000 1983.420 15.260 ;
      LAYER met2 ;
        RECT 1768.350 1219.680 1768.910 1228.680 ;
        RECT 1768.400 1210.925 1768.540 1219.680 ;
        RECT 1768.330 1210.555 1768.610 1210.925 ;
        RECT 1942.210 1210.555 1942.490 1210.925 ;
        RECT 1942.280 15.290 1942.420 1210.555 ;
        RECT 1942.220 14.970 1942.480 15.290 ;
        RECT 1983.160 14.970 1983.420 15.290 ;
        RECT 1983.220 2.400 1983.360 14.970 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1210.600 1768.610 1210.880 ;
        RECT 1942.210 1210.600 1942.490 1210.880 ;
      LAYER met3 ;
        RECT 1768.305 1210.890 1768.635 1210.905 ;
        RECT 1942.185 1210.890 1942.515 1210.905 ;
        RECT 1768.305 1210.590 1942.515 1210.890 ;
        RECT 1768.305 1210.575 1768.635 1210.590 ;
        RECT 1942.185 1210.575 1942.515 1210.590 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1779.810 19.960 1780.130 20.020 ;
        RECT 2001.070 19.960 2001.390 20.020 ;
        RECT 1779.810 19.820 2001.390 19.960 ;
        RECT 1779.810 19.760 1780.130 19.820 ;
        RECT 2001.070 19.760 2001.390 19.820 ;
      LAYER via ;
        RECT 1779.840 19.760 1780.100 20.020 ;
        RECT 2001.100 19.760 2001.360 20.020 ;
      LAYER met2 ;
        RECT 1777.550 1220.330 1778.110 1228.680 ;
        RECT 1777.550 1220.190 1780.040 1220.330 ;
        RECT 1777.550 1219.680 1778.110 1220.190 ;
        RECT 1779.900 20.050 1780.040 1220.190 ;
        RECT 1779.840 19.730 1780.100 20.050 ;
        RECT 2001.100 19.730 2001.360 20.050 ;
        RECT 2001.160 2.400 2001.300 19.730 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 1212.680 1787.030 1212.740 ;
        RECT 1835.470 1212.680 1835.790 1212.740 ;
        RECT 1786.710 1212.540 1835.790 1212.680 ;
        RECT 1786.710 1212.480 1787.030 1212.540 ;
        RECT 1835.470 1212.480 1835.790 1212.540 ;
        RECT 1837.310 1212.680 1837.630 1212.740 ;
        RECT 1955.990 1212.680 1956.310 1212.740 ;
        RECT 1837.310 1212.540 1956.310 1212.680 ;
        RECT 1837.310 1212.480 1837.630 1212.540 ;
        RECT 1955.990 1212.480 1956.310 1212.540 ;
        RECT 1955.990 16.900 1956.310 16.960 ;
        RECT 2018.550 16.900 2018.870 16.960 ;
        RECT 1955.990 16.760 2018.870 16.900 ;
        RECT 1955.990 16.700 1956.310 16.760 ;
        RECT 2018.550 16.700 2018.870 16.760 ;
      LAYER via ;
        RECT 1786.740 1212.480 1787.000 1212.740 ;
        RECT 1835.500 1212.480 1835.760 1212.740 ;
        RECT 1837.340 1212.480 1837.600 1212.740 ;
        RECT 1956.020 1212.480 1956.280 1212.740 ;
        RECT 1956.020 16.700 1956.280 16.960 ;
        RECT 2018.580 16.700 2018.840 16.960 ;
      LAYER met2 ;
        RECT 1786.750 1219.680 1787.310 1228.680 ;
        RECT 1786.800 1212.770 1786.940 1219.680 ;
        RECT 1786.740 1212.450 1787.000 1212.770 ;
        RECT 1835.490 1212.595 1835.770 1212.965 ;
        RECT 1837.330 1212.595 1837.610 1212.965 ;
        RECT 1835.500 1212.450 1835.760 1212.595 ;
        RECT 1837.340 1212.450 1837.600 1212.595 ;
        RECT 1956.020 1212.450 1956.280 1212.770 ;
        RECT 1956.080 16.990 1956.220 1212.450 ;
        RECT 1956.020 16.670 1956.280 16.990 ;
        RECT 2018.580 16.670 2018.840 16.990 ;
        RECT 2018.640 2.400 2018.780 16.670 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
      LAYER via2 ;
        RECT 1835.490 1212.640 1835.770 1212.920 ;
        RECT 1837.330 1212.640 1837.610 1212.920 ;
      LAYER met3 ;
        RECT 1835.465 1212.930 1835.795 1212.945 ;
        RECT 1837.305 1212.930 1837.635 1212.945 ;
        RECT 1835.465 1212.630 1837.635 1212.930 ;
        RECT 1835.465 1212.615 1835.795 1212.630 ;
        RECT 1837.305 1212.615 1837.635 1212.630 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1795.910 1207.580 1796.230 1207.640 ;
        RECT 1800.510 1207.580 1800.830 1207.640 ;
        RECT 1795.910 1207.440 1800.830 1207.580 ;
        RECT 1795.910 1207.380 1796.230 1207.440 ;
        RECT 1800.510 1207.380 1800.830 1207.440 ;
        RECT 1800.510 19.620 1800.830 19.680 ;
        RECT 2036.490 19.620 2036.810 19.680 ;
        RECT 1800.510 19.480 2036.810 19.620 ;
        RECT 1800.510 19.420 1800.830 19.480 ;
        RECT 2036.490 19.420 2036.810 19.480 ;
      LAYER via ;
        RECT 1795.940 1207.380 1796.200 1207.640 ;
        RECT 1800.540 1207.380 1800.800 1207.640 ;
        RECT 1800.540 19.420 1800.800 19.680 ;
        RECT 2036.520 19.420 2036.780 19.680 ;
      LAYER met2 ;
        RECT 1795.950 1219.680 1796.510 1228.680 ;
        RECT 1796.000 1207.670 1796.140 1219.680 ;
        RECT 1795.940 1207.350 1796.200 1207.670 ;
        RECT 1800.540 1207.350 1800.800 1207.670 ;
        RECT 1800.600 19.710 1800.740 1207.350 ;
        RECT 1800.540 19.390 1800.800 19.710 ;
        RECT 2036.520 19.390 2036.780 19.710 ;
        RECT 2036.580 2.400 2036.720 19.390 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1846.125 1211.505 1846.295 1212.355 ;
      LAYER mcon ;
        RECT 1846.125 1212.185 1846.295 1212.355 ;
      LAYER met1 ;
        RECT 1846.065 1212.340 1846.355 1212.385 ;
        RECT 1976.690 1212.340 1977.010 1212.400 ;
        RECT 1846.065 1212.200 1977.010 1212.340 ;
        RECT 1846.065 1212.155 1846.355 1212.200 ;
        RECT 1976.690 1212.140 1977.010 1212.200 ;
        RECT 1805.110 1211.660 1805.430 1211.720 ;
        RECT 1846.065 1211.660 1846.355 1211.705 ;
        RECT 1805.110 1211.520 1846.355 1211.660 ;
        RECT 1805.110 1211.460 1805.430 1211.520 ;
        RECT 1846.065 1211.475 1846.355 1211.520 ;
        RECT 1976.230 20.300 1976.550 20.360 ;
        RECT 2054.430 20.300 2054.750 20.360 ;
        RECT 1976.230 20.160 2054.750 20.300 ;
        RECT 1976.230 20.100 1976.550 20.160 ;
        RECT 2054.430 20.100 2054.750 20.160 ;
      LAYER via ;
        RECT 1976.720 1212.140 1976.980 1212.400 ;
        RECT 1805.140 1211.460 1805.400 1211.720 ;
        RECT 1976.260 20.100 1976.520 20.360 ;
        RECT 2054.460 20.100 2054.720 20.360 ;
      LAYER met2 ;
        RECT 1805.150 1219.680 1805.710 1228.680 ;
        RECT 1805.200 1211.750 1805.340 1219.680 ;
        RECT 1976.720 1212.110 1976.980 1212.430 ;
        RECT 1805.140 1211.430 1805.400 1211.750 ;
        RECT 1976.780 41.210 1976.920 1212.110 ;
        RECT 1976.320 41.070 1976.920 41.210 ;
        RECT 1976.320 20.390 1976.460 41.070 ;
        RECT 1976.260 20.070 1976.520 20.390 ;
        RECT 2054.460 20.070 2054.720 20.390 ;
        RECT 2054.520 2.400 2054.660 20.070 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1139.030 1196.700 1139.350 1196.760 ;
        RECT 1143.630 1196.700 1143.950 1196.760 ;
        RECT 1139.030 1196.560 1143.950 1196.700 ;
        RECT 1139.030 1196.500 1139.350 1196.560 ;
        RECT 1143.630 1196.500 1143.950 1196.560 ;
        RECT 769.650 30.840 769.970 30.900 ;
        RECT 1139.030 30.840 1139.350 30.900 ;
        RECT 769.650 30.700 1139.350 30.840 ;
        RECT 769.650 30.640 769.970 30.700 ;
        RECT 1139.030 30.640 1139.350 30.700 ;
      LAYER via ;
        RECT 1139.060 1196.500 1139.320 1196.760 ;
        RECT 1143.660 1196.500 1143.920 1196.760 ;
        RECT 769.680 30.640 769.940 30.900 ;
        RECT 1139.060 30.640 1139.320 30.900 ;
      LAYER met2 ;
        RECT 1145.050 1220.330 1145.610 1228.680 ;
        RECT 1143.720 1220.190 1145.610 1220.330 ;
        RECT 1143.720 1196.790 1143.860 1220.190 ;
        RECT 1145.050 1219.680 1145.610 1220.190 ;
        RECT 1139.060 1196.470 1139.320 1196.790 ;
        RECT 1143.660 1196.470 1143.920 1196.790 ;
        RECT 1139.120 30.930 1139.260 1196.470 ;
        RECT 769.680 30.610 769.940 30.930 ;
        RECT 1139.060 30.610 1139.320 30.930 ;
        RECT 769.740 2.400 769.880 30.610 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 19.280 1814.630 19.340 ;
        RECT 2072.370 19.280 2072.690 19.340 ;
        RECT 1814.310 19.140 2072.690 19.280 ;
        RECT 1814.310 19.080 1814.630 19.140 ;
        RECT 2072.370 19.080 2072.690 19.140 ;
      LAYER via ;
        RECT 1814.340 19.080 1814.600 19.340 ;
        RECT 2072.400 19.080 2072.660 19.340 ;
      LAYER met2 ;
        RECT 1814.350 1219.680 1814.910 1228.680 ;
        RECT 1814.400 19.370 1814.540 1219.680 ;
        RECT 1814.340 19.050 1814.600 19.370 ;
        RECT 2072.400 19.050 2072.660 19.370 ;
        RECT 2072.460 2.400 2072.600 19.050 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1850.265 1211.505 1850.435 1214.055 ;
      LAYER mcon ;
        RECT 1850.265 1213.885 1850.435 1214.055 ;
      LAYER met1 ;
        RECT 1823.510 1214.040 1823.830 1214.100 ;
        RECT 1850.205 1214.040 1850.495 1214.085 ;
        RECT 1823.510 1213.900 1850.495 1214.040 ;
        RECT 1823.510 1213.840 1823.830 1213.900 ;
        RECT 1850.205 1213.855 1850.495 1213.900 ;
        RECT 1850.205 1211.660 1850.495 1211.705 ;
        RECT 2045.690 1211.660 2046.010 1211.720 ;
        RECT 1850.205 1211.520 2046.010 1211.660 ;
        RECT 1850.205 1211.475 1850.495 1211.520 ;
        RECT 2045.690 1211.460 2046.010 1211.520 ;
        RECT 2045.690 19.620 2046.010 19.680 ;
        RECT 2089.850 19.620 2090.170 19.680 ;
        RECT 2045.690 19.480 2090.170 19.620 ;
        RECT 2045.690 19.420 2046.010 19.480 ;
        RECT 2089.850 19.420 2090.170 19.480 ;
      LAYER via ;
        RECT 1823.540 1213.840 1823.800 1214.100 ;
        RECT 2045.720 1211.460 2045.980 1211.720 ;
        RECT 2045.720 19.420 2045.980 19.680 ;
        RECT 2089.880 19.420 2090.140 19.680 ;
      LAYER met2 ;
        RECT 1823.550 1219.680 1824.110 1228.680 ;
        RECT 1823.600 1214.130 1823.740 1219.680 ;
        RECT 1823.540 1213.810 1823.800 1214.130 ;
        RECT 2045.720 1211.430 2045.980 1211.750 ;
        RECT 2045.780 19.710 2045.920 1211.430 ;
        RECT 2045.720 19.390 2045.980 19.710 ;
        RECT 2089.880 19.390 2090.140 19.710 ;
        RECT 2089.940 2.400 2090.080 19.390 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1834.550 18.600 1834.870 18.660 ;
        RECT 2107.790 18.600 2108.110 18.660 ;
        RECT 1834.550 18.460 2108.110 18.600 ;
        RECT 1834.550 18.400 1834.870 18.460 ;
        RECT 2107.790 18.400 2108.110 18.460 ;
      LAYER via ;
        RECT 1834.580 18.400 1834.840 18.660 ;
        RECT 2107.820 18.400 2108.080 18.660 ;
      LAYER met2 ;
        RECT 1832.750 1220.330 1833.310 1228.680 ;
        RECT 1832.750 1220.190 1834.780 1220.330 ;
        RECT 1832.750 1219.680 1833.310 1220.190 ;
        RECT 1834.640 18.690 1834.780 1220.190 ;
        RECT 1834.580 18.370 1834.840 18.690 ;
        RECT 2107.820 18.370 2108.080 18.690 ;
        RECT 2107.880 2.400 2108.020 18.370 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1841.910 1211.320 1842.230 1211.380 ;
        RECT 2056.270 1211.320 2056.590 1211.380 ;
        RECT 1841.910 1211.180 2056.590 1211.320 ;
        RECT 1841.910 1211.120 1842.230 1211.180 ;
        RECT 2056.270 1211.120 2056.590 1211.180 ;
        RECT 2056.270 1207.580 2056.590 1207.640 ;
        RECT 2059.490 1207.580 2059.810 1207.640 ;
        RECT 2056.270 1207.440 2059.810 1207.580 ;
        RECT 2056.270 1207.380 2056.590 1207.440 ;
        RECT 2059.490 1207.380 2059.810 1207.440 ;
        RECT 2059.490 15.200 2059.810 15.260 ;
        RECT 2125.730 15.200 2126.050 15.260 ;
        RECT 2059.490 15.060 2126.050 15.200 ;
        RECT 2059.490 15.000 2059.810 15.060 ;
        RECT 2125.730 15.000 2126.050 15.060 ;
      LAYER via ;
        RECT 1841.940 1211.120 1842.200 1211.380 ;
        RECT 2056.300 1211.120 2056.560 1211.380 ;
        RECT 2056.300 1207.380 2056.560 1207.640 ;
        RECT 2059.520 1207.380 2059.780 1207.640 ;
        RECT 2059.520 15.000 2059.780 15.260 ;
        RECT 2125.760 15.000 2126.020 15.260 ;
      LAYER met2 ;
        RECT 1841.950 1219.680 1842.510 1228.680 ;
        RECT 1842.000 1211.410 1842.140 1219.680 ;
        RECT 1841.940 1211.090 1842.200 1211.410 ;
        RECT 2056.300 1211.090 2056.560 1211.410 ;
        RECT 2056.360 1207.670 2056.500 1211.090 ;
        RECT 2056.300 1207.350 2056.560 1207.670 ;
        RECT 2059.520 1207.350 2059.780 1207.670 ;
        RECT 2059.580 15.290 2059.720 1207.350 ;
        RECT 2059.520 14.970 2059.780 15.290 ;
        RECT 2125.760 14.970 2126.020 15.290 ;
        RECT 2125.820 2.400 2125.960 14.970 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1850.650 1214.040 1850.970 1214.100 ;
        RECT 1855.710 1214.040 1856.030 1214.100 ;
        RECT 1850.650 1213.900 1856.030 1214.040 ;
        RECT 1850.650 1213.840 1850.970 1213.900 ;
        RECT 1855.710 1213.840 1856.030 1213.900 ;
        RECT 1855.710 18.260 1856.030 18.320 ;
        RECT 2143.670 18.260 2143.990 18.320 ;
        RECT 1855.710 18.120 2143.990 18.260 ;
        RECT 1855.710 18.060 1856.030 18.120 ;
        RECT 2143.670 18.060 2143.990 18.120 ;
      LAYER via ;
        RECT 1850.680 1213.840 1850.940 1214.100 ;
        RECT 1855.740 1213.840 1856.000 1214.100 ;
        RECT 1855.740 18.060 1856.000 18.320 ;
        RECT 2143.700 18.060 2143.960 18.320 ;
      LAYER met2 ;
        RECT 1850.690 1219.680 1851.250 1228.680 ;
        RECT 1850.740 1214.130 1850.880 1219.680 ;
        RECT 1850.680 1213.810 1850.940 1214.130 ;
        RECT 1855.740 1213.810 1856.000 1214.130 ;
        RECT 1855.800 18.350 1855.940 1213.810 ;
        RECT 1855.740 18.030 1856.000 18.350 ;
        RECT 2143.700 18.030 2143.960 18.350 ;
        RECT 2143.760 2.400 2143.900 18.030 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 17.920 1862.930 17.980 ;
        RECT 2161.610 17.920 2161.930 17.980 ;
        RECT 1862.610 17.780 2161.930 17.920 ;
        RECT 1862.610 17.720 1862.930 17.780 ;
        RECT 2161.610 17.720 2161.930 17.780 ;
      LAYER via ;
        RECT 1862.640 17.720 1862.900 17.980 ;
        RECT 2161.640 17.720 2161.900 17.980 ;
      LAYER met2 ;
        RECT 1859.890 1220.330 1860.450 1228.680 ;
        RECT 1859.890 1220.190 1862.840 1220.330 ;
        RECT 1859.890 1219.680 1860.450 1220.190 ;
        RECT 1862.700 18.010 1862.840 1220.190 ;
        RECT 1862.640 17.690 1862.900 18.010 ;
        RECT 2161.640 17.690 2161.900 18.010 ;
        RECT 2161.700 2.400 2161.840 17.690 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.510 17.580 1869.830 17.640 ;
        RECT 2179.090 17.580 2179.410 17.640 ;
        RECT 1869.510 17.440 2179.410 17.580 ;
        RECT 1869.510 17.380 1869.830 17.440 ;
        RECT 2179.090 17.380 2179.410 17.440 ;
      LAYER via ;
        RECT 1869.540 17.380 1869.800 17.640 ;
        RECT 2179.120 17.380 2179.380 17.640 ;
      LAYER met2 ;
        RECT 1869.090 1220.330 1869.650 1228.680 ;
        RECT 1869.090 1219.680 1869.740 1220.330 ;
        RECT 1869.600 17.670 1869.740 1219.680 ;
        RECT 1869.540 17.350 1869.800 17.670 ;
        RECT 2179.120 17.350 2179.380 17.670 ;
        RECT 2179.180 2.400 2179.320 17.350 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1878.250 1214.040 1878.570 1214.100 ;
        RECT 2195.190 1214.040 2195.510 1214.100 ;
        RECT 1878.250 1213.900 2195.510 1214.040 ;
        RECT 1878.250 1213.840 1878.570 1213.900 ;
        RECT 2195.190 1213.840 2195.510 1213.900 ;
        RECT 2195.190 2.960 2195.510 3.020 ;
        RECT 2197.030 2.960 2197.350 3.020 ;
        RECT 2195.190 2.820 2197.350 2.960 ;
        RECT 2195.190 2.760 2195.510 2.820 ;
        RECT 2197.030 2.760 2197.350 2.820 ;
      LAYER via ;
        RECT 1878.280 1213.840 1878.540 1214.100 ;
        RECT 2195.220 1213.840 2195.480 1214.100 ;
        RECT 2195.220 2.760 2195.480 3.020 ;
        RECT 2197.060 2.760 2197.320 3.020 ;
      LAYER met2 ;
        RECT 1878.290 1219.680 1878.850 1228.680 ;
        RECT 1878.340 1214.130 1878.480 1219.680 ;
        RECT 1878.280 1213.810 1878.540 1214.130 ;
        RECT 2195.220 1213.810 2195.480 1214.130 ;
        RECT 2195.280 3.050 2195.420 1213.810 ;
        RECT 2195.220 2.730 2195.480 3.050 ;
        RECT 2197.060 2.730 2197.320 3.050 ;
        RECT 2197.120 2.400 2197.260 2.730 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1887.450 1208.260 1887.770 1208.320 ;
        RECT 1901.250 1208.260 1901.570 1208.320 ;
        RECT 1887.450 1208.120 1901.570 1208.260 ;
        RECT 1887.450 1208.060 1887.770 1208.120 ;
        RECT 1901.250 1208.060 1901.570 1208.120 ;
        RECT 2214.970 17.240 2215.290 17.300 ;
        RECT 1953.780 17.100 2215.290 17.240 ;
        RECT 1901.250 16.220 1901.570 16.280 ;
        RECT 1953.780 16.220 1953.920 17.100 ;
        RECT 2214.970 17.040 2215.290 17.100 ;
        RECT 1901.250 16.080 1953.920 16.220 ;
        RECT 1901.250 16.020 1901.570 16.080 ;
      LAYER via ;
        RECT 1887.480 1208.060 1887.740 1208.320 ;
        RECT 1901.280 1208.060 1901.540 1208.320 ;
        RECT 1901.280 16.020 1901.540 16.280 ;
        RECT 2215.000 17.040 2215.260 17.300 ;
      LAYER met2 ;
        RECT 1887.490 1219.680 1888.050 1228.680 ;
        RECT 1887.540 1208.350 1887.680 1219.680 ;
        RECT 1887.480 1208.030 1887.740 1208.350 ;
        RECT 1901.280 1208.030 1901.540 1208.350 ;
        RECT 1901.340 16.310 1901.480 1208.030 ;
        RECT 2215.000 17.010 2215.260 17.330 ;
        RECT 1901.280 15.990 1901.540 16.310 ;
        RECT 2215.060 2.400 2215.200 17.010 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2213.205 1210.485 2215.675 1210.655 ;
        RECT 2213.205 1210.145 2213.375 1210.485 ;
      LAYER mcon ;
        RECT 2215.505 1210.485 2215.675 1210.655 ;
      LAYER met1 ;
        RECT 2215.445 1210.640 2215.735 1210.685 ;
        RECT 2228.770 1210.640 2229.090 1210.700 ;
        RECT 2215.445 1210.500 2229.090 1210.640 ;
        RECT 2215.445 1210.455 2215.735 1210.500 ;
        RECT 2228.770 1210.440 2229.090 1210.500 ;
        RECT 1896.650 1210.300 1896.970 1210.360 ;
        RECT 2213.145 1210.300 2213.435 1210.345 ;
        RECT 1896.650 1210.160 2213.435 1210.300 ;
        RECT 1896.650 1210.100 1896.970 1210.160 ;
        RECT 2213.145 1210.115 2213.435 1210.160 ;
        RECT 2228.770 2.960 2229.090 3.020 ;
        RECT 2232.910 2.960 2233.230 3.020 ;
        RECT 2228.770 2.820 2233.230 2.960 ;
        RECT 2228.770 2.760 2229.090 2.820 ;
        RECT 2232.910 2.760 2233.230 2.820 ;
      LAYER via ;
        RECT 2228.800 1210.440 2229.060 1210.700 ;
        RECT 1896.680 1210.100 1896.940 1210.360 ;
        RECT 2228.800 2.760 2229.060 3.020 ;
        RECT 2232.940 2.760 2233.200 3.020 ;
      LAYER met2 ;
        RECT 1896.690 1219.680 1897.250 1228.680 ;
        RECT 1896.740 1210.390 1896.880 1219.680 ;
        RECT 2228.800 1210.410 2229.060 1210.730 ;
        RECT 1896.680 1210.070 1896.940 1210.390 ;
        RECT 2228.860 3.050 2229.000 1210.410 ;
        RECT 2228.800 2.730 2229.060 3.050 ;
        RECT 2232.940 2.730 2233.200 3.050 ;
        RECT 2233.000 2.400 2233.140 2.730 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 787.590 31.180 787.910 31.240 ;
        RECT 1152.830 31.180 1153.150 31.240 ;
        RECT 787.590 31.040 1153.150 31.180 ;
        RECT 787.590 30.980 787.910 31.040 ;
        RECT 1152.830 30.980 1153.150 31.040 ;
      LAYER via ;
        RECT 787.620 30.980 787.880 31.240 ;
        RECT 1152.860 30.980 1153.120 31.240 ;
      LAYER met2 ;
        RECT 1154.250 1220.330 1154.810 1228.680 ;
        RECT 1152.920 1220.190 1154.810 1220.330 ;
        RECT 1152.920 31.270 1153.060 1220.190 ;
        RECT 1154.250 1219.680 1154.810 1220.190 ;
        RECT 787.620 30.950 787.880 31.270 ;
        RECT 1152.860 30.950 1153.120 31.270 ;
        RECT 787.680 2.400 787.820 30.950 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1932.145 13.685 1932.315 14.875 ;
        RECT 1979.985 13.685 1980.155 14.535 ;
      LAYER mcon ;
        RECT 1932.145 14.705 1932.315 14.875 ;
        RECT 1979.985 14.365 1980.155 14.535 ;
      LAYER met1 ;
        RECT 1905.850 1207.920 1906.170 1207.980 ;
        RECT 1921.950 1207.920 1922.270 1207.980 ;
        RECT 1905.850 1207.780 1922.270 1207.920 ;
        RECT 1905.850 1207.720 1906.170 1207.780 ;
        RECT 1921.950 1207.720 1922.270 1207.780 ;
        RECT 1921.950 620.540 1922.270 620.800 ;
        RECT 1922.040 619.780 1922.180 620.540 ;
        RECT 1921.950 619.520 1922.270 619.780 ;
        RECT 2250.850 15.540 2251.170 15.600 ;
        RECT 1983.680 15.400 2251.170 15.540 ;
        RECT 1921.950 14.860 1922.270 14.920 ;
        RECT 1932.085 14.860 1932.375 14.905 ;
        RECT 1921.950 14.720 1932.375 14.860 ;
        RECT 1921.950 14.660 1922.270 14.720 ;
        RECT 1932.085 14.675 1932.375 14.720 ;
        RECT 1979.925 14.520 1980.215 14.565 ;
        RECT 1983.680 14.520 1983.820 15.400 ;
        RECT 2250.850 15.340 2251.170 15.400 ;
        RECT 1979.925 14.380 1983.820 14.520 ;
        RECT 1979.925 14.335 1980.215 14.380 ;
        RECT 1932.085 13.840 1932.375 13.885 ;
        RECT 1979.925 13.840 1980.215 13.885 ;
        RECT 1932.085 13.700 1980.215 13.840 ;
        RECT 1932.085 13.655 1932.375 13.700 ;
        RECT 1979.925 13.655 1980.215 13.700 ;
      LAYER via ;
        RECT 1905.880 1207.720 1906.140 1207.980 ;
        RECT 1921.980 1207.720 1922.240 1207.980 ;
        RECT 1921.980 620.540 1922.240 620.800 ;
        RECT 1921.980 619.520 1922.240 619.780 ;
        RECT 1921.980 14.660 1922.240 14.920 ;
        RECT 2250.880 15.340 2251.140 15.600 ;
      LAYER met2 ;
        RECT 1905.890 1219.680 1906.450 1228.680 ;
        RECT 1905.940 1208.010 1906.080 1219.680 ;
        RECT 1905.880 1207.690 1906.140 1208.010 ;
        RECT 1921.980 1207.690 1922.240 1208.010 ;
        RECT 1922.040 620.830 1922.180 1207.690 ;
        RECT 1921.980 620.510 1922.240 620.830 ;
        RECT 1921.980 619.490 1922.240 619.810 ;
        RECT 1922.040 14.950 1922.180 619.490 ;
        RECT 2250.880 15.310 2251.140 15.630 ;
        RECT 1921.980 14.630 1922.240 14.950 ;
        RECT 2250.940 2.400 2251.080 15.310 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1915.050 1208.260 1915.370 1208.320 ;
        RECT 1915.050 1208.120 1943.340 1208.260 ;
        RECT 1915.050 1208.060 1915.370 1208.120 ;
        RECT 1943.200 1207.920 1943.340 1208.120 ;
        RECT 2263.270 1207.920 2263.590 1207.980 ;
        RECT 1943.200 1207.780 2263.590 1207.920 ;
        RECT 2263.270 1207.720 2263.590 1207.780 ;
      LAYER via ;
        RECT 1915.080 1208.060 1915.340 1208.320 ;
        RECT 2263.300 1207.720 2263.560 1207.980 ;
      LAYER met2 ;
        RECT 1915.090 1219.680 1915.650 1228.680 ;
        RECT 1915.140 1208.350 1915.280 1219.680 ;
        RECT 1915.080 1208.030 1915.340 1208.350 ;
        RECT 2263.300 1207.690 2263.560 1208.010 ;
        RECT 2263.360 16.730 2263.500 1207.690 ;
        RECT 2263.360 16.590 2268.560 16.730 ;
        RECT 2268.420 2.400 2268.560 16.590 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1969.865 1208.105 1970.035 1210.655 ;
      LAYER mcon ;
        RECT 1969.865 1210.485 1970.035 1210.655 ;
      LAYER met1 ;
        RECT 1924.250 1210.640 1924.570 1210.700 ;
        RECT 1969.805 1210.640 1970.095 1210.685 ;
        RECT 1924.250 1210.500 1970.095 1210.640 ;
        RECT 1924.250 1210.440 1924.570 1210.500 ;
        RECT 1969.805 1210.455 1970.095 1210.500 ;
        RECT 1969.805 1208.260 1970.095 1208.305 ;
        RECT 2283.970 1208.260 2284.290 1208.320 ;
        RECT 1969.805 1208.120 2284.290 1208.260 ;
        RECT 1969.805 1208.075 1970.095 1208.120 ;
        RECT 2283.970 1208.060 2284.290 1208.120 ;
      LAYER via ;
        RECT 1924.280 1210.440 1924.540 1210.700 ;
        RECT 2284.000 1208.060 2284.260 1208.320 ;
      LAYER met2 ;
        RECT 1924.290 1219.680 1924.850 1228.680 ;
        RECT 1924.340 1210.730 1924.480 1219.680 ;
        RECT 1924.280 1210.410 1924.540 1210.730 ;
        RECT 2284.000 1208.030 2284.260 1208.350 ;
        RECT 2284.060 16.730 2284.200 1208.030 ;
        RECT 2284.060 16.590 2286.500 16.730 ;
        RECT 2286.360 2.400 2286.500 16.590 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1933.450 1207.920 1933.770 1207.980 ;
        RECT 1942.650 1207.920 1942.970 1207.980 ;
        RECT 1933.450 1207.780 1942.970 1207.920 ;
        RECT 1933.450 1207.720 1933.770 1207.780 ;
        RECT 1942.650 1207.720 1942.970 1207.780 ;
        RECT 2304.210 15.880 2304.530 15.940 ;
        RECT 1969.880 15.740 2304.530 15.880 ;
        RECT 1942.650 15.540 1942.970 15.600 ;
        RECT 1969.880 15.540 1970.020 15.740 ;
        RECT 2304.210 15.680 2304.530 15.740 ;
        RECT 1942.650 15.400 1970.020 15.540 ;
        RECT 1942.650 15.340 1942.970 15.400 ;
      LAYER via ;
        RECT 1933.480 1207.720 1933.740 1207.980 ;
        RECT 1942.680 1207.720 1942.940 1207.980 ;
        RECT 1942.680 15.340 1942.940 15.600 ;
        RECT 2304.240 15.680 2304.500 15.940 ;
      LAYER met2 ;
        RECT 1933.490 1219.680 1934.050 1228.680 ;
        RECT 1933.540 1208.010 1933.680 1219.680 ;
        RECT 1933.480 1207.690 1933.740 1208.010 ;
        RECT 1942.680 1207.690 1942.940 1208.010 ;
        RECT 1942.740 15.630 1942.880 1207.690 ;
        RECT 2304.240 15.650 2304.500 15.970 ;
        RECT 1942.680 15.310 1942.940 15.630 ;
        RECT 2304.300 2.400 2304.440 15.650 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1942.650 1209.280 1942.970 1209.340 ;
        RECT 1942.650 1209.140 1969.560 1209.280 ;
        RECT 1942.650 1209.080 1942.970 1209.140 ;
        RECT 1969.420 1208.600 1969.560 1209.140 ;
        RECT 2318.470 1208.600 2318.790 1208.660 ;
        RECT 1969.420 1208.460 2318.790 1208.600 ;
        RECT 2318.470 1208.400 2318.790 1208.460 ;
      LAYER via ;
        RECT 1942.680 1209.080 1942.940 1209.340 ;
        RECT 2318.500 1208.400 2318.760 1208.660 ;
      LAYER met2 ;
        RECT 1942.690 1219.680 1943.250 1228.680 ;
        RECT 1942.740 1209.370 1942.880 1219.680 ;
        RECT 1942.680 1209.050 1942.940 1209.370 ;
        RECT 2318.500 1208.370 2318.760 1208.690 ;
        RECT 2318.560 16.730 2318.700 1208.370 ;
        RECT 2318.560 16.590 2322.380 16.730 ;
        RECT 2322.240 2.400 2322.380 16.590 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1951.850 1208.260 1952.170 1208.320 ;
        RECT 1962.890 1208.260 1963.210 1208.320 ;
        RECT 1951.850 1208.120 1963.210 1208.260 ;
        RECT 1951.850 1208.060 1952.170 1208.120 ;
        RECT 1962.890 1208.060 1963.210 1208.120 ;
        RECT 1962.890 16.560 1963.210 16.620 ;
        RECT 1962.890 16.420 1970.480 16.560 ;
        RECT 1962.890 16.360 1963.210 16.420 ;
        RECT 1970.340 16.220 1970.480 16.420 ;
        RECT 2339.630 16.220 2339.950 16.280 ;
        RECT 1970.340 16.080 2339.950 16.220 ;
        RECT 2339.630 16.020 2339.950 16.080 ;
      LAYER via ;
        RECT 1951.880 1208.060 1952.140 1208.320 ;
        RECT 1962.920 1208.060 1963.180 1208.320 ;
        RECT 1962.920 16.360 1963.180 16.620 ;
        RECT 2339.660 16.020 2339.920 16.280 ;
      LAYER met2 ;
        RECT 1951.890 1219.680 1952.450 1228.680 ;
        RECT 1951.940 1208.350 1952.080 1219.680 ;
        RECT 1951.880 1208.030 1952.140 1208.350 ;
        RECT 1962.920 1208.030 1963.180 1208.350 ;
        RECT 1962.980 16.650 1963.120 1208.030 ;
        RECT 1962.920 16.330 1963.180 16.650 ;
        RECT 2339.660 15.990 2339.920 16.310 ;
        RECT 2339.720 2.400 2339.860 15.990 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1977.685 1209.125 1977.855 1210.995 ;
      LAYER mcon ;
        RECT 1977.685 1210.825 1977.855 1210.995 ;
      LAYER met1 ;
        RECT 1961.050 1210.980 1961.370 1211.040 ;
        RECT 1977.625 1210.980 1977.915 1211.025 ;
        RECT 1961.050 1210.840 1977.915 1210.980 ;
        RECT 1961.050 1210.780 1961.370 1210.840 ;
        RECT 1977.625 1210.795 1977.915 1210.840 ;
        RECT 1977.625 1209.280 1977.915 1209.325 ;
        RECT 2352.970 1209.280 2353.290 1209.340 ;
        RECT 1977.625 1209.140 2353.290 1209.280 ;
        RECT 1977.625 1209.095 1977.915 1209.140 ;
        RECT 2352.970 1209.080 2353.290 1209.140 ;
        RECT 2352.970 2.960 2353.290 3.020 ;
        RECT 2357.570 2.960 2357.890 3.020 ;
        RECT 2352.970 2.820 2357.890 2.960 ;
        RECT 2352.970 2.760 2353.290 2.820 ;
        RECT 2357.570 2.760 2357.890 2.820 ;
      LAYER via ;
        RECT 1961.080 1210.780 1961.340 1211.040 ;
        RECT 2353.000 1209.080 2353.260 1209.340 ;
        RECT 2353.000 2.760 2353.260 3.020 ;
        RECT 2357.600 2.760 2357.860 3.020 ;
      LAYER met2 ;
        RECT 1961.090 1219.680 1961.650 1228.680 ;
        RECT 1961.140 1211.070 1961.280 1219.680 ;
        RECT 1961.080 1210.750 1961.340 1211.070 ;
        RECT 2353.000 1209.050 2353.260 1209.370 ;
        RECT 2353.060 3.050 2353.200 1209.050 ;
        RECT 2353.000 2.730 2353.260 3.050 ;
        RECT 2357.600 2.730 2357.860 3.050 ;
        RECT 2357.660 2.400 2357.800 2.730 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1969.790 1207.580 1970.110 1207.640 ;
        RECT 1977.150 1207.580 1977.470 1207.640 ;
        RECT 1969.790 1207.440 1977.470 1207.580 ;
        RECT 1969.790 1207.380 1970.110 1207.440 ;
        RECT 1977.150 1207.380 1977.470 1207.440 ;
        RECT 1977.150 20.640 1977.470 20.700 ;
        RECT 2375.510 20.640 2375.830 20.700 ;
        RECT 1977.150 20.500 2375.830 20.640 ;
        RECT 1977.150 20.440 1977.470 20.500 ;
        RECT 2375.510 20.440 2375.830 20.500 ;
      LAYER via ;
        RECT 1969.820 1207.380 1970.080 1207.640 ;
        RECT 1977.180 1207.380 1977.440 1207.640 ;
        RECT 1977.180 20.440 1977.440 20.700 ;
        RECT 2375.540 20.440 2375.800 20.700 ;
      LAYER met2 ;
        RECT 1969.830 1219.680 1970.390 1228.680 ;
        RECT 1969.880 1207.670 1970.020 1219.680 ;
        RECT 1969.820 1207.350 1970.080 1207.670 ;
        RECT 1977.180 1207.350 1977.440 1207.670 ;
        RECT 1977.240 20.730 1977.380 1207.350 ;
        RECT 1977.180 20.410 1977.440 20.730 ;
        RECT 2375.540 20.410 2375.800 20.730 ;
        RECT 2375.600 2.400 2375.740 20.410 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1978.990 1209.960 1979.310 1210.020 ;
        RECT 2387.930 1209.960 2388.250 1210.020 ;
        RECT 1978.990 1209.820 2388.250 1209.960 ;
        RECT 1978.990 1209.760 1979.310 1209.820 ;
        RECT 2387.930 1209.760 2388.250 1209.820 ;
        RECT 2387.930 2.960 2388.250 3.020 ;
        RECT 2393.450 2.960 2393.770 3.020 ;
        RECT 2387.930 2.820 2393.770 2.960 ;
        RECT 2387.930 2.760 2388.250 2.820 ;
        RECT 2393.450 2.760 2393.770 2.820 ;
      LAYER via ;
        RECT 1979.020 1209.760 1979.280 1210.020 ;
        RECT 2387.960 1209.760 2388.220 1210.020 ;
        RECT 2387.960 2.760 2388.220 3.020 ;
        RECT 2393.480 2.760 2393.740 3.020 ;
      LAYER met2 ;
        RECT 1979.030 1219.680 1979.590 1228.680 ;
        RECT 1979.080 1210.050 1979.220 1219.680 ;
        RECT 1979.020 1209.730 1979.280 1210.050 ;
        RECT 2387.960 1209.730 2388.220 1210.050 ;
        RECT 2388.020 3.050 2388.160 1209.730 ;
        RECT 2387.960 2.730 2388.220 3.050 ;
        RECT 2393.480 2.730 2393.740 3.050 ;
        RECT 2393.540 2.400 2393.680 2.730 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2017.705 1110.865 2017.875 1158.975 ;
        RECT 2019.085 144.925 2019.255 193.035 ;
      LAYER mcon ;
        RECT 2017.705 1158.805 2017.875 1158.975 ;
        RECT 2019.085 192.865 2019.255 193.035 ;
      LAYER met1 ;
        RECT 1988.190 1212.680 1988.510 1212.740 ;
        RECT 2018.090 1212.680 2018.410 1212.740 ;
        RECT 1988.190 1212.540 2018.410 1212.680 ;
        RECT 1988.190 1212.480 1988.510 1212.540 ;
        RECT 2018.090 1212.480 2018.410 1212.540 ;
        RECT 2018.090 1173.580 2018.410 1173.640 ;
        RECT 2017.720 1173.440 2018.410 1173.580 ;
        RECT 2017.720 1172.960 2017.860 1173.440 ;
        RECT 2018.090 1173.380 2018.410 1173.440 ;
        RECT 2017.630 1172.700 2017.950 1172.960 ;
        RECT 2017.630 1158.960 2017.950 1159.020 ;
        RECT 2017.435 1158.820 2017.950 1158.960 ;
        RECT 2017.630 1158.760 2017.950 1158.820 ;
        RECT 2017.645 1111.020 2017.935 1111.065 ;
        RECT 2018.550 1111.020 2018.870 1111.080 ;
        RECT 2017.645 1110.880 2018.870 1111.020 ;
        RECT 2017.645 1110.835 2017.935 1110.880 ;
        RECT 2018.550 1110.820 2018.870 1110.880 ;
        RECT 2017.630 1076.000 2017.950 1076.060 ;
        RECT 2018.550 1076.000 2018.870 1076.060 ;
        RECT 2017.630 1075.860 2018.870 1076.000 ;
        RECT 2017.630 1075.800 2017.950 1075.860 ;
        RECT 2018.550 1075.800 2018.870 1075.860 ;
        RECT 2017.630 1028.060 2017.950 1028.120 ;
        RECT 2018.550 1028.060 2018.870 1028.120 ;
        RECT 2017.630 1027.920 2018.870 1028.060 ;
        RECT 2017.630 1027.860 2017.950 1027.920 ;
        RECT 2018.550 1027.860 2018.870 1027.920 ;
        RECT 2019.010 966.180 2019.330 966.240 ;
        RECT 2019.930 966.180 2020.250 966.240 ;
        RECT 2019.010 966.040 2020.250 966.180 ;
        RECT 2019.010 965.980 2019.330 966.040 ;
        RECT 2019.930 965.980 2020.250 966.040 ;
        RECT 2019.010 869.620 2019.330 869.680 ;
        RECT 2019.930 869.620 2020.250 869.680 ;
        RECT 2019.010 869.480 2020.250 869.620 ;
        RECT 2019.010 869.420 2019.330 869.480 ;
        RECT 2019.930 869.420 2020.250 869.480 ;
        RECT 2017.630 821.000 2017.950 821.060 ;
        RECT 2018.550 821.000 2018.870 821.060 ;
        RECT 2017.630 820.860 2018.870 821.000 ;
        RECT 2017.630 820.800 2017.950 820.860 ;
        RECT 2018.550 820.800 2018.870 820.860 ;
        RECT 2018.090 690.440 2018.410 690.500 ;
        RECT 2017.720 690.300 2018.410 690.440 ;
        RECT 2017.720 689.820 2017.860 690.300 ;
        RECT 2018.090 690.240 2018.410 690.300 ;
        RECT 2017.630 689.560 2017.950 689.820 ;
        RECT 2016.250 676.160 2016.570 676.220 ;
        RECT 2017.630 676.160 2017.950 676.220 ;
        RECT 2016.250 676.020 2017.950 676.160 ;
        RECT 2016.250 675.960 2016.570 676.020 ;
        RECT 2017.630 675.960 2017.950 676.020 ;
        RECT 2017.170 593.340 2017.490 593.600 ;
        RECT 2017.260 593.200 2017.400 593.340 ;
        RECT 2017.630 593.200 2017.950 593.260 ;
        RECT 2017.260 593.060 2017.950 593.200 ;
        RECT 2017.630 593.000 2017.950 593.060 ;
        RECT 2016.250 579.600 2016.570 579.660 ;
        RECT 2017.630 579.600 2017.950 579.660 ;
        RECT 2016.250 579.460 2017.950 579.600 ;
        RECT 2016.250 579.400 2016.570 579.460 ;
        RECT 2017.630 579.400 2017.950 579.460 ;
        RECT 2017.170 496.780 2017.490 497.040 ;
        RECT 2017.260 496.640 2017.400 496.780 ;
        RECT 2017.630 496.640 2017.950 496.700 ;
        RECT 2017.260 496.500 2017.950 496.640 ;
        RECT 2017.630 496.440 2017.950 496.500 ;
        RECT 2016.250 483.040 2016.570 483.100 ;
        RECT 2017.630 483.040 2017.950 483.100 ;
        RECT 2016.250 482.900 2017.950 483.040 ;
        RECT 2016.250 482.840 2016.570 482.900 ;
        RECT 2017.630 482.840 2017.950 482.900 ;
        RECT 2017.170 400.220 2017.490 400.480 ;
        RECT 2017.260 399.740 2017.400 400.220 ;
        RECT 2017.630 399.740 2017.950 399.800 ;
        RECT 2017.260 399.600 2017.950 399.740 ;
        RECT 2017.630 399.540 2017.950 399.600 ;
        RECT 2017.170 310.660 2017.490 310.720 ;
        RECT 2017.630 310.660 2017.950 310.720 ;
        RECT 2017.170 310.520 2017.950 310.660 ;
        RECT 2017.170 310.460 2017.490 310.520 ;
        RECT 2017.630 310.460 2017.950 310.520 ;
        RECT 2018.090 262.380 2018.410 262.440 ;
        RECT 2018.550 262.380 2018.870 262.440 ;
        RECT 2018.090 262.240 2018.870 262.380 ;
        RECT 2018.090 262.180 2018.410 262.240 ;
        RECT 2018.550 262.180 2018.870 262.240 ;
        RECT 2018.550 241.640 2018.870 241.700 ;
        RECT 2019.010 241.640 2019.330 241.700 ;
        RECT 2018.550 241.500 2019.330 241.640 ;
        RECT 2018.550 241.440 2018.870 241.500 ;
        RECT 2019.010 241.440 2019.330 241.500 ;
        RECT 2019.010 193.020 2019.330 193.080 ;
        RECT 2018.815 192.880 2019.330 193.020 ;
        RECT 2019.010 192.820 2019.330 192.880 ;
        RECT 2019.025 145.080 2019.315 145.125 ;
        RECT 2019.470 145.080 2019.790 145.140 ;
        RECT 2019.025 144.940 2019.790 145.080 ;
        RECT 2019.025 144.895 2019.315 144.940 ;
        RECT 2019.470 144.880 2019.790 144.940 ;
        RECT 2018.550 96.800 2018.870 96.860 ;
        RECT 2019.010 96.800 2019.330 96.860 ;
        RECT 2018.550 96.660 2019.330 96.800 ;
        RECT 2018.550 96.600 2018.870 96.660 ;
        RECT 2019.010 96.600 2019.330 96.660 ;
        RECT 2019.010 16.900 2019.330 16.960 ;
        RECT 2411.390 16.900 2411.710 16.960 ;
        RECT 2019.010 16.760 2411.710 16.900 ;
        RECT 2019.010 16.700 2019.330 16.760 ;
        RECT 2411.390 16.700 2411.710 16.760 ;
      LAYER via ;
        RECT 1988.220 1212.480 1988.480 1212.740 ;
        RECT 2018.120 1212.480 2018.380 1212.740 ;
        RECT 2018.120 1173.380 2018.380 1173.640 ;
        RECT 2017.660 1172.700 2017.920 1172.960 ;
        RECT 2017.660 1158.760 2017.920 1159.020 ;
        RECT 2018.580 1110.820 2018.840 1111.080 ;
        RECT 2017.660 1075.800 2017.920 1076.060 ;
        RECT 2018.580 1075.800 2018.840 1076.060 ;
        RECT 2017.660 1027.860 2017.920 1028.120 ;
        RECT 2018.580 1027.860 2018.840 1028.120 ;
        RECT 2019.040 965.980 2019.300 966.240 ;
        RECT 2019.960 965.980 2020.220 966.240 ;
        RECT 2019.040 869.420 2019.300 869.680 ;
        RECT 2019.960 869.420 2020.220 869.680 ;
        RECT 2017.660 820.800 2017.920 821.060 ;
        RECT 2018.580 820.800 2018.840 821.060 ;
        RECT 2018.120 690.240 2018.380 690.500 ;
        RECT 2017.660 689.560 2017.920 689.820 ;
        RECT 2016.280 675.960 2016.540 676.220 ;
        RECT 2017.660 675.960 2017.920 676.220 ;
        RECT 2017.200 593.340 2017.460 593.600 ;
        RECT 2017.660 593.000 2017.920 593.260 ;
        RECT 2016.280 579.400 2016.540 579.660 ;
        RECT 2017.660 579.400 2017.920 579.660 ;
        RECT 2017.200 496.780 2017.460 497.040 ;
        RECT 2017.660 496.440 2017.920 496.700 ;
        RECT 2016.280 482.840 2016.540 483.100 ;
        RECT 2017.660 482.840 2017.920 483.100 ;
        RECT 2017.200 400.220 2017.460 400.480 ;
        RECT 2017.660 399.540 2017.920 399.800 ;
        RECT 2017.200 310.460 2017.460 310.720 ;
        RECT 2017.660 310.460 2017.920 310.720 ;
        RECT 2018.120 262.180 2018.380 262.440 ;
        RECT 2018.580 262.180 2018.840 262.440 ;
        RECT 2018.580 241.440 2018.840 241.700 ;
        RECT 2019.040 241.440 2019.300 241.700 ;
        RECT 2019.040 192.820 2019.300 193.080 ;
        RECT 2019.500 144.880 2019.760 145.140 ;
        RECT 2018.580 96.600 2018.840 96.860 ;
        RECT 2019.040 96.600 2019.300 96.860 ;
        RECT 2019.040 16.700 2019.300 16.960 ;
        RECT 2411.420 16.700 2411.680 16.960 ;
      LAYER met2 ;
        RECT 1988.230 1219.680 1988.790 1228.680 ;
        RECT 1988.280 1212.770 1988.420 1219.680 ;
        RECT 1988.220 1212.450 1988.480 1212.770 ;
        RECT 2018.120 1212.450 2018.380 1212.770 ;
        RECT 2018.180 1173.670 2018.320 1212.450 ;
        RECT 2018.120 1173.350 2018.380 1173.670 ;
        RECT 2017.660 1172.670 2017.920 1172.990 ;
        RECT 2017.720 1159.050 2017.860 1172.670 ;
        RECT 2017.660 1158.730 2017.920 1159.050 ;
        RECT 2018.580 1110.790 2018.840 1111.110 ;
        RECT 2018.640 1076.090 2018.780 1110.790 ;
        RECT 2017.660 1075.770 2017.920 1076.090 ;
        RECT 2018.580 1075.770 2018.840 1076.090 ;
        RECT 2017.720 1028.150 2017.860 1075.770 ;
        RECT 2017.660 1027.830 2017.920 1028.150 ;
        RECT 2018.580 1027.830 2018.840 1028.150 ;
        RECT 2018.640 1014.405 2018.780 1027.830 ;
        RECT 2018.570 1014.035 2018.850 1014.405 ;
        RECT 2019.950 1014.035 2020.230 1014.405 ;
        RECT 2020.020 966.270 2020.160 1014.035 ;
        RECT 2019.040 965.950 2019.300 966.270 ;
        RECT 2019.960 965.950 2020.220 966.270 ;
        RECT 2019.100 931.330 2019.240 965.950 ;
        RECT 2018.640 931.190 2019.240 931.330 ;
        RECT 2018.640 917.845 2018.780 931.190 ;
        RECT 2018.570 917.475 2018.850 917.845 ;
        RECT 2019.950 917.475 2020.230 917.845 ;
        RECT 2020.020 869.710 2020.160 917.475 ;
        RECT 2019.040 869.390 2019.300 869.710 ;
        RECT 2019.960 869.390 2020.220 869.710 ;
        RECT 2019.100 834.770 2019.240 869.390 ;
        RECT 2018.640 834.630 2019.240 834.770 ;
        RECT 2018.640 821.090 2018.780 834.630 ;
        RECT 2017.660 820.770 2017.920 821.090 ;
        RECT 2018.580 820.770 2018.840 821.090 ;
        RECT 2017.720 773.005 2017.860 820.770 ;
        RECT 2017.650 772.635 2017.930 773.005 ;
        RECT 2019.030 772.635 2019.310 773.005 ;
        RECT 2019.100 738.210 2019.240 772.635 ;
        RECT 2018.180 738.070 2019.240 738.210 ;
        RECT 2018.180 690.530 2018.320 738.070 ;
        RECT 2018.120 690.210 2018.380 690.530 ;
        RECT 2017.660 689.530 2017.920 689.850 ;
        RECT 2017.720 676.250 2017.860 689.530 ;
        RECT 2016.280 675.930 2016.540 676.250 ;
        RECT 2017.660 675.930 2017.920 676.250 ;
        RECT 2016.340 628.165 2016.480 675.930 ;
        RECT 2016.270 627.795 2016.550 628.165 ;
        RECT 2017.190 627.795 2017.470 628.165 ;
        RECT 2017.260 593.630 2017.400 627.795 ;
        RECT 2017.200 593.310 2017.460 593.630 ;
        RECT 2017.660 592.970 2017.920 593.290 ;
        RECT 2017.720 579.690 2017.860 592.970 ;
        RECT 2016.280 579.370 2016.540 579.690 ;
        RECT 2017.660 579.370 2017.920 579.690 ;
        RECT 2016.340 531.605 2016.480 579.370 ;
        RECT 2016.270 531.235 2016.550 531.605 ;
        RECT 2017.190 531.235 2017.470 531.605 ;
        RECT 2017.260 497.070 2017.400 531.235 ;
        RECT 2017.200 496.750 2017.460 497.070 ;
        RECT 2017.660 496.410 2017.920 496.730 ;
        RECT 2017.720 483.130 2017.860 496.410 ;
        RECT 2016.280 482.810 2016.540 483.130 ;
        RECT 2017.660 482.810 2017.920 483.130 ;
        RECT 2016.340 435.045 2016.480 482.810 ;
        RECT 2016.270 434.675 2016.550 435.045 ;
        RECT 2017.190 434.675 2017.470 435.045 ;
        RECT 2017.260 400.510 2017.400 434.675 ;
        RECT 2017.200 400.190 2017.460 400.510 ;
        RECT 2017.660 399.510 2017.920 399.830 ;
        RECT 2017.720 310.750 2017.860 399.510 ;
        RECT 2017.200 310.430 2017.460 310.750 ;
        RECT 2017.660 310.430 2017.920 310.750 ;
        RECT 2017.260 304.370 2017.400 310.430 ;
        RECT 2017.260 304.230 2018.320 304.370 ;
        RECT 2018.180 262.470 2018.320 304.230 ;
        RECT 2018.120 262.150 2018.380 262.470 ;
        RECT 2018.580 262.150 2018.840 262.470 ;
        RECT 2018.640 241.730 2018.780 262.150 ;
        RECT 2018.580 241.410 2018.840 241.730 ;
        RECT 2019.040 241.410 2019.300 241.730 ;
        RECT 2019.100 241.130 2019.240 241.410 ;
        RECT 2019.100 240.990 2019.700 241.130 ;
        RECT 2019.560 194.325 2019.700 240.990 ;
        RECT 2019.490 193.955 2019.770 194.325 ;
        RECT 2019.030 193.275 2019.310 193.645 ;
        RECT 2019.100 193.110 2019.240 193.275 ;
        RECT 2019.040 192.790 2019.300 193.110 ;
        RECT 2019.500 144.850 2019.760 145.170 ;
        RECT 2019.560 111.250 2019.700 144.850 ;
        RECT 2019.100 111.110 2019.700 111.250 ;
        RECT 2019.100 96.890 2019.240 111.110 ;
        RECT 2018.580 96.570 2018.840 96.890 ;
        RECT 2019.040 96.570 2019.300 96.890 ;
        RECT 2018.640 62.290 2018.780 96.570 ;
        RECT 2018.640 62.150 2019.240 62.290 ;
        RECT 2019.100 16.990 2019.240 62.150 ;
        RECT 2019.040 16.670 2019.300 16.990 ;
        RECT 2411.420 16.670 2411.680 16.990 ;
        RECT 2411.480 2.400 2411.620 16.670 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 2018.570 1014.080 2018.850 1014.360 ;
        RECT 2019.950 1014.080 2020.230 1014.360 ;
        RECT 2018.570 917.520 2018.850 917.800 ;
        RECT 2019.950 917.520 2020.230 917.800 ;
        RECT 2017.650 772.680 2017.930 772.960 ;
        RECT 2019.030 772.680 2019.310 772.960 ;
        RECT 2016.270 627.840 2016.550 628.120 ;
        RECT 2017.190 627.840 2017.470 628.120 ;
        RECT 2016.270 531.280 2016.550 531.560 ;
        RECT 2017.190 531.280 2017.470 531.560 ;
        RECT 2016.270 434.720 2016.550 435.000 ;
        RECT 2017.190 434.720 2017.470 435.000 ;
        RECT 2019.490 194.000 2019.770 194.280 ;
        RECT 2019.030 193.320 2019.310 193.600 ;
      LAYER met3 ;
        RECT 2018.545 1014.370 2018.875 1014.385 ;
        RECT 2019.925 1014.370 2020.255 1014.385 ;
        RECT 2018.545 1014.070 2020.255 1014.370 ;
        RECT 2018.545 1014.055 2018.875 1014.070 ;
        RECT 2019.925 1014.055 2020.255 1014.070 ;
        RECT 2018.545 917.810 2018.875 917.825 ;
        RECT 2019.925 917.810 2020.255 917.825 ;
        RECT 2018.545 917.510 2020.255 917.810 ;
        RECT 2018.545 917.495 2018.875 917.510 ;
        RECT 2019.925 917.495 2020.255 917.510 ;
        RECT 2017.625 772.970 2017.955 772.985 ;
        RECT 2019.005 772.970 2019.335 772.985 ;
        RECT 2017.625 772.670 2019.335 772.970 ;
        RECT 2017.625 772.655 2017.955 772.670 ;
        RECT 2019.005 772.655 2019.335 772.670 ;
        RECT 2016.245 628.130 2016.575 628.145 ;
        RECT 2017.165 628.130 2017.495 628.145 ;
        RECT 2016.245 627.830 2017.495 628.130 ;
        RECT 2016.245 627.815 2016.575 627.830 ;
        RECT 2017.165 627.815 2017.495 627.830 ;
        RECT 2016.245 531.570 2016.575 531.585 ;
        RECT 2017.165 531.570 2017.495 531.585 ;
        RECT 2016.245 531.270 2017.495 531.570 ;
        RECT 2016.245 531.255 2016.575 531.270 ;
        RECT 2017.165 531.255 2017.495 531.270 ;
        RECT 2016.245 435.010 2016.575 435.025 ;
        RECT 2017.165 435.010 2017.495 435.025 ;
        RECT 2016.245 434.710 2017.495 435.010 ;
        RECT 2016.245 434.695 2016.575 434.710 ;
        RECT 2017.165 434.695 2017.495 434.710 ;
        RECT 2019.465 194.290 2019.795 194.305 ;
        RECT 2019.465 193.975 2020.010 194.290 ;
        RECT 2019.005 193.610 2019.335 193.625 ;
        RECT 2019.710 193.610 2020.010 193.975 ;
        RECT 2019.005 193.310 2020.010 193.610 ;
        RECT 2019.005 193.295 2019.335 193.310 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1159.270 1196.700 1159.590 1196.760 ;
        RECT 1162.030 1196.700 1162.350 1196.760 ;
        RECT 1159.270 1196.560 1162.350 1196.700 ;
        RECT 1159.270 1196.500 1159.590 1196.560 ;
        RECT 1162.030 1196.500 1162.350 1196.560 ;
        RECT 805.530 31.860 805.850 31.920 ;
        RECT 1159.270 31.860 1159.590 31.920 ;
        RECT 805.530 31.720 1159.590 31.860 ;
        RECT 805.530 31.660 805.850 31.720 ;
        RECT 1159.270 31.660 1159.590 31.720 ;
      LAYER via ;
        RECT 1159.300 1196.500 1159.560 1196.760 ;
        RECT 1162.060 1196.500 1162.320 1196.760 ;
        RECT 805.560 31.660 805.820 31.920 ;
        RECT 1159.300 31.660 1159.560 31.920 ;
      LAYER met2 ;
        RECT 1163.450 1220.330 1164.010 1228.680 ;
        RECT 1162.120 1220.190 1164.010 1220.330 ;
        RECT 1162.120 1196.790 1162.260 1220.190 ;
        RECT 1163.450 1219.680 1164.010 1220.190 ;
        RECT 1159.300 1196.470 1159.560 1196.790 ;
        RECT 1162.060 1196.470 1162.320 1196.790 ;
        RECT 1159.360 31.950 1159.500 1196.470 ;
        RECT 805.560 31.630 805.820 31.950 ;
        RECT 1159.300 31.630 1159.560 31.950 ;
        RECT 805.620 2.400 805.760 31.630 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 745.270 1196.700 745.590 1196.760 ;
        RECT 749.870 1196.700 750.190 1196.760 ;
        RECT 745.270 1196.560 750.190 1196.700 ;
        RECT 745.270 1196.500 745.590 1196.560 ;
        RECT 749.870 1196.500 750.190 1196.560 ;
        RECT 2.830 24.380 3.150 24.440 ;
        RECT 745.270 24.380 745.590 24.440 ;
        RECT 2.830 24.240 745.590 24.380 ;
        RECT 2.830 24.180 3.150 24.240 ;
        RECT 745.270 24.180 745.590 24.240 ;
      LAYER via ;
        RECT 745.300 1196.500 745.560 1196.760 ;
        RECT 749.900 1196.500 750.160 1196.760 ;
        RECT 2.860 24.180 3.120 24.440 ;
        RECT 745.300 24.180 745.560 24.440 ;
      LAYER met2 ;
        RECT 751.290 1220.330 751.850 1228.680 ;
        RECT 749.960 1220.190 751.850 1220.330 ;
        RECT 749.960 1196.790 750.100 1220.190 ;
        RECT 751.290 1219.680 751.850 1220.190 ;
        RECT 745.300 1196.470 745.560 1196.790 ;
        RECT 749.900 1196.470 750.160 1196.790 ;
        RECT 745.360 24.470 745.500 1196.470 ;
        RECT 2.860 24.150 3.120 24.470 ;
        RECT 745.300 24.150 745.560 24.470 ;
        RECT 2.920 2.400 3.060 24.150 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.040 8.670 24.100 ;
        RECT 752.630 24.040 752.950 24.100 ;
        RECT 8.350 23.900 752.950 24.040 ;
        RECT 8.350 23.840 8.670 23.900 ;
        RECT 752.630 23.840 752.950 23.900 ;
      LAYER via ;
        RECT 8.380 23.840 8.640 24.100 ;
        RECT 752.660 23.840 752.920 24.100 ;
      LAYER met2 ;
        RECT 754.050 1220.330 754.610 1228.680 ;
        RECT 752.260 1220.190 754.610 1220.330 ;
        RECT 752.260 31.180 752.400 1220.190 ;
        RECT 754.050 1219.680 754.610 1220.190 ;
        RECT 752.260 31.040 752.860 31.180 ;
        RECT 752.720 24.130 752.860 31.040 ;
        RECT 8.380 23.810 8.640 24.130 ;
        RECT 752.660 23.810 752.920 24.130 ;
        RECT 8.440 2.400 8.580 23.810 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 753.625 917.745 753.795 1007.335 ;
        RECT 753.625 868.445 753.795 910.775 ;
        RECT 754.085 655.605 754.255 703.715 ;
        RECT 753.625 517.565 753.795 581.655 ;
        RECT 753.625 324.105 753.795 351.475 ;
      LAYER mcon ;
        RECT 753.625 1007.165 753.795 1007.335 ;
        RECT 753.625 910.605 753.795 910.775 ;
        RECT 754.085 703.545 754.255 703.715 ;
        RECT 753.625 581.485 753.795 581.655 ;
        RECT 753.625 351.305 753.795 351.475 ;
      LAYER met1 ;
        RECT 753.550 1196.700 753.870 1196.760 ;
        RECT 755.850 1196.700 756.170 1196.760 ;
        RECT 753.550 1196.560 756.170 1196.700 ;
        RECT 753.550 1196.500 753.870 1196.560 ;
        RECT 755.850 1196.500 756.170 1196.560 ;
        RECT 754.010 1049.140 754.330 1049.200 ;
        RECT 754.470 1049.140 754.790 1049.200 ;
        RECT 754.010 1049.000 754.790 1049.140 ;
        RECT 754.010 1048.940 754.330 1049.000 ;
        RECT 754.470 1048.940 754.790 1049.000 ;
        RECT 754.010 1028.200 754.330 1028.460 ;
        RECT 754.100 1027.780 754.240 1028.200 ;
        RECT 754.010 1027.520 754.330 1027.780 ;
        RECT 753.565 1007.320 753.855 1007.365 ;
        RECT 754.010 1007.320 754.330 1007.380 ;
        RECT 753.565 1007.180 754.330 1007.320 ;
        RECT 753.565 1007.135 753.855 1007.180 ;
        RECT 754.010 1007.120 754.330 1007.180 ;
        RECT 753.565 917.900 753.855 917.945 ;
        RECT 754.010 917.900 754.330 917.960 ;
        RECT 753.565 917.760 754.330 917.900 ;
        RECT 753.565 917.715 753.855 917.760 ;
        RECT 754.010 917.700 754.330 917.760 ;
        RECT 753.565 910.760 753.855 910.805 ;
        RECT 754.010 910.760 754.330 910.820 ;
        RECT 753.565 910.620 754.330 910.760 ;
        RECT 753.565 910.575 753.855 910.620 ;
        RECT 754.010 910.560 754.330 910.620 ;
        RECT 753.550 868.600 753.870 868.660 ;
        RECT 753.355 868.460 753.870 868.600 ;
        RECT 753.550 868.400 753.870 868.460 ;
        RECT 753.550 703.700 753.870 703.760 ;
        RECT 754.025 703.700 754.315 703.745 ;
        RECT 753.550 703.560 754.315 703.700 ;
        RECT 753.550 703.500 753.870 703.560 ;
        RECT 754.025 703.515 754.315 703.560 ;
        RECT 754.010 655.760 754.330 655.820 ;
        RECT 754.010 655.620 754.525 655.760 ;
        RECT 754.010 655.560 754.330 655.620 ;
        RECT 753.550 581.640 753.870 581.700 ;
        RECT 753.355 581.500 753.870 581.640 ;
        RECT 753.550 581.440 753.870 581.500 ;
        RECT 753.565 517.720 753.855 517.765 ;
        RECT 754.010 517.720 754.330 517.780 ;
        RECT 753.565 517.580 754.330 517.720 ;
        RECT 753.565 517.535 753.855 517.580 ;
        RECT 754.010 517.520 754.330 517.580 ;
        RECT 753.550 462.300 753.870 462.360 ;
        RECT 754.930 462.300 755.250 462.360 ;
        RECT 753.550 462.160 755.250 462.300 ;
        RECT 753.550 462.100 753.870 462.160 ;
        RECT 754.930 462.100 755.250 462.160 ;
        RECT 753.550 351.460 753.870 351.520 ;
        RECT 753.355 351.320 753.870 351.460 ;
        RECT 753.550 351.260 753.870 351.320 ;
        RECT 753.550 324.260 753.870 324.320 ;
        RECT 753.355 324.120 753.870 324.260 ;
        RECT 753.550 324.060 753.870 324.120 ;
        RECT 752.630 228.380 752.950 228.440 ;
        RECT 753.550 228.380 753.870 228.440 ;
        RECT 752.630 228.240 753.870 228.380 ;
        RECT 752.630 228.180 752.950 228.240 ;
        RECT 753.550 228.180 753.870 228.240 ;
        RECT 752.630 141.680 752.950 141.740 ;
        RECT 753.550 141.680 753.870 141.740 ;
        RECT 752.630 141.540 753.870 141.680 ;
        RECT 752.630 141.480 752.950 141.540 ;
        RECT 753.550 141.480 753.870 141.540 ;
        RECT 754.010 34.580 754.330 34.640 ;
        RECT 754.470 34.580 754.790 34.640 ;
        RECT 754.010 34.440 754.790 34.580 ;
        RECT 754.010 34.380 754.330 34.440 ;
        RECT 754.470 34.380 754.790 34.440 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 754.010 24.720 754.330 24.780 ;
        RECT 14.330 24.580 754.330 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 754.010 24.520 754.330 24.580 ;
      LAYER via ;
        RECT 753.580 1196.500 753.840 1196.760 ;
        RECT 755.880 1196.500 756.140 1196.760 ;
        RECT 754.040 1048.940 754.300 1049.200 ;
        RECT 754.500 1048.940 754.760 1049.200 ;
        RECT 754.040 1028.200 754.300 1028.460 ;
        RECT 754.040 1027.520 754.300 1027.780 ;
        RECT 754.040 1007.120 754.300 1007.380 ;
        RECT 754.040 917.700 754.300 917.960 ;
        RECT 754.040 910.560 754.300 910.820 ;
        RECT 753.580 868.400 753.840 868.660 ;
        RECT 753.580 703.500 753.840 703.760 ;
        RECT 754.040 655.560 754.300 655.820 ;
        RECT 753.580 581.440 753.840 581.700 ;
        RECT 754.040 517.520 754.300 517.780 ;
        RECT 753.580 462.100 753.840 462.360 ;
        RECT 754.960 462.100 755.220 462.360 ;
        RECT 753.580 351.260 753.840 351.520 ;
        RECT 753.580 324.060 753.840 324.320 ;
        RECT 752.660 228.180 752.920 228.440 ;
        RECT 753.580 228.180 753.840 228.440 ;
        RECT 752.660 141.480 752.920 141.740 ;
        RECT 753.580 141.480 753.840 141.740 ;
        RECT 754.040 34.380 754.300 34.640 ;
        RECT 754.500 34.380 754.760 34.640 ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 754.040 24.520 754.300 24.780 ;
      LAYER met2 ;
        RECT 757.270 1220.330 757.830 1228.680 ;
        RECT 755.940 1220.190 757.830 1220.330 ;
        RECT 755.940 1196.790 756.080 1220.190 ;
        RECT 757.270 1219.680 757.830 1220.190 ;
        RECT 753.580 1196.470 753.840 1196.790 ;
        RECT 755.880 1196.470 756.140 1196.790 ;
        RECT 753.640 1135.330 753.780 1196.470 ;
        RECT 753.640 1135.190 754.700 1135.330 ;
        RECT 754.560 1049.230 754.700 1135.190 ;
        RECT 754.040 1048.910 754.300 1049.230 ;
        RECT 754.500 1048.910 754.760 1049.230 ;
        RECT 754.100 1028.490 754.240 1048.910 ;
        RECT 754.040 1028.170 754.300 1028.490 ;
        RECT 754.040 1027.490 754.300 1027.810 ;
        RECT 754.100 1007.410 754.240 1027.490 ;
        RECT 754.040 1007.090 754.300 1007.410 ;
        RECT 754.040 917.670 754.300 917.990 ;
        RECT 754.100 910.850 754.240 917.670 ;
        RECT 754.040 910.530 754.300 910.850 ;
        RECT 753.580 868.370 753.840 868.690 ;
        RECT 753.640 821.965 753.780 868.370 ;
        RECT 753.570 821.595 753.850 821.965 ;
        RECT 754.030 820.915 754.310 821.285 ;
        RECT 754.100 783.090 754.240 820.915 ;
        RECT 753.640 782.950 754.240 783.090 ;
        RECT 753.640 735.490 753.780 782.950 ;
        RECT 753.640 735.350 754.240 735.490 ;
        RECT 754.100 711.010 754.240 735.350 ;
        RECT 753.640 710.870 754.240 711.010 ;
        RECT 753.640 703.790 753.780 710.870 ;
        RECT 753.580 703.470 753.840 703.790 ;
        RECT 754.040 655.530 754.300 655.850 ;
        RECT 754.100 606.970 754.240 655.530 ;
        RECT 753.640 606.830 754.240 606.970 ;
        RECT 753.640 581.730 753.780 606.830 ;
        RECT 753.580 581.410 753.840 581.730 ;
        RECT 754.040 517.490 754.300 517.810 ;
        RECT 754.100 517.210 754.240 517.490 ;
        RECT 754.100 517.070 755.160 517.210 ;
        RECT 755.020 463.605 755.160 517.070 ;
        RECT 754.950 463.235 755.230 463.605 ;
        RECT 753.570 462.555 753.850 462.925 ;
        RECT 753.640 462.390 753.780 462.555 ;
        RECT 753.580 462.070 753.840 462.390 ;
        RECT 754.960 462.070 755.220 462.390 ;
        RECT 755.020 390.050 755.160 462.070 ;
        RECT 754.100 389.910 755.160 390.050 ;
        RECT 754.100 351.970 754.240 389.910 ;
        RECT 753.640 351.830 754.240 351.970 ;
        RECT 753.640 351.550 753.780 351.830 ;
        RECT 753.580 351.230 753.840 351.550 ;
        RECT 753.580 324.030 753.840 324.350 ;
        RECT 753.640 303.690 753.780 324.030 ;
        RECT 753.640 303.550 754.240 303.690 ;
        RECT 754.100 256.090 754.240 303.550 ;
        RECT 753.640 255.950 754.240 256.090 ;
        RECT 753.640 255.525 753.780 255.950 ;
        RECT 752.650 255.155 752.930 255.525 ;
        RECT 753.570 255.155 753.850 255.525 ;
        RECT 752.720 228.470 752.860 255.155 ;
        RECT 752.660 228.150 752.920 228.470 ;
        RECT 753.580 228.150 753.840 228.470 ;
        RECT 753.640 165.765 753.780 228.150 ;
        RECT 752.650 165.395 752.930 165.765 ;
        RECT 753.570 165.395 753.850 165.765 ;
        RECT 752.720 141.770 752.860 165.395 ;
        RECT 752.660 141.450 752.920 141.770 ;
        RECT 753.580 141.450 753.840 141.770 ;
        RECT 753.640 117.370 753.780 141.450 ;
        RECT 753.640 117.230 754.240 117.370 ;
        RECT 754.100 82.690 754.240 117.230 ;
        RECT 754.100 82.550 754.700 82.690 ;
        RECT 754.560 34.670 754.700 82.550 ;
        RECT 754.040 34.350 754.300 34.670 ;
        RECT 754.500 34.350 754.760 34.670 ;
        RECT 754.100 24.810 754.240 34.350 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 754.040 24.490 754.300 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 753.570 821.640 753.850 821.920 ;
        RECT 754.030 820.960 754.310 821.240 ;
        RECT 754.950 463.280 755.230 463.560 ;
        RECT 753.570 462.600 753.850 462.880 ;
        RECT 752.650 255.200 752.930 255.480 ;
        RECT 753.570 255.200 753.850 255.480 ;
        RECT 752.650 165.440 752.930 165.720 ;
        RECT 753.570 165.440 753.850 165.720 ;
      LAYER met3 ;
        RECT 753.545 821.930 753.875 821.945 ;
        RECT 753.545 821.615 754.090 821.930 ;
        RECT 753.790 821.265 754.090 821.615 ;
        RECT 753.790 820.950 754.335 821.265 ;
        RECT 754.005 820.935 754.335 820.950 ;
        RECT 754.925 463.570 755.255 463.585 ;
        RECT 752.870 463.270 755.255 463.570 ;
        RECT 752.870 462.890 753.170 463.270 ;
        RECT 754.925 463.255 755.255 463.270 ;
        RECT 753.545 462.890 753.875 462.905 ;
        RECT 752.870 462.590 753.875 462.890 ;
        RECT 753.545 462.575 753.875 462.590 ;
        RECT 752.625 255.490 752.955 255.505 ;
        RECT 753.545 255.490 753.875 255.505 ;
        RECT 752.625 255.190 753.875 255.490 ;
        RECT 752.625 255.175 752.955 255.190 ;
        RECT 753.545 255.175 753.875 255.190 ;
        RECT 752.625 165.730 752.955 165.745 ;
        RECT 753.545 165.730 753.875 165.745 ;
        RECT 752.625 165.430 753.875 165.730 ;
        RECT 752.625 165.415 752.955 165.430 ;
        RECT 753.545 165.415 753.875 165.430 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 710.770 25.060 711.090 25.120 ;
        RECT 38.250 24.920 711.090 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 710.770 24.860 711.090 24.920 ;
        RECT 754.470 24.720 754.790 24.780 ;
        RECT 765.970 24.720 766.290 24.780 ;
        RECT 754.470 24.580 766.290 24.720 ;
        RECT 754.470 24.520 754.790 24.580 ;
        RECT 765.970 24.520 766.290 24.580 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 710.800 24.860 711.060 25.120 ;
        RECT 754.500 24.520 754.760 24.780 ;
        RECT 766.000 24.520 766.260 24.780 ;
      LAYER met2 ;
        RECT 769.230 1220.330 769.790 1228.680 ;
        RECT 767.440 1220.190 769.790 1220.330 ;
        RECT 767.440 1196.530 767.580 1220.190 ;
        RECT 769.230 1219.680 769.790 1220.190 ;
        RECT 766.060 1196.390 767.580 1196.530 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 710.800 25.005 711.060 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 710.790 24.635 711.070 25.005 ;
        RECT 754.490 24.635 754.770 25.005 ;
        RECT 766.060 24.810 766.200 1196.390 ;
        RECT 754.500 24.490 754.760 24.635 ;
        RECT 766.000 24.490 766.260 24.810 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 710.790 24.680 711.070 24.960 ;
        RECT 754.490 24.680 754.770 24.960 ;
      LAYER met3 ;
        RECT 710.765 24.970 711.095 24.985 ;
        RECT 754.465 24.970 754.795 24.985 ;
        RECT 710.765 24.670 754.795 24.970 ;
        RECT 710.765 24.655 711.095 24.670 ;
        RECT 754.465 24.655 754.795 24.670 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 870.005 786.505 870.175 821.015 ;
        RECT 870.005 689.605 870.175 724.455 ;
        RECT 870.005 593.045 870.175 627.895 ;
        RECT 870.005 496.485 870.175 531.335 ;
        RECT 870.005 386.325 870.175 434.775 ;
        RECT 870.005 241.485 870.175 289.595 ;
        RECT 870.005 144.925 870.175 169.235 ;
        RECT 870.005 110.245 870.175 137.955 ;
      LAYER mcon ;
        RECT 870.005 820.845 870.175 821.015 ;
        RECT 870.005 724.285 870.175 724.455 ;
        RECT 870.005 627.725 870.175 627.895 ;
        RECT 870.005 531.165 870.175 531.335 ;
        RECT 870.005 434.605 870.175 434.775 ;
        RECT 870.005 289.425 870.175 289.595 ;
        RECT 870.005 169.065 870.175 169.235 ;
        RECT 870.005 137.785 870.175 137.955 ;
      LAYER met1 ;
        RECT 870.390 1159.300 870.710 1159.360 ;
        RECT 871.770 1159.300 872.090 1159.360 ;
        RECT 870.390 1159.160 872.090 1159.300 ;
        RECT 870.390 1159.100 870.710 1159.160 ;
        RECT 871.770 1159.100 872.090 1159.160 ;
        RECT 869.470 1028.400 869.790 1028.460 ;
        RECT 870.390 1028.400 870.710 1028.460 ;
        RECT 869.470 1028.260 870.710 1028.400 ;
        RECT 869.470 1028.200 869.790 1028.260 ;
        RECT 870.390 1028.200 870.710 1028.260 ;
        RECT 869.470 931.840 869.790 931.900 ;
        RECT 870.390 931.840 870.710 931.900 ;
        RECT 869.470 931.700 870.710 931.840 ;
        RECT 869.470 931.640 869.790 931.700 ;
        RECT 870.390 931.640 870.710 931.700 ;
        RECT 870.390 869.620 870.710 869.680 ;
        RECT 871.310 869.620 871.630 869.680 ;
        RECT 870.390 869.480 871.630 869.620 ;
        RECT 870.390 869.420 870.710 869.480 ;
        RECT 871.310 869.420 871.630 869.480 ;
        RECT 869.470 835.280 869.790 835.340 ;
        RECT 870.390 835.280 870.710 835.340 ;
        RECT 869.470 835.140 870.710 835.280 ;
        RECT 869.470 835.080 869.790 835.140 ;
        RECT 870.390 835.080 870.710 835.140 ;
        RECT 869.930 821.000 870.250 821.060 ;
        RECT 869.735 820.860 870.250 821.000 ;
        RECT 869.930 820.800 870.250 820.860 ;
        RECT 869.930 786.660 870.250 786.720 ;
        RECT 869.735 786.520 870.250 786.660 ;
        RECT 869.930 786.460 870.250 786.520 ;
        RECT 869.470 738.380 869.790 738.440 ;
        RECT 870.390 738.380 870.710 738.440 ;
        RECT 869.470 738.240 870.710 738.380 ;
        RECT 869.470 738.180 869.790 738.240 ;
        RECT 870.390 738.180 870.710 738.240 ;
        RECT 869.930 724.440 870.250 724.500 ;
        RECT 869.735 724.300 870.250 724.440 ;
        RECT 869.930 724.240 870.250 724.300 ;
        RECT 869.930 689.760 870.250 689.820 ;
        RECT 869.735 689.620 870.250 689.760 ;
        RECT 869.930 689.560 870.250 689.620 ;
        RECT 869.470 641.820 869.790 641.880 ;
        RECT 870.390 641.820 870.710 641.880 ;
        RECT 869.470 641.680 870.710 641.820 ;
        RECT 869.470 641.620 869.790 641.680 ;
        RECT 870.390 641.620 870.710 641.680 ;
        RECT 869.930 627.880 870.250 627.940 ;
        RECT 869.735 627.740 870.250 627.880 ;
        RECT 869.930 627.680 870.250 627.740 ;
        RECT 869.930 593.200 870.250 593.260 ;
        RECT 869.735 593.060 870.250 593.200 ;
        RECT 869.930 593.000 870.250 593.060 ;
        RECT 869.470 545.260 869.790 545.320 ;
        RECT 870.390 545.260 870.710 545.320 ;
        RECT 869.470 545.120 870.710 545.260 ;
        RECT 869.470 545.060 869.790 545.120 ;
        RECT 870.390 545.060 870.710 545.120 ;
        RECT 869.930 531.320 870.250 531.380 ;
        RECT 869.735 531.180 870.250 531.320 ;
        RECT 869.930 531.120 870.250 531.180 ;
        RECT 869.930 496.640 870.250 496.700 ;
        RECT 869.735 496.500 870.250 496.640 ;
        RECT 869.930 496.440 870.250 496.500 ;
        RECT 869.470 448.700 869.790 448.760 ;
        RECT 870.390 448.700 870.710 448.760 ;
        RECT 869.470 448.560 870.710 448.700 ;
        RECT 869.470 448.500 869.790 448.560 ;
        RECT 870.390 448.500 870.710 448.560 ;
        RECT 869.930 434.760 870.250 434.820 ;
        RECT 869.735 434.620 870.250 434.760 ;
        RECT 869.930 434.560 870.250 434.620 ;
        RECT 869.945 386.480 870.235 386.525 ;
        RECT 870.390 386.480 870.710 386.540 ;
        RECT 869.945 386.340 870.710 386.480 ;
        RECT 869.945 386.295 870.235 386.340 ;
        RECT 870.390 386.280 870.710 386.340 ;
        RECT 869.930 338.200 870.250 338.260 ;
        RECT 870.390 338.200 870.710 338.260 ;
        RECT 869.930 338.060 870.710 338.200 ;
        RECT 869.930 338.000 870.250 338.060 ;
        RECT 870.390 338.000 870.710 338.060 ;
        RECT 869.945 289.580 870.235 289.625 ;
        RECT 870.390 289.580 870.710 289.640 ;
        RECT 869.945 289.440 870.710 289.580 ;
        RECT 869.945 289.395 870.235 289.440 ;
        RECT 870.390 289.380 870.710 289.440 ;
        RECT 869.930 241.640 870.250 241.700 ;
        RECT 869.735 241.500 870.250 241.640 ;
        RECT 869.930 241.440 870.250 241.500 ;
        RECT 869.945 169.220 870.235 169.265 ;
        RECT 870.390 169.220 870.710 169.280 ;
        RECT 869.945 169.080 870.710 169.220 ;
        RECT 869.945 169.035 870.235 169.080 ;
        RECT 870.390 169.020 870.710 169.080 ;
        RECT 869.930 145.080 870.250 145.140 ;
        RECT 869.735 144.940 870.250 145.080 ;
        RECT 869.930 144.880 870.250 144.940 ;
        RECT 869.930 137.940 870.250 138.000 ;
        RECT 869.735 137.800 870.250 137.940 ;
        RECT 869.930 137.740 870.250 137.800 ;
        RECT 869.930 110.400 870.250 110.460 ;
        RECT 869.735 110.260 870.250 110.400 ;
        RECT 869.930 110.200 870.250 110.260 ;
        RECT 240.650 27.100 240.970 27.160 ;
        RECT 869.930 27.100 870.250 27.160 ;
        RECT 240.650 26.960 870.250 27.100 ;
        RECT 240.650 26.900 240.970 26.960 ;
        RECT 869.930 26.900 870.250 26.960 ;
      LAYER via ;
        RECT 870.420 1159.100 870.680 1159.360 ;
        RECT 871.800 1159.100 872.060 1159.360 ;
        RECT 869.500 1028.200 869.760 1028.460 ;
        RECT 870.420 1028.200 870.680 1028.460 ;
        RECT 869.500 931.640 869.760 931.900 ;
        RECT 870.420 931.640 870.680 931.900 ;
        RECT 870.420 869.420 870.680 869.680 ;
        RECT 871.340 869.420 871.600 869.680 ;
        RECT 869.500 835.080 869.760 835.340 ;
        RECT 870.420 835.080 870.680 835.340 ;
        RECT 869.960 820.800 870.220 821.060 ;
        RECT 869.960 786.460 870.220 786.720 ;
        RECT 869.500 738.180 869.760 738.440 ;
        RECT 870.420 738.180 870.680 738.440 ;
        RECT 869.960 724.240 870.220 724.500 ;
        RECT 869.960 689.560 870.220 689.820 ;
        RECT 869.500 641.620 869.760 641.880 ;
        RECT 870.420 641.620 870.680 641.880 ;
        RECT 869.960 627.680 870.220 627.940 ;
        RECT 869.960 593.000 870.220 593.260 ;
        RECT 869.500 545.060 869.760 545.320 ;
        RECT 870.420 545.060 870.680 545.320 ;
        RECT 869.960 531.120 870.220 531.380 ;
        RECT 869.960 496.440 870.220 496.700 ;
        RECT 869.500 448.500 869.760 448.760 ;
        RECT 870.420 448.500 870.680 448.760 ;
        RECT 869.960 434.560 870.220 434.820 ;
        RECT 870.420 386.280 870.680 386.540 ;
        RECT 869.960 338.000 870.220 338.260 ;
        RECT 870.420 338.000 870.680 338.260 ;
        RECT 870.420 289.380 870.680 289.640 ;
        RECT 869.960 241.440 870.220 241.700 ;
        RECT 870.420 169.020 870.680 169.280 ;
        RECT 869.960 144.880 870.220 145.140 ;
        RECT 869.960 137.740 870.220 138.000 ;
        RECT 869.960 110.200 870.220 110.460 ;
        RECT 240.680 26.900 240.940 27.160 ;
        RECT 869.960 26.900 870.220 27.160 ;
      LAYER met2 ;
        RECT 873.190 1220.330 873.750 1228.680 ;
        RECT 871.860 1220.190 873.750 1220.330 ;
        RECT 871.860 1159.390 872.000 1220.190 ;
        RECT 873.190 1219.680 873.750 1220.190 ;
        RECT 870.420 1159.070 870.680 1159.390 ;
        RECT 871.800 1159.070 872.060 1159.390 ;
        RECT 870.480 1028.490 870.620 1159.070 ;
        RECT 869.500 1028.170 869.760 1028.490 ;
        RECT 870.420 1028.170 870.680 1028.490 ;
        RECT 869.560 1027.890 869.700 1028.170 ;
        RECT 869.560 1027.750 870.160 1027.890 ;
        RECT 870.020 980.290 870.160 1027.750 ;
        RECT 870.020 980.150 870.620 980.290 ;
        RECT 870.480 931.930 870.620 980.150 ;
        RECT 869.500 931.610 869.760 931.930 ;
        RECT 870.420 931.610 870.680 931.930 ;
        RECT 869.560 931.330 869.700 931.610 ;
        RECT 869.560 931.190 870.160 931.330 ;
        RECT 870.020 917.845 870.160 931.190 ;
        RECT 869.950 917.475 870.230 917.845 ;
        RECT 871.330 917.475 871.610 917.845 ;
        RECT 871.400 869.710 871.540 917.475 ;
        RECT 870.420 869.390 870.680 869.710 ;
        RECT 871.340 869.390 871.600 869.710 ;
        RECT 870.480 835.370 870.620 869.390 ;
        RECT 869.500 835.050 869.760 835.370 ;
        RECT 870.420 835.050 870.680 835.370 ;
        RECT 869.560 834.770 869.700 835.050 ;
        RECT 869.560 834.630 870.160 834.770 ;
        RECT 870.020 821.090 870.160 834.630 ;
        RECT 869.960 820.770 870.220 821.090 ;
        RECT 869.960 786.430 870.220 786.750 ;
        RECT 870.020 772.890 870.160 786.430 ;
        RECT 870.020 772.750 870.620 772.890 ;
        RECT 870.480 738.470 870.620 772.750 ;
        RECT 869.500 738.210 869.760 738.470 ;
        RECT 869.500 738.150 870.160 738.210 ;
        RECT 870.420 738.150 870.680 738.470 ;
        RECT 869.560 738.070 870.160 738.150 ;
        RECT 870.020 724.530 870.160 738.070 ;
        RECT 869.960 724.210 870.220 724.530 ;
        RECT 869.960 689.530 870.220 689.850 ;
        RECT 870.020 676.330 870.160 689.530 ;
        RECT 870.020 676.190 870.620 676.330 ;
        RECT 870.480 641.910 870.620 676.190 ;
        RECT 869.500 641.650 869.760 641.910 ;
        RECT 869.500 641.590 870.160 641.650 ;
        RECT 870.420 641.590 870.680 641.910 ;
        RECT 869.560 641.510 870.160 641.590 ;
        RECT 870.020 627.970 870.160 641.510 ;
        RECT 869.960 627.650 870.220 627.970 ;
        RECT 869.960 592.970 870.220 593.290 ;
        RECT 870.020 579.770 870.160 592.970 ;
        RECT 870.020 579.630 870.620 579.770 ;
        RECT 870.480 545.350 870.620 579.630 ;
        RECT 869.500 545.090 869.760 545.350 ;
        RECT 869.500 545.030 870.160 545.090 ;
        RECT 870.420 545.030 870.680 545.350 ;
        RECT 869.560 544.950 870.160 545.030 ;
        RECT 870.020 531.410 870.160 544.950 ;
        RECT 869.960 531.090 870.220 531.410 ;
        RECT 869.960 496.410 870.220 496.730 ;
        RECT 870.020 483.210 870.160 496.410 ;
        RECT 870.020 483.070 870.620 483.210 ;
        RECT 870.480 448.790 870.620 483.070 ;
        RECT 869.500 448.530 869.760 448.790 ;
        RECT 869.500 448.470 870.160 448.530 ;
        RECT 870.420 448.470 870.680 448.790 ;
        RECT 869.560 448.390 870.160 448.470 ;
        RECT 870.020 434.850 870.160 448.390 ;
        RECT 869.960 434.530 870.220 434.850 ;
        RECT 870.420 386.250 870.680 386.570 ;
        RECT 870.480 338.290 870.620 386.250 ;
        RECT 869.960 337.970 870.220 338.290 ;
        RECT 870.420 337.970 870.680 338.290 ;
        RECT 870.020 303.690 870.160 337.970 ;
        RECT 870.020 303.550 870.620 303.690 ;
        RECT 870.480 289.670 870.620 303.550 ;
        RECT 870.420 289.350 870.680 289.670 ;
        RECT 869.960 241.410 870.220 241.730 ;
        RECT 870.020 207.130 870.160 241.410 ;
        RECT 870.020 206.990 870.620 207.130 ;
        RECT 870.480 169.310 870.620 206.990 ;
        RECT 870.420 168.990 870.680 169.310 ;
        RECT 869.960 144.850 870.220 145.170 ;
        RECT 870.020 138.030 870.160 144.850 ;
        RECT 869.960 137.710 870.220 138.030 ;
        RECT 869.960 110.170 870.220 110.490 ;
        RECT 870.020 27.190 870.160 110.170 ;
        RECT 240.680 26.870 240.940 27.190 ;
        RECT 869.960 26.870 870.220 27.190 ;
        RECT 240.740 2.400 240.880 26.870 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 869.950 917.520 870.230 917.800 ;
        RECT 871.330 917.520 871.610 917.800 ;
      LAYER met3 ;
        RECT 869.925 917.810 870.255 917.825 ;
        RECT 871.305 917.810 871.635 917.825 ;
        RECT 869.925 917.510 871.635 917.810 ;
        RECT 869.925 917.495 870.255 917.510 ;
        RECT 871.305 917.495 871.635 917.510 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 27.440 258.450 27.500 ;
        RECT 877.290 27.440 877.610 27.500 ;
        RECT 258.130 27.300 877.610 27.440 ;
        RECT 258.130 27.240 258.450 27.300 ;
        RECT 877.290 27.240 877.610 27.300 ;
      LAYER via ;
        RECT 258.160 27.240 258.420 27.500 ;
        RECT 877.320 27.240 877.580 27.500 ;
      LAYER met2 ;
        RECT 882.390 1220.330 882.950 1228.680 ;
        RECT 880.140 1220.190 882.950 1220.330 ;
        RECT 880.140 1196.530 880.280 1220.190 ;
        RECT 882.390 1219.680 882.950 1220.190 ;
        RECT 877.380 1196.390 880.280 1196.530 ;
        RECT 877.380 27.530 877.520 1196.390 ;
        RECT 258.160 27.210 258.420 27.530 ;
        RECT 877.320 27.210 877.580 27.530 ;
        RECT 258.220 2.400 258.360 27.210 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 23.700 276.390 23.760 ;
        RECT 890.170 23.700 890.490 23.760 ;
        RECT 276.070 23.560 890.490 23.700 ;
        RECT 276.070 23.500 276.390 23.560 ;
        RECT 890.170 23.500 890.490 23.560 ;
      LAYER via ;
        RECT 276.100 23.500 276.360 23.760 ;
        RECT 890.200 23.500 890.460 23.760 ;
      LAYER met2 ;
        RECT 891.590 1220.330 892.150 1228.680 ;
        RECT 890.260 1220.190 892.150 1220.330 ;
        RECT 890.260 23.790 890.400 1220.190 ;
        RECT 891.590 1219.680 892.150 1220.190 ;
        RECT 276.100 23.470 276.360 23.790 ;
        RECT 890.200 23.470 890.460 23.790 ;
        RECT 276.160 2.400 276.300 23.470 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 897.605 1062.585 897.775 1077.035 ;
        RECT 897.605 89.845 897.775 137.955 ;
      LAYER mcon ;
        RECT 897.605 1076.865 897.775 1077.035 ;
        RECT 897.605 137.785 897.775 137.955 ;
      LAYER met1 ;
        RECT 897.990 1159.300 898.310 1159.360 ;
        RECT 899.370 1159.300 899.690 1159.360 ;
        RECT 897.990 1159.160 899.690 1159.300 ;
        RECT 897.990 1159.100 898.310 1159.160 ;
        RECT 899.370 1159.100 899.690 1159.160 ;
        RECT 897.990 1111.020 898.310 1111.080 ;
        RECT 898.910 1111.020 899.230 1111.080 ;
        RECT 897.990 1110.880 899.230 1111.020 ;
        RECT 897.990 1110.820 898.310 1110.880 ;
        RECT 898.910 1110.820 899.230 1110.880 ;
        RECT 897.545 1077.020 897.835 1077.065 ;
        RECT 897.990 1077.020 898.310 1077.080 ;
        RECT 897.545 1076.880 898.310 1077.020 ;
        RECT 897.545 1076.835 897.835 1076.880 ;
        RECT 897.990 1076.820 898.310 1076.880 ;
        RECT 897.530 1062.740 897.850 1062.800 ;
        RECT 897.335 1062.600 897.850 1062.740 ;
        RECT 897.530 1062.540 897.850 1062.600 ;
        RECT 897.530 255.720 897.850 255.980 ;
        RECT 897.620 255.300 897.760 255.720 ;
        RECT 897.530 255.040 897.850 255.300 ;
        RECT 897.990 145.420 898.310 145.480 ;
        RECT 897.620 145.280 898.310 145.420 ;
        RECT 897.620 145.140 897.760 145.280 ;
        RECT 897.990 145.220 898.310 145.280 ;
        RECT 897.530 144.880 897.850 145.140 ;
        RECT 897.530 137.940 897.850 138.000 ;
        RECT 897.335 137.800 897.850 137.940 ;
        RECT 897.530 137.740 897.850 137.800 ;
        RECT 897.530 90.000 897.850 90.060 ;
        RECT 897.335 89.860 897.850 90.000 ;
        RECT 897.530 89.800 897.850 89.860 ;
        RECT 294.010 23.360 294.330 23.420 ;
        RECT 897.530 23.360 897.850 23.420 ;
        RECT 294.010 23.220 897.850 23.360 ;
        RECT 294.010 23.160 294.330 23.220 ;
        RECT 897.530 23.160 897.850 23.220 ;
      LAYER via ;
        RECT 898.020 1159.100 898.280 1159.360 ;
        RECT 899.400 1159.100 899.660 1159.360 ;
        RECT 898.020 1110.820 898.280 1111.080 ;
        RECT 898.940 1110.820 899.200 1111.080 ;
        RECT 898.020 1076.820 898.280 1077.080 ;
        RECT 897.560 1062.540 897.820 1062.800 ;
        RECT 897.560 255.720 897.820 255.980 ;
        RECT 897.560 255.040 897.820 255.300 ;
        RECT 898.020 145.220 898.280 145.480 ;
        RECT 897.560 144.880 897.820 145.140 ;
        RECT 897.560 137.740 897.820 138.000 ;
        RECT 897.560 89.800 897.820 90.060 ;
        RECT 294.040 23.160 294.300 23.420 ;
        RECT 897.560 23.160 897.820 23.420 ;
      LAYER met2 ;
        RECT 900.790 1221.010 901.350 1228.680 ;
        RECT 898.540 1220.870 901.350 1221.010 ;
        RECT 898.540 1207.525 898.680 1220.870 ;
        RECT 900.790 1219.680 901.350 1220.870 ;
        RECT 898.470 1207.155 898.750 1207.525 ;
        RECT 899.390 1207.155 899.670 1207.525 ;
        RECT 899.460 1159.390 899.600 1207.155 ;
        RECT 898.020 1159.245 898.280 1159.390 ;
        RECT 898.010 1158.875 898.290 1159.245 ;
        RECT 898.930 1158.875 899.210 1159.245 ;
        RECT 899.400 1159.070 899.660 1159.390 ;
        RECT 899.000 1111.110 899.140 1158.875 ;
        RECT 898.020 1110.790 898.280 1111.110 ;
        RECT 898.940 1110.790 899.200 1111.110 ;
        RECT 898.080 1077.110 898.220 1110.790 ;
        RECT 898.020 1076.790 898.280 1077.110 ;
        RECT 897.560 1062.510 897.820 1062.830 ;
        RECT 897.620 1028.570 897.760 1062.510 ;
        RECT 897.160 1028.430 897.760 1028.570 ;
        RECT 897.160 1027.890 897.300 1028.430 ;
        RECT 897.160 1027.750 897.760 1027.890 ;
        RECT 897.620 932.010 897.760 1027.750 ;
        RECT 897.160 931.870 897.760 932.010 ;
        RECT 897.160 931.330 897.300 931.870 ;
        RECT 897.160 931.190 897.760 931.330 ;
        RECT 897.620 835.450 897.760 931.190 ;
        RECT 897.160 835.310 897.760 835.450 ;
        RECT 897.160 834.770 897.300 835.310 ;
        RECT 897.160 834.630 897.760 834.770 ;
        RECT 897.620 738.890 897.760 834.630 ;
        RECT 897.160 738.750 897.760 738.890 ;
        RECT 897.160 738.210 897.300 738.750 ;
        RECT 897.160 738.070 897.760 738.210 ;
        RECT 897.620 642.330 897.760 738.070 ;
        RECT 897.160 642.190 897.760 642.330 ;
        RECT 897.160 641.650 897.300 642.190 ;
        RECT 897.160 641.510 897.760 641.650 ;
        RECT 897.620 545.770 897.760 641.510 ;
        RECT 897.160 545.630 897.760 545.770 ;
        RECT 897.160 545.090 897.300 545.630 ;
        RECT 897.160 544.950 897.760 545.090 ;
        RECT 897.620 449.210 897.760 544.950 ;
        RECT 897.160 449.070 897.760 449.210 ;
        RECT 897.160 448.530 897.300 449.070 ;
        RECT 897.160 448.390 897.760 448.530 ;
        RECT 897.620 351.970 897.760 448.390 ;
        RECT 897.160 351.830 897.760 351.970 ;
        RECT 897.160 351.290 897.300 351.830 ;
        RECT 897.160 351.150 897.760 351.290 ;
        RECT 897.620 256.010 897.760 351.150 ;
        RECT 897.560 255.690 897.820 256.010 ;
        RECT 897.560 255.010 897.820 255.330 ;
        RECT 897.620 207.130 897.760 255.010 ;
        RECT 897.620 206.990 898.220 207.130 ;
        RECT 898.080 145.510 898.220 206.990 ;
        RECT 898.020 145.190 898.280 145.510 ;
        RECT 897.560 144.850 897.820 145.170 ;
        RECT 897.620 138.030 897.760 144.850 ;
        RECT 897.560 137.710 897.820 138.030 ;
        RECT 897.560 89.770 897.820 90.090 ;
        RECT 897.620 23.450 897.760 89.770 ;
        RECT 294.040 23.130 294.300 23.450 ;
        RECT 897.560 23.130 897.820 23.450 ;
        RECT 294.100 2.400 294.240 23.130 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 898.470 1207.200 898.750 1207.480 ;
        RECT 899.390 1207.200 899.670 1207.480 ;
        RECT 898.010 1158.920 898.290 1159.200 ;
        RECT 898.930 1158.920 899.210 1159.200 ;
      LAYER met3 ;
        RECT 898.445 1207.490 898.775 1207.505 ;
        RECT 899.365 1207.490 899.695 1207.505 ;
        RECT 898.445 1207.190 899.695 1207.490 ;
        RECT 898.445 1207.175 898.775 1207.190 ;
        RECT 899.365 1207.175 899.695 1207.190 ;
        RECT 897.985 1159.210 898.315 1159.225 ;
        RECT 898.905 1159.210 899.235 1159.225 ;
        RECT 897.985 1158.910 899.235 1159.210 ;
        RECT 897.985 1158.895 898.315 1158.910 ;
        RECT 898.905 1158.895 899.235 1158.910 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 22.680 312.270 22.740 ;
        RECT 904.890 22.680 905.210 22.740 ;
        RECT 311.950 22.540 905.210 22.680 ;
        RECT 311.950 22.480 312.270 22.540 ;
        RECT 904.890 22.480 905.210 22.540 ;
      LAYER via ;
        RECT 311.980 22.480 312.240 22.740 ;
        RECT 904.920 22.480 905.180 22.740 ;
      LAYER met2 ;
        RECT 909.990 1220.330 910.550 1228.680 ;
        RECT 907.740 1220.190 910.550 1220.330 ;
        RECT 907.740 1196.530 907.880 1220.190 ;
        RECT 909.990 1219.680 910.550 1220.190 ;
        RECT 904.980 1196.390 907.880 1196.530 ;
        RECT 904.980 22.770 905.120 1196.390 ;
        RECT 311.980 22.450 312.240 22.770 ;
        RECT 904.920 22.450 905.180 22.770 ;
        RECT 312.040 2.400 312.180 22.450 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 23.020 330.210 23.080 ;
        RECT 917.770 23.020 918.090 23.080 ;
        RECT 329.890 22.880 918.090 23.020 ;
        RECT 329.890 22.820 330.210 22.880 ;
        RECT 917.770 22.820 918.090 22.880 ;
      LAYER via ;
        RECT 329.920 22.820 330.180 23.080 ;
        RECT 917.800 22.820 918.060 23.080 ;
      LAYER met2 ;
        RECT 919.190 1220.330 919.750 1228.680 ;
        RECT 917.860 1220.190 919.750 1220.330 ;
        RECT 917.860 23.110 918.000 1220.190 ;
        RECT 919.190 1219.680 919.750 1220.190 ;
        RECT 329.920 22.790 330.180 23.110 ;
        RECT 917.800 22.790 918.060 23.110 ;
        RECT 329.980 2.400 330.120 22.790 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 925.590 1159.300 925.910 1159.360 ;
        RECT 926.970 1159.300 927.290 1159.360 ;
        RECT 925.590 1159.160 927.290 1159.300 ;
        RECT 925.590 1159.100 925.910 1159.160 ;
        RECT 926.970 1159.100 927.290 1159.160 ;
        RECT 925.590 1111.020 925.910 1111.080 ;
        RECT 926.510 1111.020 926.830 1111.080 ;
        RECT 925.590 1110.880 926.830 1111.020 ;
        RECT 925.590 1110.820 925.910 1110.880 ;
        RECT 926.510 1110.820 926.830 1110.880 ;
        RECT 925.590 1062.740 925.910 1062.800 ;
        RECT 926.050 1062.740 926.370 1062.800 ;
        RECT 925.590 1062.600 926.370 1062.740 ;
        RECT 925.590 1062.540 925.910 1062.600 ;
        RECT 926.050 1062.540 926.370 1062.600 ;
        RECT 347.370 22.340 347.690 22.400 ;
        RECT 926.050 22.340 926.370 22.400 ;
        RECT 347.370 22.200 926.370 22.340 ;
        RECT 347.370 22.140 347.690 22.200 ;
        RECT 926.050 22.140 926.370 22.200 ;
      LAYER via ;
        RECT 925.620 1159.100 925.880 1159.360 ;
        RECT 927.000 1159.100 927.260 1159.360 ;
        RECT 925.620 1110.820 925.880 1111.080 ;
        RECT 926.540 1110.820 926.800 1111.080 ;
        RECT 925.620 1062.540 925.880 1062.800 ;
        RECT 926.080 1062.540 926.340 1062.800 ;
        RECT 347.400 22.140 347.660 22.400 ;
        RECT 926.080 22.140 926.340 22.400 ;
      LAYER met2 ;
        RECT 928.390 1221.010 928.950 1228.680 ;
        RECT 926.140 1220.870 928.950 1221.010 ;
        RECT 926.140 1207.525 926.280 1220.870 ;
        RECT 928.390 1219.680 928.950 1220.870 ;
        RECT 926.070 1207.155 926.350 1207.525 ;
        RECT 926.990 1207.155 927.270 1207.525 ;
        RECT 927.060 1159.390 927.200 1207.155 ;
        RECT 925.620 1159.245 925.880 1159.390 ;
        RECT 925.610 1158.875 925.890 1159.245 ;
        RECT 926.530 1158.875 926.810 1159.245 ;
        RECT 927.000 1159.070 927.260 1159.390 ;
        RECT 926.600 1111.110 926.740 1158.875 ;
        RECT 925.620 1110.790 925.880 1111.110 ;
        RECT 926.540 1110.790 926.800 1111.110 ;
        RECT 925.680 1062.830 925.820 1110.790 ;
        RECT 925.620 1062.510 925.880 1062.830 ;
        RECT 926.080 1062.510 926.340 1062.830 ;
        RECT 926.140 883.050 926.280 1062.510 ;
        RECT 925.680 882.910 926.280 883.050 ;
        RECT 925.680 881.690 925.820 882.910 ;
        RECT 925.680 881.550 926.280 881.690 ;
        RECT 926.140 787.170 926.280 881.550 ;
        RECT 925.680 787.030 926.280 787.170 ;
        RECT 925.680 786.490 925.820 787.030 ;
        RECT 925.680 786.350 926.280 786.490 ;
        RECT 926.140 690.610 926.280 786.350 ;
        RECT 925.680 690.470 926.280 690.610 ;
        RECT 925.680 688.570 925.820 690.470 ;
        RECT 925.680 688.430 926.280 688.570 ;
        RECT 926.140 594.050 926.280 688.430 ;
        RECT 925.680 593.910 926.280 594.050 ;
        RECT 925.680 593.370 925.820 593.910 ;
        RECT 925.680 593.230 926.280 593.370 ;
        RECT 926.140 303.690 926.280 593.230 ;
        RECT 925.680 303.550 926.280 303.690 ;
        RECT 925.680 303.010 925.820 303.550 ;
        RECT 925.680 302.870 926.280 303.010 ;
        RECT 926.140 110.570 926.280 302.870 ;
        RECT 925.680 110.430 926.280 110.570 ;
        RECT 925.680 109.890 925.820 110.430 ;
        RECT 925.680 109.750 926.280 109.890 ;
        RECT 926.140 22.430 926.280 109.750 ;
        RECT 347.400 22.110 347.660 22.430 ;
        RECT 926.080 22.110 926.340 22.430 ;
        RECT 347.460 2.400 347.600 22.110 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 926.070 1207.200 926.350 1207.480 ;
        RECT 926.990 1207.200 927.270 1207.480 ;
        RECT 925.610 1158.920 925.890 1159.200 ;
        RECT 926.530 1158.920 926.810 1159.200 ;
      LAYER met3 ;
        RECT 926.045 1207.490 926.375 1207.505 ;
        RECT 926.965 1207.490 927.295 1207.505 ;
        RECT 926.045 1207.190 927.295 1207.490 ;
        RECT 926.045 1207.175 926.375 1207.190 ;
        RECT 926.965 1207.175 927.295 1207.190 ;
        RECT 925.585 1159.210 925.915 1159.225 ;
        RECT 926.505 1159.210 926.835 1159.225 ;
        RECT 925.585 1158.910 926.835 1159.210 ;
        RECT 925.585 1158.895 925.915 1158.910 ;
        RECT 926.505 1158.895 926.835 1158.910 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 22.000 365.630 22.060 ;
        RECT 932.030 22.000 932.350 22.060 ;
        RECT 365.310 21.860 932.350 22.000 ;
        RECT 365.310 21.800 365.630 21.860 ;
        RECT 932.030 21.800 932.350 21.860 ;
      LAYER via ;
        RECT 365.340 21.800 365.600 22.060 ;
        RECT 932.060 21.800 932.320 22.060 ;
      LAYER met2 ;
        RECT 937.590 1220.330 938.150 1228.680 ;
        RECT 935.340 1220.190 938.150 1220.330 ;
        RECT 935.340 1196.530 935.480 1220.190 ;
        RECT 937.590 1219.680 938.150 1220.190 ;
        RECT 932.120 1196.390 935.480 1196.530 ;
        RECT 932.120 22.090 932.260 1196.390 ;
        RECT 365.340 21.770 365.600 22.090 ;
        RECT 932.060 21.770 932.320 22.090 ;
        RECT 365.400 2.400 365.540 21.770 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 945.370 434.900 945.690 435.160 ;
        RECT 945.460 434.480 945.600 434.900 ;
        RECT 945.370 434.220 945.690 434.480 ;
        RECT 383.250 21.660 383.570 21.720 ;
        RECT 945.370 21.660 945.690 21.720 ;
        RECT 383.250 21.520 945.690 21.660 ;
        RECT 383.250 21.460 383.570 21.520 ;
        RECT 945.370 21.460 945.690 21.520 ;
      LAYER via ;
        RECT 945.400 434.900 945.660 435.160 ;
        RECT 945.400 434.220 945.660 434.480 ;
        RECT 383.280 21.460 383.540 21.720 ;
        RECT 945.400 21.460 945.660 21.720 ;
      LAYER met2 ;
        RECT 946.790 1220.330 947.350 1228.680 ;
        RECT 945.460 1220.190 947.350 1220.330 ;
        RECT 945.460 435.190 945.600 1220.190 ;
        RECT 946.790 1219.680 947.350 1220.190 ;
        RECT 945.400 434.870 945.660 435.190 ;
        RECT 945.400 434.190 945.660 434.510 ;
        RECT 945.460 21.750 945.600 434.190 ;
        RECT 383.280 21.430 383.540 21.750 ;
        RECT 945.400 21.430 945.660 21.750 ;
        RECT 383.340 2.400 383.480 21.430 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 953.725 869.465 953.895 917.575 ;
        RECT 953.265 506.685 953.435 531.335 ;
        RECT 953.265 403.325 953.435 434.775 ;
        RECT 953.265 331.245 953.435 352.495 ;
        RECT 953.265 282.965 953.435 323.255 ;
        RECT 953.265 138.465 953.435 186.235 ;
      LAYER mcon ;
        RECT 953.725 917.405 953.895 917.575 ;
        RECT 953.265 531.165 953.435 531.335 ;
        RECT 953.265 434.605 953.435 434.775 ;
        RECT 953.265 352.325 953.435 352.495 ;
        RECT 953.265 323.085 953.435 323.255 ;
        RECT 953.265 186.065 953.435 186.235 ;
      LAYER met1 ;
        RECT 953.190 1159.300 953.510 1159.360 ;
        RECT 953.650 1159.300 953.970 1159.360 ;
        RECT 953.190 1159.160 953.970 1159.300 ;
        RECT 953.190 1159.100 953.510 1159.160 ;
        RECT 953.650 1159.100 953.970 1159.160 ;
        RECT 953.650 1062.740 953.970 1062.800 ;
        RECT 954.570 1062.740 954.890 1062.800 ;
        RECT 953.650 1062.600 954.890 1062.740 ;
        RECT 953.650 1062.540 953.970 1062.600 ;
        RECT 954.570 1062.540 954.890 1062.600 ;
        RECT 952.270 1014.460 952.590 1014.520 ;
        RECT 953.190 1014.460 953.510 1014.520 ;
        RECT 952.270 1014.320 953.510 1014.460 ;
        RECT 952.270 1014.260 952.590 1014.320 ;
        RECT 953.190 1014.260 953.510 1014.320 ;
        RECT 952.270 966.180 952.590 966.240 ;
        RECT 953.650 966.180 953.970 966.240 ;
        RECT 952.270 966.040 953.970 966.180 ;
        RECT 952.270 965.980 952.590 966.040 ;
        RECT 953.650 965.980 953.970 966.040 ;
        RECT 953.650 917.560 953.970 917.620 ;
        RECT 953.455 917.420 953.970 917.560 ;
        RECT 953.650 917.360 953.970 917.420 ;
        RECT 953.650 869.620 953.970 869.680 ;
        RECT 953.455 869.480 953.970 869.620 ;
        RECT 953.650 869.420 953.970 869.480 ;
        RECT 952.270 814.200 952.590 814.260 ;
        RECT 953.190 814.200 953.510 814.260 ;
        RECT 952.270 814.060 953.510 814.200 ;
        RECT 952.270 814.000 952.590 814.060 ;
        RECT 953.190 814.000 953.510 814.060 ;
        RECT 953.190 724.240 953.510 724.500 ;
        RECT 953.280 724.100 953.420 724.240 ;
        RECT 953.650 724.100 953.970 724.160 ;
        RECT 953.280 723.960 953.970 724.100 ;
        RECT 953.650 723.900 953.970 723.960 ;
        RECT 951.810 717.640 952.130 717.700 ;
        RECT 953.650 717.640 953.970 717.700 ;
        RECT 951.810 717.500 953.970 717.640 ;
        RECT 951.810 717.440 952.130 717.500 ;
        RECT 953.650 717.440 953.970 717.500 ;
        RECT 952.270 669.360 952.590 669.420 ;
        RECT 953.190 669.360 953.510 669.420 ;
        RECT 952.270 669.220 953.510 669.360 ;
        RECT 952.270 669.160 952.590 669.220 ;
        RECT 953.190 669.160 953.510 669.220 ;
        RECT 953.190 620.540 953.510 620.800 ;
        RECT 953.280 620.400 953.420 620.540 ;
        RECT 954.570 620.400 954.890 620.460 ;
        RECT 953.280 620.260 954.890 620.400 ;
        RECT 954.570 620.200 954.890 620.260 ;
        RECT 953.190 531.320 953.510 531.380 ;
        RECT 952.995 531.180 953.510 531.320 ;
        RECT 953.190 531.120 953.510 531.180 ;
        RECT 953.190 506.840 953.510 506.900 ;
        RECT 952.995 506.700 953.510 506.840 ;
        RECT 953.190 506.640 953.510 506.700 ;
        RECT 953.190 458.900 953.510 458.960 ;
        RECT 954.110 458.900 954.430 458.960 ;
        RECT 953.190 458.760 954.430 458.900 ;
        RECT 953.190 458.700 953.510 458.760 ;
        RECT 954.110 458.700 954.430 458.760 ;
        RECT 953.190 434.760 953.510 434.820 ;
        RECT 952.995 434.620 953.510 434.760 ;
        RECT 953.190 434.560 953.510 434.620 ;
        RECT 953.190 403.480 953.510 403.540 ;
        RECT 952.995 403.340 953.510 403.480 ;
        RECT 953.190 403.280 953.510 403.340 ;
        RECT 953.190 352.480 953.510 352.540 ;
        RECT 952.995 352.340 953.510 352.480 ;
        RECT 953.190 352.280 953.510 352.340 ;
        RECT 953.190 331.400 953.510 331.460 ;
        RECT 952.995 331.260 953.510 331.400 ;
        RECT 953.190 331.200 953.510 331.260 ;
        RECT 953.190 323.240 953.510 323.300 ;
        RECT 952.995 323.100 953.510 323.240 ;
        RECT 953.190 323.040 953.510 323.100 ;
        RECT 953.205 283.120 953.495 283.165 ;
        RECT 953.650 283.120 953.970 283.180 ;
        RECT 953.205 282.980 953.970 283.120 ;
        RECT 953.205 282.935 953.495 282.980 ;
        RECT 953.650 282.920 953.970 282.980 ;
        RECT 953.190 241.640 953.510 241.700 ;
        RECT 953.650 241.640 953.970 241.700 ;
        RECT 953.190 241.500 953.970 241.640 ;
        RECT 953.190 241.440 953.510 241.500 ;
        RECT 953.650 241.440 953.970 241.500 ;
        RECT 953.190 193.360 953.510 193.420 ;
        RECT 953.650 193.360 953.970 193.420 ;
        RECT 953.190 193.220 953.970 193.360 ;
        RECT 953.190 193.160 953.510 193.220 ;
        RECT 953.650 193.160 953.970 193.220 ;
        RECT 953.205 186.220 953.495 186.265 ;
        RECT 953.650 186.220 953.970 186.280 ;
        RECT 953.205 186.080 953.970 186.220 ;
        RECT 953.205 186.035 953.495 186.080 ;
        RECT 953.650 186.020 953.970 186.080 ;
        RECT 953.190 138.620 953.510 138.680 ;
        RECT 952.995 138.480 953.510 138.620 ;
        RECT 953.190 138.420 953.510 138.480 ;
        RECT 953.190 110.540 953.510 110.800 ;
        RECT 953.280 110.060 953.420 110.540 ;
        RECT 953.650 110.060 953.970 110.120 ;
        RECT 953.280 109.920 953.970 110.060 ;
        RECT 953.650 109.860 953.970 109.920 ;
        RECT 952.270 67.560 952.590 67.620 ;
        RECT 953.650 67.560 953.970 67.620 ;
        RECT 952.270 67.420 953.970 67.560 ;
        RECT 952.270 67.360 952.590 67.420 ;
        RECT 953.650 67.360 953.970 67.420 ;
        RECT 401.190 21.320 401.510 21.380 ;
        RECT 952.270 21.320 952.590 21.380 ;
        RECT 401.190 21.180 952.590 21.320 ;
        RECT 401.190 21.120 401.510 21.180 ;
        RECT 952.270 21.120 952.590 21.180 ;
      LAYER via ;
        RECT 953.220 1159.100 953.480 1159.360 ;
        RECT 953.680 1159.100 953.940 1159.360 ;
        RECT 953.680 1062.540 953.940 1062.800 ;
        RECT 954.600 1062.540 954.860 1062.800 ;
        RECT 952.300 1014.260 952.560 1014.520 ;
        RECT 953.220 1014.260 953.480 1014.520 ;
        RECT 952.300 965.980 952.560 966.240 ;
        RECT 953.680 965.980 953.940 966.240 ;
        RECT 953.680 917.360 953.940 917.620 ;
        RECT 953.680 869.420 953.940 869.680 ;
        RECT 952.300 814.000 952.560 814.260 ;
        RECT 953.220 814.000 953.480 814.260 ;
        RECT 953.220 724.240 953.480 724.500 ;
        RECT 953.680 723.900 953.940 724.160 ;
        RECT 951.840 717.440 952.100 717.700 ;
        RECT 953.680 717.440 953.940 717.700 ;
        RECT 952.300 669.160 952.560 669.420 ;
        RECT 953.220 669.160 953.480 669.420 ;
        RECT 953.220 620.540 953.480 620.800 ;
        RECT 954.600 620.200 954.860 620.460 ;
        RECT 953.220 531.120 953.480 531.380 ;
        RECT 953.220 506.640 953.480 506.900 ;
        RECT 953.220 458.700 953.480 458.960 ;
        RECT 954.140 458.700 954.400 458.960 ;
        RECT 953.220 434.560 953.480 434.820 ;
        RECT 953.220 403.280 953.480 403.540 ;
        RECT 953.220 352.280 953.480 352.540 ;
        RECT 953.220 331.200 953.480 331.460 ;
        RECT 953.220 323.040 953.480 323.300 ;
        RECT 953.680 282.920 953.940 283.180 ;
        RECT 953.220 241.440 953.480 241.700 ;
        RECT 953.680 241.440 953.940 241.700 ;
        RECT 953.220 193.160 953.480 193.420 ;
        RECT 953.680 193.160 953.940 193.420 ;
        RECT 953.680 186.020 953.940 186.280 ;
        RECT 953.220 138.420 953.480 138.680 ;
        RECT 953.220 110.540 953.480 110.800 ;
        RECT 953.680 109.860 953.940 110.120 ;
        RECT 952.300 67.360 952.560 67.620 ;
        RECT 953.680 67.360 953.940 67.620 ;
        RECT 401.220 21.120 401.480 21.380 ;
        RECT 952.300 21.120 952.560 21.380 ;
      LAYER met2 ;
        RECT 955.530 1221.010 956.090 1228.680 ;
        RECT 953.740 1220.870 956.090 1221.010 ;
        RECT 953.740 1159.390 953.880 1220.870 ;
        RECT 955.530 1219.680 956.090 1220.870 ;
        RECT 953.220 1159.070 953.480 1159.390 ;
        RECT 953.680 1159.070 953.940 1159.390 ;
        RECT 953.280 1124.450 953.420 1159.070 ;
        RECT 953.280 1124.310 953.880 1124.450 ;
        RECT 953.740 1110.965 953.880 1124.310 ;
        RECT 953.670 1110.595 953.950 1110.965 ;
        RECT 954.590 1110.595 954.870 1110.965 ;
        RECT 954.660 1062.830 954.800 1110.595 ;
        RECT 953.680 1062.685 953.940 1062.830 ;
        RECT 952.290 1062.315 952.570 1062.685 ;
        RECT 953.670 1062.315 953.950 1062.685 ;
        RECT 954.600 1062.510 954.860 1062.830 ;
        RECT 952.360 1014.550 952.500 1062.315 ;
        RECT 952.300 1014.405 952.560 1014.550 ;
        RECT 953.220 1014.405 953.480 1014.550 ;
        RECT 952.290 1014.035 952.570 1014.405 ;
        RECT 953.210 1014.035 953.490 1014.405 ;
        RECT 952.360 966.270 952.500 1014.035 ;
        RECT 952.300 965.950 952.560 966.270 ;
        RECT 953.680 966.125 953.940 966.270 ;
        RECT 953.670 965.755 953.950 966.125 ;
        RECT 954.590 965.755 954.870 966.125 ;
        RECT 954.660 930.650 954.800 965.755 ;
        RECT 953.740 930.510 954.800 930.650 ;
        RECT 953.740 917.650 953.880 930.510 ;
        RECT 953.680 917.330 953.940 917.650 ;
        RECT 953.680 869.390 953.940 869.710 ;
        RECT 953.740 845.650 953.880 869.390 ;
        RECT 953.280 845.510 953.880 845.650 ;
        RECT 953.280 814.290 953.420 845.510 ;
        RECT 952.300 813.970 952.560 814.290 ;
        RECT 953.220 813.970 953.480 814.290 ;
        RECT 952.360 766.205 952.500 813.970 ;
        RECT 952.290 765.835 952.570 766.205 ;
        RECT 953.670 765.835 953.950 766.205 ;
        RECT 953.740 724.610 953.880 765.835 ;
        RECT 953.280 724.530 953.880 724.610 ;
        RECT 953.220 724.470 953.880 724.530 ;
        RECT 953.220 724.210 953.480 724.470 ;
        RECT 953.680 723.870 953.940 724.190 ;
        RECT 953.740 717.730 953.880 723.870 ;
        RECT 951.840 717.410 952.100 717.730 ;
        RECT 953.680 717.410 953.940 717.730 ;
        RECT 951.900 669.645 952.040 717.410 ;
        RECT 951.830 669.275 952.110 669.645 ;
        RECT 952.300 669.130 952.560 669.450 ;
        RECT 953.210 669.275 953.490 669.645 ;
        RECT 953.220 669.130 953.480 669.275 ;
        RECT 952.360 621.365 952.500 669.130 ;
        RECT 952.290 620.995 952.570 621.365 ;
        RECT 953.210 620.995 953.490 621.365 ;
        RECT 953.280 620.830 953.420 620.995 ;
        RECT 953.220 620.510 953.480 620.830 ;
        RECT 954.600 620.170 954.860 620.490 ;
        RECT 954.660 579.090 954.800 620.170 ;
        RECT 954.200 578.950 954.800 579.090 ;
        RECT 954.200 531.605 954.340 578.950 ;
        RECT 953.210 531.235 953.490 531.605 ;
        RECT 954.130 531.235 954.410 531.605 ;
        RECT 953.220 531.090 953.480 531.235 ;
        RECT 953.220 506.610 953.480 506.930 ;
        RECT 953.280 458.990 953.420 506.610 ;
        RECT 953.220 458.670 953.480 458.990 ;
        RECT 954.140 458.670 954.400 458.990 ;
        RECT 954.200 435.045 954.340 458.670 ;
        RECT 953.210 434.675 953.490 435.045 ;
        RECT 954.130 434.675 954.410 435.045 ;
        RECT 953.220 434.530 953.480 434.675 ;
        RECT 953.220 403.250 953.480 403.570 ;
        RECT 953.280 352.570 953.420 403.250 ;
        RECT 953.220 352.250 953.480 352.570 ;
        RECT 953.220 331.170 953.480 331.490 ;
        RECT 953.280 323.330 953.420 331.170 ;
        RECT 953.220 323.010 953.480 323.330 ;
        RECT 953.680 282.890 953.940 283.210 ;
        RECT 953.740 241.730 953.880 282.890 ;
        RECT 953.220 241.410 953.480 241.730 ;
        RECT 953.680 241.410 953.940 241.730 ;
        RECT 953.280 193.450 953.420 241.410 ;
        RECT 953.220 193.130 953.480 193.450 ;
        RECT 953.680 193.130 953.940 193.450 ;
        RECT 953.740 186.310 953.880 193.130 ;
        RECT 953.680 185.990 953.940 186.310 ;
        RECT 953.220 138.390 953.480 138.710 ;
        RECT 953.280 110.830 953.420 138.390 ;
        RECT 953.220 110.510 953.480 110.830 ;
        RECT 953.680 109.830 953.940 110.150 ;
        RECT 953.740 67.650 953.880 109.830 ;
        RECT 952.300 67.330 952.560 67.650 ;
        RECT 953.680 67.330 953.940 67.650 ;
        RECT 952.360 21.410 952.500 67.330 ;
        RECT 401.220 21.090 401.480 21.410 ;
        RECT 952.300 21.090 952.560 21.410 ;
        RECT 401.280 2.400 401.420 21.090 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 953.670 1110.640 953.950 1110.920 ;
        RECT 954.590 1110.640 954.870 1110.920 ;
        RECT 952.290 1062.360 952.570 1062.640 ;
        RECT 953.670 1062.360 953.950 1062.640 ;
        RECT 952.290 1014.080 952.570 1014.360 ;
        RECT 953.210 1014.080 953.490 1014.360 ;
        RECT 953.670 965.800 953.950 966.080 ;
        RECT 954.590 965.800 954.870 966.080 ;
        RECT 952.290 765.880 952.570 766.160 ;
        RECT 953.670 765.880 953.950 766.160 ;
        RECT 951.830 669.320 952.110 669.600 ;
        RECT 953.210 669.320 953.490 669.600 ;
        RECT 952.290 621.040 952.570 621.320 ;
        RECT 953.210 621.040 953.490 621.320 ;
        RECT 953.210 531.280 953.490 531.560 ;
        RECT 954.130 531.280 954.410 531.560 ;
        RECT 953.210 434.720 953.490 435.000 ;
        RECT 954.130 434.720 954.410 435.000 ;
      LAYER met3 ;
        RECT 953.645 1110.930 953.975 1110.945 ;
        RECT 954.565 1110.930 954.895 1110.945 ;
        RECT 953.645 1110.630 954.895 1110.930 ;
        RECT 953.645 1110.615 953.975 1110.630 ;
        RECT 954.565 1110.615 954.895 1110.630 ;
        RECT 952.265 1062.650 952.595 1062.665 ;
        RECT 953.645 1062.650 953.975 1062.665 ;
        RECT 952.265 1062.350 953.975 1062.650 ;
        RECT 952.265 1062.335 952.595 1062.350 ;
        RECT 953.645 1062.335 953.975 1062.350 ;
        RECT 952.265 1014.370 952.595 1014.385 ;
        RECT 953.185 1014.370 953.515 1014.385 ;
        RECT 952.265 1014.070 953.515 1014.370 ;
        RECT 952.265 1014.055 952.595 1014.070 ;
        RECT 953.185 1014.055 953.515 1014.070 ;
        RECT 953.645 966.090 953.975 966.105 ;
        RECT 954.565 966.090 954.895 966.105 ;
        RECT 953.645 965.790 954.895 966.090 ;
        RECT 953.645 965.775 953.975 965.790 ;
        RECT 954.565 965.775 954.895 965.790 ;
        RECT 952.265 766.170 952.595 766.185 ;
        RECT 953.645 766.170 953.975 766.185 ;
        RECT 952.265 765.870 953.975 766.170 ;
        RECT 952.265 765.855 952.595 765.870 ;
        RECT 953.645 765.855 953.975 765.870 ;
        RECT 951.805 669.610 952.135 669.625 ;
        RECT 953.185 669.610 953.515 669.625 ;
        RECT 951.805 669.310 953.515 669.610 ;
        RECT 951.805 669.295 952.135 669.310 ;
        RECT 953.185 669.295 953.515 669.310 ;
        RECT 952.265 621.330 952.595 621.345 ;
        RECT 953.185 621.330 953.515 621.345 ;
        RECT 952.265 621.030 953.515 621.330 ;
        RECT 952.265 621.015 952.595 621.030 ;
        RECT 953.185 621.015 953.515 621.030 ;
        RECT 953.185 531.570 953.515 531.585 ;
        RECT 954.105 531.570 954.435 531.585 ;
        RECT 953.185 531.270 954.435 531.570 ;
        RECT 953.185 531.255 953.515 531.270 ;
        RECT 954.105 531.255 954.435 531.270 ;
        RECT 953.185 435.010 953.515 435.025 ;
        RECT 954.105 435.010 954.435 435.025 ;
        RECT 953.185 434.710 954.435 435.010 ;
        RECT 953.185 434.695 953.515 434.710 ;
        RECT 954.105 434.695 954.435 434.710 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.650 1220.330 782.210 1228.680 ;
        RECT 779.860 1220.190 782.210 1220.330 ;
        RECT 779.860 24.325 780.000 1220.190 ;
        RECT 781.650 1219.680 782.210 1220.190 ;
        RECT 62.190 23.955 62.470 24.325 ;
        RECT 779.790 23.955 780.070 24.325 ;
        RECT 62.260 2.400 62.400 23.955 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 62.190 24.000 62.470 24.280 ;
        RECT 779.790 24.000 780.070 24.280 ;
      LAYER met3 ;
        RECT 62.165 24.290 62.495 24.305 ;
        RECT 779.765 24.290 780.095 24.305 ;
        RECT 62.165 23.990 780.095 24.290 ;
        RECT 62.165 23.975 62.495 23.990 ;
        RECT 779.765 23.975 780.095 23.990 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 959.705 1110.865 959.875 1124.975 ;
        RECT 960.165 869.465 960.335 917.235 ;
        RECT 960.165 620.585 960.335 662.235 ;
        RECT 959.705 559.045 959.875 566.355 ;
        RECT 959.705 379.525 959.875 434.775 ;
        RECT 960.165 269.025 960.335 276.675 ;
        RECT 959.705 131.325 959.875 138.295 ;
        RECT 959.705 48.365 959.875 107.015 ;
      LAYER mcon ;
        RECT 959.705 1124.805 959.875 1124.975 ;
        RECT 960.165 917.065 960.335 917.235 ;
        RECT 960.165 662.065 960.335 662.235 ;
        RECT 959.705 566.185 959.875 566.355 ;
        RECT 959.705 434.605 959.875 434.775 ;
        RECT 960.165 276.505 960.335 276.675 ;
        RECT 959.705 138.125 959.875 138.295 ;
        RECT 959.705 106.845 959.875 107.015 ;
      LAYER met1 ;
        RECT 959.630 1124.960 959.950 1125.020 ;
        RECT 959.435 1124.820 959.950 1124.960 ;
        RECT 959.630 1124.760 959.950 1124.820 ;
        RECT 959.630 1111.020 959.950 1111.080 ;
        RECT 959.435 1110.880 959.950 1111.020 ;
        RECT 959.630 1110.820 959.950 1110.880 ;
        RECT 958.710 1062.740 959.030 1062.800 ;
        RECT 960.090 1062.740 960.410 1062.800 ;
        RECT 958.710 1062.600 960.410 1062.740 ;
        RECT 958.710 1062.540 959.030 1062.600 ;
        RECT 960.090 1062.540 960.410 1062.600 ;
        RECT 960.090 1028.540 960.410 1028.800 ;
        RECT 960.180 1028.120 960.320 1028.540 ;
        RECT 960.090 1027.860 960.410 1028.120 ;
        RECT 959.170 966.180 959.490 966.240 ;
        RECT 960.090 966.180 960.410 966.240 ;
        RECT 959.170 966.040 960.410 966.180 ;
        RECT 959.170 965.980 959.490 966.040 ;
        RECT 960.090 965.980 960.410 966.040 ;
        RECT 960.090 917.220 960.410 917.280 ;
        RECT 959.895 917.080 960.410 917.220 ;
        RECT 960.090 917.020 960.410 917.080 ;
        RECT 960.090 869.620 960.410 869.680 ;
        RECT 959.895 869.480 960.410 869.620 ;
        RECT 960.090 869.420 960.410 869.480 ;
        RECT 959.170 724.440 959.490 724.500 ;
        RECT 959.630 724.440 959.950 724.500 ;
        RECT 959.170 724.300 959.950 724.440 ;
        RECT 959.170 724.240 959.490 724.300 ;
        RECT 959.630 724.240 959.950 724.300 ;
        RECT 960.090 662.220 960.410 662.280 ;
        RECT 959.895 662.080 960.410 662.220 ;
        RECT 960.090 662.020 960.410 662.080 ;
        RECT 960.090 620.740 960.410 620.800 ;
        RECT 959.895 620.600 960.410 620.740 ;
        RECT 960.090 620.540 960.410 620.600 ;
        RECT 959.645 566.340 959.935 566.385 ;
        RECT 960.090 566.340 960.410 566.400 ;
        RECT 959.645 566.200 960.410 566.340 ;
        RECT 959.645 566.155 959.935 566.200 ;
        RECT 960.090 566.140 960.410 566.200 ;
        RECT 959.630 559.200 959.950 559.260 ;
        RECT 959.435 559.060 959.950 559.200 ;
        RECT 959.630 559.000 959.950 559.060 ;
        RECT 958.710 510.920 959.030 510.980 ;
        RECT 961.010 510.920 961.330 510.980 ;
        RECT 958.710 510.780 961.330 510.920 ;
        RECT 958.710 510.720 959.030 510.780 ;
        RECT 961.010 510.720 961.330 510.780 ;
        RECT 960.090 462.640 960.410 462.700 ;
        RECT 960.550 462.640 960.870 462.700 ;
        RECT 960.090 462.500 960.870 462.640 ;
        RECT 960.090 462.440 960.410 462.500 ;
        RECT 960.550 462.440 960.870 462.500 ;
        RECT 959.630 434.760 959.950 434.820 ;
        RECT 959.435 434.620 959.950 434.760 ;
        RECT 959.630 434.560 959.950 434.620 ;
        RECT 959.645 379.680 959.935 379.725 ;
        RECT 960.090 379.680 960.410 379.740 ;
        RECT 959.645 379.540 960.410 379.680 ;
        RECT 959.645 379.495 959.935 379.540 ;
        RECT 960.090 379.480 960.410 379.540 ;
        RECT 960.090 352.480 960.410 352.540 ;
        RECT 959.720 352.340 960.410 352.480 ;
        RECT 959.720 351.860 959.860 352.340 ;
        RECT 960.090 352.280 960.410 352.340 ;
        RECT 959.630 351.600 959.950 351.860 ;
        RECT 959.630 331.060 959.950 331.120 ;
        RECT 960.550 331.060 960.870 331.120 ;
        RECT 959.630 330.920 960.870 331.060 ;
        RECT 959.630 330.860 959.950 330.920 ;
        RECT 960.550 330.860 960.870 330.920 ;
        RECT 960.105 276.660 960.395 276.705 ;
        RECT 960.550 276.660 960.870 276.720 ;
        RECT 960.105 276.520 960.870 276.660 ;
        RECT 960.105 276.475 960.395 276.520 ;
        RECT 960.550 276.460 960.870 276.520 ;
        RECT 960.090 269.180 960.410 269.240 ;
        RECT 959.895 269.040 960.410 269.180 ;
        RECT 960.090 268.980 960.410 269.040 ;
        RECT 959.630 138.280 959.950 138.340 ;
        RECT 959.435 138.140 959.950 138.280 ;
        RECT 959.630 138.080 959.950 138.140 ;
        RECT 959.630 131.480 959.950 131.540 ;
        RECT 959.435 131.340 959.950 131.480 ;
        RECT 959.630 131.280 959.950 131.340 ;
        RECT 958.710 107.000 959.030 107.060 ;
        RECT 959.645 107.000 959.935 107.045 ;
        RECT 958.710 106.860 959.935 107.000 ;
        RECT 958.710 106.800 959.030 106.860 ;
        RECT 959.645 106.815 959.935 106.860 ;
        RECT 959.630 48.520 959.950 48.580 ;
        RECT 959.435 48.380 959.950 48.520 ;
        RECT 959.630 48.320 959.950 48.380 ;
        RECT 419.130 20.980 419.450 21.040 ;
        RECT 959.170 20.980 959.490 21.040 ;
        RECT 419.130 20.840 959.490 20.980 ;
        RECT 419.130 20.780 419.450 20.840 ;
        RECT 959.170 20.780 959.490 20.840 ;
      LAYER via ;
        RECT 959.660 1124.760 959.920 1125.020 ;
        RECT 959.660 1110.820 959.920 1111.080 ;
        RECT 958.740 1062.540 959.000 1062.800 ;
        RECT 960.120 1062.540 960.380 1062.800 ;
        RECT 960.120 1028.540 960.380 1028.800 ;
        RECT 960.120 1027.860 960.380 1028.120 ;
        RECT 959.200 965.980 959.460 966.240 ;
        RECT 960.120 965.980 960.380 966.240 ;
        RECT 960.120 917.020 960.380 917.280 ;
        RECT 960.120 869.420 960.380 869.680 ;
        RECT 959.200 724.240 959.460 724.500 ;
        RECT 959.660 724.240 959.920 724.500 ;
        RECT 960.120 662.020 960.380 662.280 ;
        RECT 960.120 620.540 960.380 620.800 ;
        RECT 960.120 566.140 960.380 566.400 ;
        RECT 959.660 559.000 959.920 559.260 ;
        RECT 958.740 510.720 959.000 510.980 ;
        RECT 961.040 510.720 961.300 510.980 ;
        RECT 960.120 462.440 960.380 462.700 ;
        RECT 960.580 462.440 960.840 462.700 ;
        RECT 959.660 434.560 959.920 434.820 ;
        RECT 960.120 379.480 960.380 379.740 ;
        RECT 960.120 352.280 960.380 352.540 ;
        RECT 959.660 351.600 959.920 351.860 ;
        RECT 959.660 330.860 959.920 331.120 ;
        RECT 960.580 330.860 960.840 331.120 ;
        RECT 960.580 276.460 960.840 276.720 ;
        RECT 960.120 268.980 960.380 269.240 ;
        RECT 959.660 138.080 959.920 138.340 ;
        RECT 959.660 131.280 959.920 131.540 ;
        RECT 958.740 106.800 959.000 107.060 ;
        RECT 959.660 48.320 959.920 48.580 ;
        RECT 419.160 20.780 419.420 21.040 ;
        RECT 959.200 20.780 959.460 21.040 ;
      LAYER met2 ;
        RECT 964.730 1221.010 965.290 1228.680 ;
        RECT 962.940 1220.870 965.290 1221.010 ;
        RECT 962.940 1196.530 963.080 1220.870 ;
        RECT 964.730 1219.680 965.290 1220.870 ;
        RECT 960.180 1196.390 963.080 1196.530 ;
        RECT 960.180 1159.130 960.320 1196.390 ;
        RECT 959.720 1158.990 960.320 1159.130 ;
        RECT 959.720 1125.050 959.860 1158.990 ;
        RECT 959.660 1124.730 959.920 1125.050 ;
        RECT 959.660 1110.965 959.920 1111.110 ;
        RECT 958.730 1110.595 959.010 1110.965 ;
        RECT 959.650 1110.595 959.930 1110.965 ;
        RECT 958.800 1062.830 958.940 1110.595 ;
        RECT 958.740 1062.510 959.000 1062.830 ;
        RECT 960.120 1062.510 960.380 1062.830 ;
        RECT 960.180 1028.830 960.320 1062.510 ;
        RECT 960.120 1028.510 960.380 1028.830 ;
        RECT 960.120 1027.830 960.380 1028.150 ;
        RECT 960.180 1015.085 960.320 1027.830 ;
        RECT 960.110 1014.715 960.390 1015.085 ;
        RECT 959.190 1014.035 959.470 1014.405 ;
        RECT 959.260 966.270 959.400 1014.035 ;
        RECT 959.200 965.950 959.460 966.270 ;
        RECT 960.120 966.125 960.380 966.270 ;
        RECT 960.110 965.755 960.390 966.125 ;
        RECT 961.030 965.755 961.310 966.125 ;
        RECT 961.100 930.650 961.240 965.755 ;
        RECT 960.180 930.510 961.240 930.650 ;
        RECT 960.180 917.310 960.320 930.510 ;
        RECT 960.120 916.990 960.380 917.310 ;
        RECT 960.120 869.390 960.380 869.710 ;
        RECT 960.180 814.485 960.320 869.390 ;
        RECT 960.110 814.115 960.390 814.485 ;
        RECT 960.570 813.435 960.850 813.805 ;
        RECT 960.640 724.725 960.780 813.435 ;
        RECT 959.200 724.210 959.460 724.530 ;
        RECT 959.650 724.355 959.930 724.725 ;
        RECT 960.570 724.355 960.850 724.725 ;
        RECT 959.660 724.210 959.920 724.355 ;
        RECT 959.260 676.445 959.400 724.210 ;
        RECT 959.190 676.075 959.470 676.445 ;
        RECT 960.110 676.075 960.390 676.445 ;
        RECT 960.180 662.310 960.320 676.075 ;
        RECT 960.120 661.990 960.380 662.310 ;
        RECT 960.120 620.510 960.380 620.830 ;
        RECT 960.180 566.430 960.320 620.510 ;
        RECT 960.120 566.110 960.380 566.430 ;
        RECT 959.660 558.970 959.920 559.290 ;
        RECT 959.720 558.805 959.860 558.970 ;
        RECT 958.730 558.435 959.010 558.805 ;
        RECT 959.650 558.435 959.930 558.805 ;
        RECT 958.800 511.010 958.940 558.435 ;
        RECT 958.740 510.690 959.000 511.010 ;
        RECT 961.040 510.690 961.300 511.010 ;
        RECT 961.100 496.130 961.240 510.690 ;
        RECT 960.640 495.990 961.240 496.130 ;
        RECT 960.640 462.730 960.780 495.990 ;
        RECT 960.120 462.410 960.380 462.730 ;
        RECT 960.580 462.410 960.840 462.730 ;
        RECT 960.180 458.050 960.320 462.410 ;
        RECT 959.720 457.910 960.320 458.050 ;
        RECT 959.720 434.850 959.860 457.910 ;
        RECT 959.660 434.530 959.920 434.850 ;
        RECT 960.120 379.450 960.380 379.770 ;
        RECT 960.180 352.570 960.320 379.450 ;
        RECT 960.120 352.250 960.380 352.570 ;
        RECT 959.660 351.570 959.920 351.890 ;
        RECT 959.720 331.150 959.860 351.570 ;
        RECT 959.660 330.830 959.920 331.150 ;
        RECT 960.580 330.830 960.840 331.150 ;
        RECT 960.640 276.750 960.780 330.830 ;
        RECT 960.580 276.430 960.840 276.750 ;
        RECT 960.120 268.950 960.380 269.270 ;
        RECT 960.180 229.570 960.320 268.950 ;
        RECT 959.720 229.430 960.320 229.570 ;
        RECT 959.720 220.845 959.860 229.430 ;
        RECT 959.650 220.475 959.930 220.845 ;
        RECT 960.570 220.475 960.850 220.845 ;
        RECT 960.640 178.570 960.780 220.475 ;
        RECT 959.720 178.430 960.780 178.570 ;
        RECT 959.720 138.370 959.860 178.430 ;
        RECT 959.660 138.050 959.920 138.370 ;
        RECT 959.660 131.250 959.920 131.570 ;
        RECT 959.720 131.085 959.860 131.250 ;
        RECT 958.730 130.715 959.010 131.085 ;
        RECT 959.650 130.715 959.930 131.085 ;
        RECT 958.800 107.090 958.940 130.715 ;
        RECT 958.740 106.770 959.000 107.090 ;
        RECT 959.660 48.290 959.920 48.610 ;
        RECT 959.720 48.010 959.860 48.290 ;
        RECT 959.260 47.870 959.860 48.010 ;
        RECT 959.260 21.070 959.400 47.870 ;
        RECT 419.160 20.750 419.420 21.070 ;
        RECT 959.200 20.750 959.460 21.070 ;
        RECT 419.220 2.400 419.360 20.750 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 958.730 1110.640 959.010 1110.920 ;
        RECT 959.650 1110.640 959.930 1110.920 ;
        RECT 960.110 1014.760 960.390 1015.040 ;
        RECT 959.190 1014.080 959.470 1014.360 ;
        RECT 960.110 965.800 960.390 966.080 ;
        RECT 961.030 965.800 961.310 966.080 ;
        RECT 960.110 814.160 960.390 814.440 ;
        RECT 960.570 813.480 960.850 813.760 ;
        RECT 959.650 724.400 959.930 724.680 ;
        RECT 960.570 724.400 960.850 724.680 ;
        RECT 959.190 676.120 959.470 676.400 ;
        RECT 960.110 676.120 960.390 676.400 ;
        RECT 958.730 558.480 959.010 558.760 ;
        RECT 959.650 558.480 959.930 558.760 ;
        RECT 959.650 220.520 959.930 220.800 ;
        RECT 960.570 220.520 960.850 220.800 ;
        RECT 958.730 130.760 959.010 131.040 ;
        RECT 959.650 130.760 959.930 131.040 ;
      LAYER met3 ;
        RECT 958.705 1110.930 959.035 1110.945 ;
        RECT 959.625 1110.930 959.955 1110.945 ;
        RECT 958.705 1110.630 959.955 1110.930 ;
        RECT 958.705 1110.615 959.035 1110.630 ;
        RECT 959.625 1110.615 959.955 1110.630 ;
        RECT 960.085 1015.050 960.415 1015.065 ;
        RECT 959.870 1014.735 960.415 1015.050 ;
        RECT 959.165 1014.370 959.495 1014.385 ;
        RECT 959.870 1014.370 960.170 1014.735 ;
        RECT 959.165 1014.070 960.170 1014.370 ;
        RECT 959.165 1014.055 959.495 1014.070 ;
        RECT 960.085 966.090 960.415 966.105 ;
        RECT 961.005 966.090 961.335 966.105 ;
        RECT 960.085 965.790 961.335 966.090 ;
        RECT 960.085 965.775 960.415 965.790 ;
        RECT 961.005 965.775 961.335 965.790 ;
        RECT 960.085 814.450 960.415 814.465 ;
        RECT 959.870 814.135 960.415 814.450 ;
        RECT 959.870 813.770 960.170 814.135 ;
        RECT 960.545 813.770 960.875 813.785 ;
        RECT 959.870 813.470 960.875 813.770 ;
        RECT 960.545 813.455 960.875 813.470 ;
        RECT 959.625 724.690 959.955 724.705 ;
        RECT 960.545 724.690 960.875 724.705 ;
        RECT 959.625 724.390 960.875 724.690 ;
        RECT 959.625 724.375 959.955 724.390 ;
        RECT 960.545 724.375 960.875 724.390 ;
        RECT 959.165 676.410 959.495 676.425 ;
        RECT 960.085 676.410 960.415 676.425 ;
        RECT 959.165 676.110 960.415 676.410 ;
        RECT 959.165 676.095 959.495 676.110 ;
        RECT 960.085 676.095 960.415 676.110 ;
        RECT 958.705 558.770 959.035 558.785 ;
        RECT 959.625 558.770 959.955 558.785 ;
        RECT 958.705 558.470 959.955 558.770 ;
        RECT 958.705 558.455 959.035 558.470 ;
        RECT 959.625 558.455 959.955 558.470 ;
        RECT 959.625 220.810 959.955 220.825 ;
        RECT 960.545 220.810 960.875 220.825 ;
        RECT 959.625 220.510 960.875 220.810 ;
        RECT 959.625 220.495 959.955 220.510 ;
        RECT 960.545 220.495 960.875 220.510 ;
        RECT 958.705 131.050 959.035 131.065 ;
        RECT 959.625 131.050 959.955 131.065 ;
        RECT 958.705 130.750 959.955 131.050 ;
        RECT 958.705 130.735 959.035 130.750 ;
        RECT 959.625 130.735 959.955 130.750 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 38.320 436.930 38.380 ;
        RECT 972.970 38.320 973.290 38.380 ;
        RECT 436.610 38.180 973.290 38.320 ;
        RECT 436.610 38.120 436.930 38.180 ;
        RECT 972.970 38.120 973.290 38.180 ;
      LAYER via ;
        RECT 436.640 38.120 436.900 38.380 ;
        RECT 973.000 38.120 973.260 38.380 ;
      LAYER met2 ;
        RECT 973.930 1220.330 974.490 1228.680 ;
        RECT 973.060 1220.190 974.490 1220.330 ;
        RECT 973.060 38.410 973.200 1220.190 ;
        RECT 973.930 1219.680 974.490 1220.190 ;
        RECT 436.640 38.090 436.900 38.410 ;
        RECT 973.000 38.090 973.260 38.410 ;
        RECT 436.700 2.400 436.840 38.090 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 981.325 897.005 981.495 945.115 ;
      LAYER mcon ;
        RECT 981.325 944.945 981.495 945.115 ;
      LAYER met1 ;
        RECT 980.790 1159.300 981.110 1159.360 ;
        RECT 981.250 1159.300 981.570 1159.360 ;
        RECT 980.790 1159.160 981.570 1159.300 ;
        RECT 980.790 1159.100 981.110 1159.160 ;
        RECT 981.250 1159.100 981.570 1159.160 ;
        RECT 980.790 1111.020 981.110 1111.080 ;
        RECT 981.710 1111.020 982.030 1111.080 ;
        RECT 980.790 1110.880 982.030 1111.020 ;
        RECT 980.790 1110.820 981.110 1110.880 ;
        RECT 981.710 1110.820 982.030 1110.880 ;
        RECT 981.250 1056.280 981.570 1056.340 ;
        RECT 981.710 1056.280 982.030 1056.340 ;
        RECT 981.250 1056.140 982.030 1056.280 ;
        RECT 981.250 1056.080 981.570 1056.140 ;
        RECT 981.710 1056.080 982.030 1056.140 ;
        RECT 979.870 1008.000 980.190 1008.060 ;
        RECT 981.250 1008.000 981.570 1008.060 ;
        RECT 979.870 1007.860 981.570 1008.000 ;
        RECT 979.870 1007.800 980.190 1007.860 ;
        RECT 981.250 1007.800 981.570 1007.860 ;
        RECT 981.265 945.100 981.555 945.145 ;
        RECT 981.710 945.100 982.030 945.160 ;
        RECT 981.265 944.960 982.030 945.100 ;
        RECT 981.265 944.915 981.555 944.960 ;
        RECT 981.710 944.900 982.030 944.960 ;
        RECT 981.250 897.160 981.570 897.220 ;
        RECT 981.055 897.020 981.570 897.160 ;
        RECT 981.250 896.960 981.570 897.020 ;
        RECT 981.250 814.340 981.570 814.600 ;
        RECT 981.340 813.920 981.480 814.340 ;
        RECT 981.250 813.660 981.570 813.920 ;
        RECT 981.250 711.180 981.570 711.240 ;
        RECT 980.880 711.040 981.570 711.180 ;
        RECT 980.880 710.560 981.020 711.040 ;
        RECT 981.250 710.980 981.570 711.040 ;
        RECT 980.790 710.300 981.110 710.560 ;
        RECT 980.790 614.280 981.110 614.340 ;
        RECT 981.250 614.280 981.570 614.340 ;
        RECT 980.790 614.140 981.570 614.280 ;
        RECT 980.790 614.080 981.110 614.140 ;
        RECT 981.250 614.080 981.570 614.140 ;
        RECT 980.790 566.000 981.110 566.060 ;
        RECT 981.250 566.000 981.570 566.060 ;
        RECT 980.790 565.860 981.570 566.000 ;
        RECT 980.790 565.800 981.110 565.860 ;
        RECT 981.250 565.800 981.570 565.860 ;
        RECT 981.250 379.340 981.570 379.400 ;
        RECT 981.710 379.340 982.030 379.400 ;
        RECT 981.250 379.200 982.030 379.340 ;
        RECT 981.250 379.140 981.570 379.200 ;
        RECT 981.710 379.140 982.030 379.200 ;
        RECT 981.250 255.580 981.570 255.640 ;
        RECT 980.880 255.440 981.570 255.580 ;
        RECT 980.880 255.300 981.020 255.440 ;
        RECT 981.250 255.380 981.570 255.440 ;
        RECT 980.790 255.040 981.110 255.300 ;
        RECT 980.790 227.700 981.110 227.760 ;
        RECT 981.710 227.700 982.030 227.760 ;
        RECT 980.790 227.560 982.030 227.700 ;
        RECT 980.790 227.500 981.110 227.560 ;
        RECT 981.710 227.500 982.030 227.560 ;
        RECT 980.790 110.400 981.110 110.460 ;
        RECT 981.710 110.400 982.030 110.460 ;
        RECT 980.790 110.260 982.030 110.400 ;
        RECT 980.790 110.200 981.110 110.260 ;
        RECT 981.710 110.200 982.030 110.260 ;
        RECT 454.550 38.660 454.870 38.720 ;
        RECT 981.710 38.660 982.030 38.720 ;
        RECT 454.550 38.520 982.030 38.660 ;
        RECT 454.550 38.460 454.870 38.520 ;
        RECT 981.710 38.460 982.030 38.520 ;
      LAYER via ;
        RECT 980.820 1159.100 981.080 1159.360 ;
        RECT 981.280 1159.100 981.540 1159.360 ;
        RECT 980.820 1110.820 981.080 1111.080 ;
        RECT 981.740 1110.820 982.000 1111.080 ;
        RECT 981.280 1056.080 981.540 1056.340 ;
        RECT 981.740 1056.080 982.000 1056.340 ;
        RECT 979.900 1007.800 980.160 1008.060 ;
        RECT 981.280 1007.800 981.540 1008.060 ;
        RECT 981.740 944.900 982.000 945.160 ;
        RECT 981.280 896.960 981.540 897.220 ;
        RECT 981.280 814.340 981.540 814.600 ;
        RECT 981.280 813.660 981.540 813.920 ;
        RECT 981.280 710.980 981.540 711.240 ;
        RECT 980.820 710.300 981.080 710.560 ;
        RECT 980.820 614.080 981.080 614.340 ;
        RECT 981.280 614.080 981.540 614.340 ;
        RECT 980.820 565.800 981.080 566.060 ;
        RECT 981.280 565.800 981.540 566.060 ;
        RECT 981.280 379.140 981.540 379.400 ;
        RECT 981.740 379.140 982.000 379.400 ;
        RECT 981.280 255.380 981.540 255.640 ;
        RECT 980.820 255.040 981.080 255.300 ;
        RECT 980.820 227.500 981.080 227.760 ;
        RECT 981.740 227.500 982.000 227.760 ;
        RECT 980.820 110.200 981.080 110.460 ;
        RECT 981.740 110.200 982.000 110.460 ;
        RECT 454.580 38.460 454.840 38.720 ;
        RECT 981.740 38.460 982.000 38.720 ;
      LAYER met2 ;
        RECT 983.130 1221.010 983.690 1228.680 ;
        RECT 981.340 1220.870 983.690 1221.010 ;
        RECT 981.340 1159.390 981.480 1220.870 ;
        RECT 983.130 1219.680 983.690 1220.870 ;
        RECT 980.820 1159.070 981.080 1159.390 ;
        RECT 981.280 1159.070 981.540 1159.390 ;
        RECT 980.880 1111.110 981.020 1159.070 ;
        RECT 980.820 1110.790 981.080 1111.110 ;
        RECT 981.740 1110.790 982.000 1111.110 ;
        RECT 981.800 1056.370 981.940 1110.790 ;
        RECT 981.280 1056.050 981.540 1056.370 ;
        RECT 981.740 1056.050 982.000 1056.370 ;
        RECT 981.340 1008.090 981.480 1056.050 ;
        RECT 979.900 1007.770 980.160 1008.090 ;
        RECT 981.280 1007.770 981.540 1008.090 ;
        RECT 979.960 994.005 980.100 1007.770 ;
        RECT 979.890 993.635 980.170 994.005 ;
        RECT 981.730 992.275 982.010 992.645 ;
        RECT 981.800 945.190 981.940 992.275 ;
        RECT 981.740 944.870 982.000 945.190 ;
        RECT 981.280 896.930 981.540 897.250 ;
        RECT 981.340 814.630 981.480 896.930 ;
        RECT 981.280 814.310 981.540 814.630 ;
        RECT 981.280 813.630 981.540 813.950 ;
        RECT 981.340 711.270 981.480 813.630 ;
        RECT 981.280 710.950 981.540 711.270 ;
        RECT 980.820 710.270 981.080 710.590 ;
        RECT 980.880 703.645 981.020 710.270 ;
        RECT 980.810 703.275 981.090 703.645 ;
        RECT 981.270 702.595 981.550 702.965 ;
        RECT 981.340 614.370 981.480 702.595 ;
        RECT 980.820 614.050 981.080 614.370 ;
        RECT 981.280 614.050 981.540 614.370 ;
        RECT 980.880 566.090 981.020 614.050 ;
        RECT 980.820 565.770 981.080 566.090 ;
        RECT 981.280 565.770 981.540 566.090 ;
        RECT 981.340 451.930 981.480 565.770 ;
        RECT 981.340 451.790 981.940 451.930 ;
        RECT 981.800 412.490 981.940 451.790 ;
        RECT 981.340 412.350 981.940 412.490 ;
        RECT 981.340 379.430 981.480 412.350 ;
        RECT 981.280 379.110 981.540 379.430 ;
        RECT 981.740 379.110 982.000 379.430 ;
        RECT 981.800 306.410 981.940 379.110 ;
        RECT 981.340 306.270 981.940 306.410 ;
        RECT 981.340 255.670 981.480 306.270 ;
        RECT 981.280 255.350 981.540 255.670 ;
        RECT 980.820 255.010 981.080 255.330 ;
        RECT 980.880 227.790 981.020 255.010 ;
        RECT 980.820 227.470 981.080 227.790 ;
        RECT 981.740 227.470 982.000 227.790 ;
        RECT 981.800 110.570 981.940 227.470 ;
        RECT 980.880 110.490 981.940 110.570 ;
        RECT 980.820 110.430 982.000 110.490 ;
        RECT 980.820 110.170 981.080 110.430 ;
        RECT 981.740 110.170 982.000 110.430 ;
        RECT 981.800 60.250 981.940 110.170 ;
        RECT 981.800 60.110 982.400 60.250 ;
        RECT 982.260 58.890 982.400 60.110 ;
        RECT 981.800 58.750 982.400 58.890 ;
        RECT 981.800 38.750 981.940 58.750 ;
        RECT 454.580 38.430 454.840 38.750 ;
        RECT 981.740 38.430 982.000 38.750 ;
        RECT 454.640 2.400 454.780 38.430 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 979.890 993.680 980.170 993.960 ;
        RECT 981.730 992.320 982.010 992.600 ;
        RECT 980.810 703.320 981.090 703.600 ;
        RECT 981.270 702.640 981.550 702.920 ;
      LAYER met3 ;
        RECT 979.865 993.970 980.195 993.985 ;
        RECT 979.865 993.655 980.410 993.970 ;
        RECT 980.110 992.610 980.410 993.655 ;
        RECT 981.705 992.610 982.035 992.625 ;
        RECT 980.110 992.310 982.035 992.610 ;
        RECT 981.705 992.295 982.035 992.310 ;
        RECT 980.785 703.610 981.115 703.625 ;
        RECT 980.110 703.310 981.115 703.610 ;
        RECT 980.110 702.930 980.410 703.310 ;
        RECT 980.785 703.295 981.115 703.310 ;
        RECT 981.245 702.930 981.575 702.945 ;
        RECT 980.110 702.630 981.575 702.930 ;
        RECT 981.245 702.615 981.575 702.630 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 39.000 472.810 39.060 ;
        RECT 987.230 39.000 987.550 39.060 ;
        RECT 472.490 38.860 987.550 39.000 ;
        RECT 472.490 38.800 472.810 38.860 ;
        RECT 987.230 38.800 987.550 38.860 ;
      LAYER via ;
        RECT 472.520 38.800 472.780 39.060 ;
        RECT 987.260 38.800 987.520 39.060 ;
      LAYER met2 ;
        RECT 992.330 1220.330 992.890 1228.680 ;
        RECT 990.540 1220.190 992.890 1220.330 ;
        RECT 990.540 1196.530 990.680 1220.190 ;
        RECT 992.330 1219.680 992.890 1220.190 ;
        RECT 987.320 1196.390 990.680 1196.530 ;
        RECT 987.320 39.090 987.460 1196.390 ;
        RECT 472.520 38.770 472.780 39.090 ;
        RECT 987.260 38.770 987.520 39.090 ;
        RECT 472.580 2.400 472.720 38.770 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 39.340 490.750 39.400 ;
        RECT 1001.030 39.340 1001.350 39.400 ;
        RECT 490.430 39.200 1001.350 39.340 ;
        RECT 490.430 39.140 490.750 39.200 ;
        RECT 1001.030 39.140 1001.350 39.200 ;
      LAYER via ;
        RECT 490.460 39.140 490.720 39.400 ;
        RECT 1001.060 39.140 1001.320 39.400 ;
      LAYER met2 ;
        RECT 1001.530 1220.330 1002.090 1228.680 ;
        RECT 1001.120 1220.190 1002.090 1220.330 ;
        RECT 1001.120 39.430 1001.260 1220.190 ;
        RECT 1001.530 1219.680 1002.090 1220.190 ;
        RECT 490.460 39.110 490.720 39.430 ;
        RECT 1001.060 39.110 1001.320 39.430 ;
        RECT 490.520 2.400 490.660 39.110 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 39.680 508.230 39.740 ;
        RECT 1008.390 39.680 1008.710 39.740 ;
        RECT 507.910 39.540 1008.710 39.680 ;
        RECT 507.910 39.480 508.230 39.540 ;
        RECT 1008.390 39.480 1008.710 39.540 ;
      LAYER via ;
        RECT 507.940 39.480 508.200 39.740 ;
        RECT 1008.420 39.480 1008.680 39.740 ;
      LAYER met2 ;
        RECT 1010.730 1220.330 1011.290 1228.680 ;
        RECT 1008.480 1220.190 1011.290 1220.330 ;
        RECT 1008.480 39.770 1008.620 1220.190 ;
        RECT 1010.730 1219.680 1011.290 1220.190 ;
        RECT 507.940 39.450 508.200 39.770 ;
        RECT 1008.420 39.450 1008.680 39.770 ;
        RECT 508.000 2.400 508.140 39.450 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 40.020 526.170 40.080 ;
        RECT 1014.830 40.020 1015.150 40.080 ;
        RECT 525.850 39.880 1015.150 40.020 ;
        RECT 525.850 39.820 526.170 39.880 ;
        RECT 1014.830 39.820 1015.150 39.880 ;
      LAYER via ;
        RECT 525.880 39.820 526.140 40.080 ;
        RECT 1014.860 39.820 1015.120 40.080 ;
      LAYER met2 ;
        RECT 1019.930 1220.330 1020.490 1228.680 ;
        RECT 1017.680 1220.190 1020.490 1220.330 ;
        RECT 1017.680 1196.530 1017.820 1220.190 ;
        RECT 1019.930 1219.680 1020.490 1220.190 ;
        RECT 1014.920 1196.390 1017.820 1196.530 ;
        RECT 1014.920 40.110 1015.060 1196.390 ;
        RECT 525.880 39.790 526.140 40.110 ;
        RECT 1014.860 39.790 1015.120 40.110 ;
        RECT 525.940 2.400 526.080 39.790 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 40.360 544.110 40.420 ;
        RECT 1028.170 40.360 1028.490 40.420 ;
        RECT 543.790 40.220 1028.490 40.360 ;
        RECT 543.790 40.160 544.110 40.220 ;
        RECT 1028.170 40.160 1028.490 40.220 ;
      LAYER via ;
        RECT 543.820 40.160 544.080 40.420 ;
        RECT 1028.200 40.160 1028.460 40.420 ;
      LAYER met2 ;
        RECT 1029.130 1220.330 1029.690 1228.680 ;
        RECT 1028.260 1220.190 1029.690 1220.330 ;
        RECT 1028.260 40.450 1028.400 1220.190 ;
        RECT 1029.130 1219.680 1029.690 1220.190 ;
        RECT 543.820 40.130 544.080 40.450 ;
        RECT 1028.200 40.130 1028.460 40.450 ;
        RECT 543.880 2.400 544.020 40.130 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1035.145 524.365 1035.315 572.475 ;
        RECT 1035.145 331.245 1035.315 420.835 ;
        RECT 1035.605 281.605 1035.775 324.275 ;
        RECT 1035.605 186.405 1035.775 234.515 ;
        RECT 1036.065 138.465 1036.235 185.895 ;
        RECT 1035.605 89.845 1035.775 137.955 ;
      LAYER mcon ;
        RECT 1035.145 572.305 1035.315 572.475 ;
        RECT 1035.145 420.665 1035.315 420.835 ;
        RECT 1035.605 324.105 1035.775 324.275 ;
        RECT 1035.605 234.345 1035.775 234.515 ;
        RECT 1036.065 185.725 1036.235 185.895 ;
        RECT 1035.605 137.785 1035.775 137.955 ;
      LAYER met1 ;
        RECT 1035.530 1152.500 1035.850 1152.560 ;
        RECT 1035.990 1152.500 1036.310 1152.560 ;
        RECT 1035.530 1152.360 1036.310 1152.500 ;
        RECT 1035.530 1152.300 1035.850 1152.360 ;
        RECT 1035.990 1152.300 1036.310 1152.360 ;
        RECT 1035.070 966.180 1035.390 966.240 ;
        RECT 1035.990 966.180 1036.310 966.240 ;
        RECT 1035.070 966.040 1036.310 966.180 ;
        RECT 1035.070 965.980 1035.390 966.040 ;
        RECT 1035.990 965.980 1036.310 966.040 ;
        RECT 1035.070 869.620 1035.390 869.680 ;
        RECT 1035.990 869.620 1036.310 869.680 ;
        RECT 1035.070 869.480 1036.310 869.620 ;
        RECT 1035.070 869.420 1035.390 869.480 ;
        RECT 1035.990 869.420 1036.310 869.480 ;
        RECT 1035.530 787.140 1035.850 787.400 ;
        RECT 1035.620 786.720 1035.760 787.140 ;
        RECT 1035.530 786.460 1035.850 786.720 ;
        RECT 1035.530 724.440 1035.850 724.500 ;
        RECT 1035.990 724.440 1036.310 724.500 ;
        RECT 1035.530 724.300 1036.310 724.440 ;
        RECT 1035.530 724.240 1035.850 724.300 ;
        RECT 1035.990 724.240 1036.310 724.300 ;
        RECT 1035.070 572.460 1035.390 572.520 ;
        RECT 1034.875 572.320 1035.390 572.460 ;
        RECT 1035.070 572.260 1035.390 572.320 ;
        RECT 1035.085 524.520 1035.375 524.565 ;
        RECT 1035.530 524.520 1035.850 524.580 ;
        RECT 1035.085 524.380 1035.850 524.520 ;
        RECT 1035.085 524.335 1035.375 524.380 ;
        RECT 1035.530 524.320 1035.850 524.380 ;
        RECT 1035.530 476.040 1035.850 476.300 ;
        RECT 1035.620 475.560 1035.760 476.040 ;
        RECT 1035.990 475.560 1036.310 475.620 ;
        RECT 1035.620 475.420 1036.310 475.560 ;
        RECT 1035.990 475.360 1036.310 475.420 ;
        RECT 1035.070 427.960 1035.390 428.020 ;
        RECT 1035.990 427.960 1036.310 428.020 ;
        RECT 1035.070 427.820 1036.310 427.960 ;
        RECT 1035.070 427.760 1035.390 427.820 ;
        RECT 1035.990 427.760 1036.310 427.820 ;
        RECT 1035.070 420.820 1035.390 420.880 ;
        RECT 1034.875 420.680 1035.390 420.820 ;
        RECT 1035.070 420.620 1035.390 420.680 ;
        RECT 1035.085 331.400 1035.375 331.445 ;
        RECT 1035.530 331.400 1035.850 331.460 ;
        RECT 1035.085 331.260 1035.850 331.400 ;
        RECT 1035.085 331.215 1035.375 331.260 ;
        RECT 1035.530 331.200 1035.850 331.260 ;
        RECT 1035.530 324.260 1035.850 324.320 ;
        RECT 1035.335 324.120 1035.850 324.260 ;
        RECT 1035.530 324.060 1035.850 324.120 ;
        RECT 1035.530 281.760 1035.850 281.820 ;
        RECT 1035.335 281.620 1035.850 281.760 ;
        RECT 1035.530 281.560 1035.850 281.620 ;
        RECT 1035.530 234.500 1035.850 234.560 ;
        RECT 1035.335 234.360 1035.850 234.500 ;
        RECT 1035.530 234.300 1035.850 234.360 ;
        RECT 1035.545 186.375 1035.835 186.605 ;
        RECT 1035.620 185.880 1035.760 186.375 ;
        RECT 1036.005 185.880 1036.295 185.925 ;
        RECT 1035.620 185.740 1036.295 185.880 ;
        RECT 1036.005 185.695 1036.295 185.740 ;
        RECT 1035.530 138.620 1035.850 138.680 ;
        RECT 1036.005 138.620 1036.295 138.665 ;
        RECT 1035.530 138.480 1036.295 138.620 ;
        RECT 1035.530 138.420 1035.850 138.480 ;
        RECT 1036.005 138.435 1036.295 138.480 ;
        RECT 1035.530 137.940 1035.850 138.000 ;
        RECT 1035.335 137.800 1035.850 137.940 ;
        RECT 1035.530 137.740 1035.850 137.800 ;
        RECT 1035.545 90.000 1035.835 90.045 ;
        RECT 1035.990 90.000 1036.310 90.060 ;
        RECT 1035.545 89.860 1036.310 90.000 ;
        RECT 1035.545 89.815 1035.835 89.860 ;
        RECT 1035.990 89.800 1036.310 89.860 ;
        RECT 561.730 40.700 562.050 40.760 ;
        RECT 1035.990 40.700 1036.310 40.760 ;
        RECT 561.730 40.560 1036.310 40.700 ;
        RECT 561.730 40.500 562.050 40.560 ;
        RECT 1035.990 40.500 1036.310 40.560 ;
      LAYER via ;
        RECT 1035.560 1152.300 1035.820 1152.560 ;
        RECT 1036.020 1152.300 1036.280 1152.560 ;
        RECT 1035.100 965.980 1035.360 966.240 ;
        RECT 1036.020 965.980 1036.280 966.240 ;
        RECT 1035.100 869.420 1035.360 869.680 ;
        RECT 1036.020 869.420 1036.280 869.680 ;
        RECT 1035.560 787.140 1035.820 787.400 ;
        RECT 1035.560 786.460 1035.820 786.720 ;
        RECT 1035.560 724.240 1035.820 724.500 ;
        RECT 1036.020 724.240 1036.280 724.500 ;
        RECT 1035.100 572.260 1035.360 572.520 ;
        RECT 1035.560 524.320 1035.820 524.580 ;
        RECT 1035.560 476.040 1035.820 476.300 ;
        RECT 1036.020 475.360 1036.280 475.620 ;
        RECT 1035.100 427.760 1035.360 428.020 ;
        RECT 1036.020 427.760 1036.280 428.020 ;
        RECT 1035.100 420.620 1035.360 420.880 ;
        RECT 1035.560 331.200 1035.820 331.460 ;
        RECT 1035.560 324.060 1035.820 324.320 ;
        RECT 1035.560 281.560 1035.820 281.820 ;
        RECT 1035.560 234.300 1035.820 234.560 ;
        RECT 1035.560 138.420 1035.820 138.680 ;
        RECT 1035.560 137.740 1035.820 138.000 ;
        RECT 1036.020 89.800 1036.280 90.060 ;
        RECT 561.760 40.500 562.020 40.760 ;
        RECT 1036.020 40.500 1036.280 40.760 ;
      LAYER met2 ;
        RECT 1038.330 1221.010 1038.890 1228.680 ;
        RECT 1036.080 1220.870 1038.890 1221.010 ;
        RECT 1036.080 1152.590 1036.220 1220.870 ;
        RECT 1038.330 1219.680 1038.890 1220.870 ;
        RECT 1035.560 1152.270 1035.820 1152.590 ;
        RECT 1036.020 1152.270 1036.280 1152.590 ;
        RECT 1035.620 1104.165 1035.760 1152.270 ;
        RECT 1034.630 1103.795 1034.910 1104.165 ;
        RECT 1035.550 1103.795 1035.830 1104.165 ;
        RECT 1034.700 1055.885 1034.840 1103.795 ;
        RECT 1034.630 1055.515 1034.910 1055.885 ;
        RECT 1035.550 1055.515 1035.830 1055.885 ;
        RECT 1035.620 1038.770 1035.760 1055.515 ;
        RECT 1035.620 1038.630 1036.220 1038.770 ;
        RECT 1036.080 966.270 1036.220 1038.630 ;
        RECT 1035.100 965.950 1035.360 966.270 ;
        RECT 1036.020 965.950 1036.280 966.270 ;
        RECT 1035.160 947.650 1035.300 965.950 ;
        RECT 1035.160 947.510 1036.220 947.650 ;
        RECT 1036.080 869.710 1036.220 947.510 ;
        RECT 1035.100 869.390 1035.360 869.710 ;
        RECT 1036.020 869.390 1036.280 869.710 ;
        RECT 1035.160 847.010 1035.300 869.390 ;
        RECT 1035.160 846.870 1035.760 847.010 ;
        RECT 1035.620 787.430 1035.760 846.870 ;
        RECT 1035.560 787.110 1035.820 787.430 ;
        RECT 1035.560 786.430 1035.820 786.750 ;
        RECT 1035.620 724.530 1035.760 786.430 ;
        RECT 1035.560 724.210 1035.820 724.530 ;
        RECT 1036.020 724.210 1036.280 724.530 ;
        RECT 1036.080 676.445 1036.220 724.210 ;
        RECT 1035.090 676.075 1035.370 676.445 ;
        RECT 1036.010 676.075 1036.290 676.445 ;
        RECT 1035.160 651.850 1035.300 676.075 ;
        RECT 1035.160 651.710 1035.760 651.850 ;
        RECT 1035.620 580.565 1035.760 651.710 ;
        RECT 1035.550 580.195 1035.830 580.565 ;
        RECT 1035.090 579.515 1035.370 579.885 ;
        RECT 1035.160 572.550 1035.300 579.515 ;
        RECT 1035.100 572.230 1035.360 572.550 ;
        RECT 1035.560 524.290 1035.820 524.610 ;
        RECT 1035.620 476.330 1035.760 524.290 ;
        RECT 1035.560 476.010 1035.820 476.330 ;
        RECT 1036.020 475.330 1036.280 475.650 ;
        RECT 1036.080 428.050 1036.220 475.330 ;
        RECT 1035.100 427.730 1035.360 428.050 ;
        RECT 1036.020 427.730 1036.280 428.050 ;
        RECT 1035.160 420.910 1035.300 427.730 ;
        RECT 1035.100 420.590 1035.360 420.910 ;
        RECT 1035.560 331.170 1035.820 331.490 ;
        RECT 1035.620 324.350 1035.760 331.170 ;
        RECT 1035.560 324.030 1035.820 324.350 ;
        RECT 1035.560 281.530 1035.820 281.850 ;
        RECT 1035.620 234.590 1035.760 281.530 ;
        RECT 1035.560 234.270 1035.820 234.590 ;
        RECT 1035.560 138.390 1035.820 138.710 ;
        RECT 1035.620 138.030 1035.760 138.390 ;
        RECT 1035.560 137.710 1035.820 138.030 ;
        RECT 1036.020 89.770 1036.280 90.090 ;
        RECT 1036.080 40.790 1036.220 89.770 ;
        RECT 561.760 40.470 562.020 40.790 ;
        RECT 1036.020 40.470 1036.280 40.790 ;
        RECT 561.820 2.400 561.960 40.470 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 1034.630 1103.840 1034.910 1104.120 ;
        RECT 1035.550 1103.840 1035.830 1104.120 ;
        RECT 1034.630 1055.560 1034.910 1055.840 ;
        RECT 1035.550 1055.560 1035.830 1055.840 ;
        RECT 1035.090 676.120 1035.370 676.400 ;
        RECT 1036.010 676.120 1036.290 676.400 ;
        RECT 1035.550 580.240 1035.830 580.520 ;
        RECT 1035.090 579.560 1035.370 579.840 ;
      LAYER met3 ;
        RECT 1034.605 1104.130 1034.935 1104.145 ;
        RECT 1035.525 1104.130 1035.855 1104.145 ;
        RECT 1034.605 1103.830 1035.855 1104.130 ;
        RECT 1034.605 1103.815 1034.935 1103.830 ;
        RECT 1035.525 1103.815 1035.855 1103.830 ;
        RECT 1034.605 1055.850 1034.935 1055.865 ;
        RECT 1035.525 1055.850 1035.855 1055.865 ;
        RECT 1034.605 1055.550 1035.855 1055.850 ;
        RECT 1034.605 1055.535 1034.935 1055.550 ;
        RECT 1035.525 1055.535 1035.855 1055.550 ;
        RECT 1035.065 676.410 1035.395 676.425 ;
        RECT 1035.985 676.410 1036.315 676.425 ;
        RECT 1035.065 676.110 1036.315 676.410 ;
        RECT 1035.065 676.095 1035.395 676.110 ;
        RECT 1035.985 676.095 1036.315 676.110 ;
        RECT 1035.525 580.530 1035.855 580.545 ;
        RECT 1035.310 580.215 1035.855 580.530 ;
        RECT 1035.310 579.865 1035.610 580.215 ;
        RECT 1035.065 579.550 1035.610 579.865 ;
        RECT 1035.065 579.535 1035.395 579.550 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1042.045 524.365 1042.215 531.675 ;
        RECT 1042.045 475.405 1042.215 517.395 ;
        RECT 1042.505 331.585 1042.675 420.835 ;
        RECT 1042.505 276.165 1042.675 324.275 ;
        RECT 1042.965 144.925 1043.135 210.375 ;
      LAYER mcon ;
        RECT 1042.045 531.505 1042.215 531.675 ;
        RECT 1042.045 517.225 1042.215 517.395 ;
        RECT 1042.505 420.665 1042.675 420.835 ;
        RECT 1042.505 324.105 1042.675 324.275 ;
        RECT 1042.965 210.205 1043.135 210.375 ;
      LAYER met1 ;
        RECT 1042.430 1159.300 1042.750 1159.360 ;
        RECT 1045.650 1159.300 1045.970 1159.360 ;
        RECT 1042.430 1159.160 1045.970 1159.300 ;
        RECT 1042.430 1159.100 1042.750 1159.160 ;
        RECT 1045.650 1159.100 1045.970 1159.160 ;
        RECT 1042.430 1014.460 1042.750 1014.520 ;
        RECT 1042.890 1014.460 1043.210 1014.520 ;
        RECT 1042.430 1014.320 1043.210 1014.460 ;
        RECT 1042.430 1014.260 1042.750 1014.320 ;
        RECT 1042.890 1014.260 1043.210 1014.320 ;
        RECT 1041.970 1007.320 1042.290 1007.380 ;
        RECT 1042.890 1007.320 1043.210 1007.380 ;
        RECT 1041.970 1007.180 1043.210 1007.320 ;
        RECT 1041.970 1007.120 1042.290 1007.180 ;
        RECT 1042.890 1007.120 1043.210 1007.180 ;
        RECT 1042.430 869.620 1042.750 869.680 ;
        RECT 1042.890 869.620 1043.210 869.680 ;
        RECT 1042.430 869.480 1043.210 869.620 ;
        RECT 1042.430 869.420 1042.750 869.480 ;
        RECT 1042.890 869.420 1043.210 869.480 ;
        RECT 1042.430 787.140 1042.750 787.400 ;
        RECT 1042.520 786.720 1042.660 787.140 ;
        RECT 1042.430 786.460 1042.750 786.720 ;
        RECT 1042.430 724.440 1042.750 724.500 ;
        RECT 1043.350 724.440 1043.670 724.500 ;
        RECT 1042.430 724.300 1043.670 724.440 ;
        RECT 1042.430 724.240 1042.750 724.300 ;
        RECT 1043.350 724.240 1043.670 724.300 ;
        RECT 1042.430 627.880 1042.750 627.940 ;
        RECT 1043.350 627.880 1043.670 627.940 ;
        RECT 1042.430 627.740 1043.670 627.880 ;
        RECT 1042.430 627.680 1042.750 627.740 ;
        RECT 1043.350 627.680 1043.670 627.740 ;
        RECT 1042.890 602.720 1043.210 602.780 ;
        RECT 1043.350 602.720 1043.670 602.780 ;
        RECT 1042.890 602.580 1043.670 602.720 ;
        RECT 1042.890 602.520 1043.210 602.580 ;
        RECT 1043.350 602.520 1043.670 602.580 ;
        RECT 1041.985 531.660 1042.275 531.705 ;
        RECT 1042.890 531.660 1043.210 531.720 ;
        RECT 1041.985 531.520 1043.210 531.660 ;
        RECT 1041.985 531.475 1042.275 531.520 ;
        RECT 1042.890 531.460 1043.210 531.520 ;
        RECT 1041.970 524.520 1042.290 524.580 ;
        RECT 1041.775 524.380 1042.290 524.520 ;
        RECT 1041.970 524.320 1042.290 524.380 ;
        RECT 1041.970 517.380 1042.290 517.440 ;
        RECT 1041.775 517.240 1042.290 517.380 ;
        RECT 1041.970 517.180 1042.290 517.240 ;
        RECT 1041.985 475.560 1042.275 475.605 ;
        RECT 1043.810 475.560 1044.130 475.620 ;
        RECT 1041.985 475.420 1044.130 475.560 ;
        RECT 1041.985 475.375 1042.275 475.420 ;
        RECT 1043.810 475.360 1044.130 475.420 ;
        RECT 1042.445 420.820 1042.735 420.865 ;
        RECT 1042.890 420.820 1043.210 420.880 ;
        RECT 1042.445 420.680 1043.210 420.820 ;
        RECT 1042.445 420.635 1042.735 420.680 ;
        RECT 1042.890 420.620 1043.210 420.680 ;
        RECT 1042.430 331.740 1042.750 331.800 ;
        RECT 1042.235 331.600 1042.750 331.740 ;
        RECT 1042.430 331.540 1042.750 331.600 ;
        RECT 1042.430 324.260 1042.750 324.320 ;
        RECT 1042.235 324.120 1042.750 324.260 ;
        RECT 1042.430 324.060 1042.750 324.120 ;
        RECT 1042.430 276.320 1042.750 276.380 ;
        RECT 1042.235 276.180 1042.750 276.320 ;
        RECT 1042.430 276.120 1042.750 276.180 ;
        RECT 1042.890 210.360 1043.210 210.420 ;
        RECT 1042.695 210.220 1043.210 210.360 ;
        RECT 1042.890 210.160 1043.210 210.220 ;
        RECT 1042.890 145.080 1043.210 145.140 ;
        RECT 1042.695 144.940 1043.210 145.080 ;
        RECT 1042.890 144.880 1043.210 144.940 ;
        RECT 579.670 41.040 579.990 41.100 ;
        RECT 1042.890 41.040 1043.210 41.100 ;
        RECT 579.670 40.900 1043.210 41.040 ;
        RECT 579.670 40.840 579.990 40.900 ;
        RECT 1042.890 40.840 1043.210 40.900 ;
      LAYER via ;
        RECT 1042.460 1159.100 1042.720 1159.360 ;
        RECT 1045.680 1159.100 1045.940 1159.360 ;
        RECT 1042.460 1014.260 1042.720 1014.520 ;
        RECT 1042.920 1014.260 1043.180 1014.520 ;
        RECT 1042.000 1007.120 1042.260 1007.380 ;
        RECT 1042.920 1007.120 1043.180 1007.380 ;
        RECT 1042.460 869.420 1042.720 869.680 ;
        RECT 1042.920 869.420 1043.180 869.680 ;
        RECT 1042.460 787.140 1042.720 787.400 ;
        RECT 1042.460 786.460 1042.720 786.720 ;
        RECT 1042.460 724.240 1042.720 724.500 ;
        RECT 1043.380 724.240 1043.640 724.500 ;
        RECT 1042.460 627.680 1042.720 627.940 ;
        RECT 1043.380 627.680 1043.640 627.940 ;
        RECT 1042.920 602.520 1043.180 602.780 ;
        RECT 1043.380 602.520 1043.640 602.780 ;
        RECT 1042.920 531.460 1043.180 531.720 ;
        RECT 1042.000 524.320 1042.260 524.580 ;
        RECT 1042.000 517.180 1042.260 517.440 ;
        RECT 1043.840 475.360 1044.100 475.620 ;
        RECT 1042.920 420.620 1043.180 420.880 ;
        RECT 1042.460 331.540 1042.720 331.800 ;
        RECT 1042.460 324.060 1042.720 324.320 ;
        RECT 1042.460 276.120 1042.720 276.380 ;
        RECT 1042.920 210.160 1043.180 210.420 ;
        RECT 1042.920 144.880 1043.180 145.140 ;
        RECT 579.700 40.840 579.960 41.100 ;
        RECT 1042.920 40.840 1043.180 41.100 ;
      LAYER met2 ;
        RECT 1047.530 1220.330 1048.090 1228.680 ;
        RECT 1045.740 1220.190 1048.090 1220.330 ;
        RECT 1045.740 1159.390 1045.880 1220.190 ;
        RECT 1047.530 1219.680 1048.090 1220.190 ;
        RECT 1042.460 1159.070 1042.720 1159.390 ;
        RECT 1045.680 1159.070 1045.940 1159.390 ;
        RECT 1042.520 1014.550 1042.660 1159.070 ;
        RECT 1042.460 1014.230 1042.720 1014.550 ;
        RECT 1042.920 1014.230 1043.180 1014.550 ;
        RECT 1042.980 1007.410 1043.120 1014.230 ;
        RECT 1042.000 1007.090 1042.260 1007.410 ;
        RECT 1042.920 1007.090 1043.180 1007.410 ;
        RECT 1042.060 959.325 1042.200 1007.090 ;
        RECT 1041.990 958.955 1042.270 959.325 ;
        RECT 1042.910 958.955 1043.190 959.325 ;
        RECT 1042.980 942.210 1043.120 958.955 ;
        RECT 1042.520 942.070 1043.120 942.210 ;
        RECT 1042.520 869.710 1042.660 942.070 ;
        RECT 1042.460 869.390 1042.720 869.710 ;
        RECT 1042.920 869.390 1043.180 869.710 ;
        RECT 1042.980 821.170 1043.120 869.390 ;
        RECT 1042.520 821.030 1043.120 821.170 ;
        RECT 1042.520 787.430 1042.660 821.030 ;
        RECT 1042.460 787.110 1042.720 787.430 ;
        RECT 1042.460 786.430 1042.720 786.750 ;
        RECT 1042.520 724.530 1042.660 786.430 ;
        RECT 1042.460 724.210 1042.720 724.530 ;
        RECT 1043.380 724.210 1043.640 724.530 ;
        RECT 1043.440 699.450 1043.580 724.210 ;
        RECT 1042.980 699.310 1043.580 699.450 ;
        RECT 1042.980 628.050 1043.120 699.310 ;
        RECT 1042.520 627.970 1043.120 628.050 ;
        RECT 1042.460 627.910 1043.120 627.970 ;
        RECT 1042.460 627.650 1042.720 627.910 ;
        RECT 1043.380 627.650 1043.640 627.970 ;
        RECT 1043.440 602.810 1043.580 627.650 ;
        RECT 1042.920 602.490 1043.180 602.810 ;
        RECT 1043.380 602.490 1043.640 602.810 ;
        RECT 1042.980 531.750 1043.120 602.490 ;
        RECT 1042.920 531.430 1043.180 531.750 ;
        RECT 1042.000 524.290 1042.260 524.610 ;
        RECT 1042.060 517.470 1042.200 524.290 ;
        RECT 1042.000 517.150 1042.260 517.470 ;
        RECT 1043.840 475.330 1044.100 475.650 ;
        RECT 1043.900 428.245 1044.040 475.330 ;
        RECT 1042.910 427.875 1043.190 428.245 ;
        RECT 1043.830 427.875 1044.110 428.245 ;
        RECT 1042.980 420.910 1043.120 427.875 ;
        RECT 1042.920 420.590 1043.180 420.910 ;
        RECT 1042.460 331.510 1042.720 331.830 ;
        RECT 1042.520 324.350 1042.660 331.510 ;
        RECT 1042.460 324.030 1042.720 324.350 ;
        RECT 1042.460 276.090 1042.720 276.410 ;
        RECT 1042.520 258.810 1042.660 276.090 ;
        RECT 1042.520 258.670 1043.120 258.810 ;
        RECT 1042.980 210.450 1043.120 258.670 ;
        RECT 1042.920 210.130 1043.180 210.450 ;
        RECT 1042.920 144.850 1043.180 145.170 ;
        RECT 1042.980 110.570 1043.120 144.850 ;
        RECT 1042.520 110.430 1043.120 110.570 ;
        RECT 1042.520 109.890 1042.660 110.430 ;
        RECT 1042.520 109.750 1043.120 109.890 ;
        RECT 1042.980 41.130 1043.120 109.750 ;
        RECT 579.700 40.810 579.960 41.130 ;
        RECT 1042.920 40.810 1043.180 41.130 ;
        RECT 579.760 2.400 579.900 40.810 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 1041.990 959.000 1042.270 959.280 ;
        RECT 1042.910 959.000 1043.190 959.280 ;
        RECT 1042.910 427.920 1043.190 428.200 ;
        RECT 1043.830 427.920 1044.110 428.200 ;
      LAYER met3 ;
        RECT 1041.965 959.290 1042.295 959.305 ;
        RECT 1042.885 959.290 1043.215 959.305 ;
        RECT 1041.965 958.990 1043.215 959.290 ;
        RECT 1041.965 958.975 1042.295 958.990 ;
        RECT 1042.885 958.975 1043.215 958.990 ;
        RECT 1042.885 428.210 1043.215 428.225 ;
        RECT 1043.805 428.210 1044.135 428.225 ;
        RECT 1042.885 427.910 1044.135 428.210 ;
        RECT 1042.885 427.895 1043.215 427.910 ;
        RECT 1043.805 427.895 1044.135 427.910 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.550 25.400 86.870 25.460 ;
        RECT 794.030 25.400 794.350 25.460 ;
        RECT 86.550 25.260 794.350 25.400 ;
        RECT 86.550 25.200 86.870 25.260 ;
        RECT 794.030 25.200 794.350 25.260 ;
      LAYER via ;
        RECT 86.580 25.200 86.840 25.460 ;
        RECT 794.060 25.200 794.320 25.460 ;
      LAYER met2 ;
        RECT 793.610 1220.330 794.170 1228.680 ;
        RECT 793.610 1219.680 794.260 1220.330 ;
        RECT 794.120 25.490 794.260 1219.680 ;
        RECT 86.580 25.170 86.840 25.490 ;
        RECT 794.060 25.170 794.320 25.490 ;
        RECT 86.640 12.650 86.780 25.170 ;
        RECT 86.180 12.510 86.780 12.650 ;
        RECT 86.180 2.400 86.320 12.510 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 41.380 597.470 41.440 ;
        RECT 1055.770 41.380 1056.090 41.440 ;
        RECT 597.150 41.240 1056.090 41.380 ;
        RECT 597.150 41.180 597.470 41.240 ;
        RECT 1055.770 41.180 1056.090 41.240 ;
      LAYER via ;
        RECT 597.180 41.180 597.440 41.440 ;
        RECT 1055.800 41.180 1056.060 41.440 ;
      LAYER met2 ;
        RECT 1056.730 1220.330 1057.290 1228.680 ;
        RECT 1055.860 1220.190 1057.290 1220.330 ;
        RECT 1055.860 41.470 1056.000 1220.190 ;
        RECT 1056.730 1219.680 1057.290 1220.190 ;
        RECT 597.180 41.150 597.440 41.470 ;
        RECT 1055.800 41.150 1056.060 41.470 ;
        RECT 597.240 2.400 597.380 41.150 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 37.640 615.410 37.700 ;
        RECT 1063.590 37.640 1063.910 37.700 ;
        RECT 615.090 37.500 1063.910 37.640 ;
        RECT 615.090 37.440 615.410 37.500 ;
        RECT 1063.590 37.440 1063.910 37.500 ;
      LAYER via ;
        RECT 615.120 37.440 615.380 37.700 ;
        RECT 1063.620 37.440 1063.880 37.700 ;
      LAYER met2 ;
        RECT 1065.930 1220.330 1066.490 1228.680 ;
        RECT 1063.680 1220.190 1066.490 1220.330 ;
        RECT 1063.680 37.730 1063.820 1220.190 ;
        RECT 1065.930 1219.680 1066.490 1220.190 ;
        RECT 615.120 37.410 615.380 37.730 ;
        RECT 1063.620 37.410 1063.880 37.730 ;
        RECT 615.180 2.400 615.320 37.410 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 744.885 24.905 745.055 25.755 ;
      LAYER mcon ;
        RECT 744.885 25.585 745.055 25.755 ;
      LAYER met1 ;
        RECT 109.550 25.740 109.870 25.800 ;
        RECT 744.825 25.740 745.115 25.785 ;
        RECT 109.550 25.600 745.115 25.740 ;
        RECT 109.550 25.540 109.870 25.600 ;
        RECT 744.825 25.555 745.115 25.600 ;
        RECT 800.930 25.400 801.250 25.460 ;
        RECT 794.580 25.260 801.250 25.400 ;
        RECT 744.825 25.060 745.115 25.105 ;
        RECT 794.580 25.060 794.720 25.260 ;
        RECT 800.930 25.200 801.250 25.260 ;
        RECT 744.825 24.920 794.720 25.060 ;
        RECT 744.825 24.875 745.115 24.920 ;
      LAYER via ;
        RECT 109.580 25.540 109.840 25.800 ;
        RECT 800.960 25.200 801.220 25.460 ;
      LAYER met2 ;
        RECT 806.030 1220.330 806.590 1228.680 ;
        RECT 803.780 1220.190 806.590 1220.330 ;
        RECT 803.780 1195.850 803.920 1220.190 ;
        RECT 806.030 1219.680 806.590 1220.190 ;
        RECT 801.020 1195.710 803.920 1195.850 ;
        RECT 109.580 25.510 109.840 25.830 ;
        RECT 109.640 2.400 109.780 25.510 ;
        RECT 801.020 25.490 801.160 1195.710 ;
        RECT 800.960 25.170 801.220 25.490 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 814.805 689.605 814.975 717.655 ;
        RECT 814.805 572.645 814.975 620.755 ;
        RECT 814.805 379.525 814.975 427.635 ;
        RECT 814.345 282.965 814.515 331.075 ;
        RECT 276.145 22.865 276.315 26.095 ;
        RECT 323.985 22.865 324.155 26.095 ;
        RECT 372.745 20.825 372.915 26.095 ;
        RECT 418.745 25.925 420.755 26.095 ;
        RECT 469.345 25.925 469.515 27.795 ;
        RECT 517.185 25.925 517.355 27.795 ;
        RECT 565.945 25.925 566.115 28.475 ;
        RECT 613.785 25.925 613.955 28.475 ;
        RECT 662.545 25.925 662.715 28.475 ;
        RECT 710.385 25.925 710.555 28.475 ;
        RECT 418.745 20.825 418.915 25.925 ;
      LAYER mcon ;
        RECT 814.805 717.485 814.975 717.655 ;
        RECT 814.805 620.585 814.975 620.755 ;
        RECT 814.805 427.465 814.975 427.635 ;
        RECT 814.345 330.905 814.515 331.075 ;
        RECT 565.945 28.305 566.115 28.475 ;
        RECT 469.345 27.625 469.515 27.795 ;
        RECT 276.145 25.925 276.315 26.095 ;
        RECT 323.985 25.925 324.155 26.095 ;
        RECT 372.745 25.925 372.915 26.095 ;
        RECT 420.585 25.925 420.755 26.095 ;
        RECT 517.185 27.625 517.355 27.795 ;
        RECT 613.785 28.305 613.955 28.475 ;
        RECT 662.545 28.305 662.715 28.475 ;
        RECT 710.385 28.305 710.555 28.475 ;
      LAYER met1 ;
        RECT 815.190 1159.300 815.510 1159.360 ;
        RECT 816.110 1159.300 816.430 1159.360 ;
        RECT 815.190 1159.160 816.430 1159.300 ;
        RECT 815.190 1159.100 815.510 1159.160 ;
        RECT 816.110 1159.100 816.430 1159.160 ;
        RECT 814.270 1028.400 814.590 1028.460 ;
        RECT 815.190 1028.400 815.510 1028.460 ;
        RECT 814.270 1028.260 815.510 1028.400 ;
        RECT 814.270 1028.200 814.590 1028.260 ;
        RECT 815.190 1028.200 815.510 1028.260 ;
        RECT 814.270 931.840 814.590 931.900 ;
        RECT 815.190 931.840 815.510 931.900 ;
        RECT 814.270 931.700 815.510 931.840 ;
        RECT 814.270 931.640 814.590 931.700 ;
        RECT 815.190 931.640 815.510 931.700 ;
        RECT 814.730 883.360 815.050 883.620 ;
        RECT 814.820 882.880 814.960 883.360 ;
        RECT 815.190 882.880 815.510 882.940 ;
        RECT 814.820 882.740 815.510 882.880 ;
        RECT 815.190 882.680 815.510 882.740 ;
        RECT 814.270 835.280 814.590 835.340 ;
        RECT 815.190 835.280 815.510 835.340 ;
        RECT 814.270 835.140 815.510 835.280 ;
        RECT 814.270 835.080 814.590 835.140 ;
        RECT 815.190 835.080 815.510 835.140 ;
        RECT 814.730 786.800 815.050 787.060 ;
        RECT 814.820 786.320 814.960 786.800 ;
        RECT 815.190 786.320 815.510 786.380 ;
        RECT 814.820 786.180 815.510 786.320 ;
        RECT 815.190 786.120 815.510 786.180 ;
        RECT 814.270 738.380 814.590 738.440 ;
        RECT 815.190 738.380 815.510 738.440 ;
        RECT 814.270 738.240 815.510 738.380 ;
        RECT 814.270 738.180 814.590 738.240 ;
        RECT 815.190 738.180 815.510 738.240 ;
        RECT 814.730 717.640 815.050 717.700 ;
        RECT 814.535 717.500 815.050 717.640 ;
        RECT 814.730 717.440 815.050 717.500 ;
        RECT 814.730 689.760 815.050 689.820 ;
        RECT 814.535 689.620 815.050 689.760 ;
        RECT 814.730 689.560 815.050 689.620 ;
        RECT 814.270 641.820 814.590 641.880 ;
        RECT 815.190 641.820 815.510 641.880 ;
        RECT 814.270 641.680 815.510 641.820 ;
        RECT 814.270 641.620 814.590 641.680 ;
        RECT 815.190 641.620 815.510 641.680 ;
        RECT 814.730 620.740 815.050 620.800 ;
        RECT 814.535 620.600 815.050 620.740 ;
        RECT 814.730 620.540 815.050 620.600 ;
        RECT 814.745 572.800 815.035 572.845 ;
        RECT 815.190 572.800 815.510 572.860 ;
        RECT 814.745 572.660 815.510 572.800 ;
        RECT 814.745 572.615 815.035 572.660 ;
        RECT 815.190 572.600 815.510 572.660 ;
        RECT 814.270 545.260 814.590 545.320 ;
        RECT 815.190 545.260 815.510 545.320 ;
        RECT 814.270 545.120 815.510 545.260 ;
        RECT 814.270 545.060 814.590 545.120 ;
        RECT 815.190 545.060 815.510 545.120 ;
        RECT 814.730 496.780 815.050 497.040 ;
        RECT 814.820 496.640 814.960 496.780 ;
        RECT 815.190 496.640 815.510 496.700 ;
        RECT 814.820 496.500 815.510 496.640 ;
        RECT 815.190 496.440 815.510 496.500 ;
        RECT 814.270 483.040 814.590 483.100 ;
        RECT 815.190 483.040 815.510 483.100 ;
        RECT 814.270 482.900 815.510 483.040 ;
        RECT 814.270 482.840 814.590 482.900 ;
        RECT 815.190 482.840 815.510 482.900 ;
        RECT 814.730 427.620 815.050 427.680 ;
        RECT 814.535 427.480 815.050 427.620 ;
        RECT 814.730 427.420 815.050 427.480 ;
        RECT 814.745 379.680 815.035 379.725 ;
        RECT 816.110 379.680 816.430 379.740 ;
        RECT 814.745 379.540 816.430 379.680 ;
        RECT 814.745 379.495 815.035 379.540 ;
        RECT 816.110 379.480 816.430 379.540 ;
        RECT 814.730 338.540 815.050 338.600 ;
        RECT 816.110 338.540 816.430 338.600 ;
        RECT 814.730 338.400 816.430 338.540 ;
        RECT 814.730 338.340 815.050 338.400 ;
        RECT 816.110 338.340 816.430 338.400 ;
        RECT 814.285 331.060 814.575 331.105 ;
        RECT 814.730 331.060 815.050 331.120 ;
        RECT 814.285 330.920 815.050 331.060 ;
        RECT 814.285 330.875 814.575 330.920 ;
        RECT 814.730 330.860 815.050 330.920 ;
        RECT 814.270 283.120 814.590 283.180 ;
        RECT 814.270 282.980 814.785 283.120 ;
        RECT 814.270 282.920 814.590 282.980 ;
        RECT 565.885 28.460 566.175 28.505 ;
        RECT 613.725 28.460 614.015 28.505 ;
        RECT 565.885 28.320 614.015 28.460 ;
        RECT 565.885 28.275 566.175 28.320 ;
        RECT 613.725 28.275 614.015 28.320 ;
        RECT 662.485 28.460 662.775 28.505 ;
        RECT 710.325 28.460 710.615 28.505 ;
        RECT 662.485 28.320 710.615 28.460 ;
        RECT 662.485 28.275 662.775 28.320 ;
        RECT 710.325 28.275 710.615 28.320 ;
        RECT 469.285 27.780 469.575 27.825 ;
        RECT 517.125 27.780 517.415 27.825 ;
        RECT 469.285 27.640 517.415 27.780 ;
        RECT 469.285 27.595 469.575 27.640 ;
        RECT 517.125 27.595 517.415 27.640 ;
        RECT 133.470 26.080 133.790 26.140 ;
        RECT 276.085 26.080 276.375 26.125 ;
        RECT 133.470 25.940 276.375 26.080 ;
        RECT 133.470 25.880 133.790 25.940 ;
        RECT 276.085 25.895 276.375 25.940 ;
        RECT 323.925 26.080 324.215 26.125 ;
        RECT 372.685 26.080 372.975 26.125 ;
        RECT 323.925 25.940 372.975 26.080 ;
        RECT 323.925 25.895 324.215 25.940 ;
        RECT 372.685 25.895 372.975 25.940 ;
        RECT 420.525 26.080 420.815 26.125 ;
        RECT 469.285 26.080 469.575 26.125 ;
        RECT 420.525 25.940 469.575 26.080 ;
        RECT 420.525 25.895 420.815 25.940 ;
        RECT 469.285 25.895 469.575 25.940 ;
        RECT 517.125 26.080 517.415 26.125 ;
        RECT 565.885 26.080 566.175 26.125 ;
        RECT 517.125 25.940 566.175 26.080 ;
        RECT 517.125 25.895 517.415 25.940 ;
        RECT 565.885 25.895 566.175 25.940 ;
        RECT 613.725 26.080 614.015 26.125 ;
        RECT 662.485 26.080 662.775 26.125 ;
        RECT 613.725 25.940 662.775 26.080 ;
        RECT 613.725 25.895 614.015 25.940 ;
        RECT 662.485 25.895 662.775 25.940 ;
        RECT 710.325 26.080 710.615 26.125 ;
        RECT 710.325 25.940 745.500 26.080 ;
        RECT 710.325 25.895 710.615 25.940 ;
        RECT 745.360 25.740 745.500 25.940 ;
        RECT 814.270 25.740 814.590 25.800 ;
        RECT 745.360 25.600 814.590 25.740 ;
        RECT 814.270 25.540 814.590 25.600 ;
        RECT 276.085 23.020 276.375 23.065 ;
        RECT 323.925 23.020 324.215 23.065 ;
        RECT 276.085 22.880 324.215 23.020 ;
        RECT 276.085 22.835 276.375 22.880 ;
        RECT 323.925 22.835 324.215 22.880 ;
        RECT 372.685 20.980 372.975 21.025 ;
        RECT 418.685 20.980 418.975 21.025 ;
        RECT 372.685 20.840 418.975 20.980 ;
        RECT 372.685 20.795 372.975 20.840 ;
        RECT 418.685 20.795 418.975 20.840 ;
      LAYER via ;
        RECT 815.220 1159.100 815.480 1159.360 ;
        RECT 816.140 1159.100 816.400 1159.360 ;
        RECT 814.300 1028.200 814.560 1028.460 ;
        RECT 815.220 1028.200 815.480 1028.460 ;
        RECT 814.300 931.640 814.560 931.900 ;
        RECT 815.220 931.640 815.480 931.900 ;
        RECT 814.760 883.360 815.020 883.620 ;
        RECT 815.220 882.680 815.480 882.940 ;
        RECT 814.300 835.080 814.560 835.340 ;
        RECT 815.220 835.080 815.480 835.340 ;
        RECT 814.760 786.800 815.020 787.060 ;
        RECT 815.220 786.120 815.480 786.380 ;
        RECT 814.300 738.180 814.560 738.440 ;
        RECT 815.220 738.180 815.480 738.440 ;
        RECT 814.760 717.440 815.020 717.700 ;
        RECT 814.760 689.560 815.020 689.820 ;
        RECT 814.300 641.620 814.560 641.880 ;
        RECT 815.220 641.620 815.480 641.880 ;
        RECT 814.760 620.540 815.020 620.800 ;
        RECT 815.220 572.600 815.480 572.860 ;
        RECT 814.300 545.060 814.560 545.320 ;
        RECT 815.220 545.060 815.480 545.320 ;
        RECT 814.760 496.780 815.020 497.040 ;
        RECT 815.220 496.440 815.480 496.700 ;
        RECT 814.300 482.840 814.560 483.100 ;
        RECT 815.220 482.840 815.480 483.100 ;
        RECT 814.760 427.420 815.020 427.680 ;
        RECT 816.140 379.480 816.400 379.740 ;
        RECT 814.760 338.340 815.020 338.600 ;
        RECT 816.140 338.340 816.400 338.600 ;
        RECT 814.760 330.860 815.020 331.120 ;
        RECT 814.300 282.920 814.560 283.180 ;
        RECT 133.500 25.880 133.760 26.140 ;
        RECT 814.300 25.540 814.560 25.800 ;
      LAYER met2 ;
        RECT 818.450 1221.010 819.010 1228.680 ;
        RECT 816.200 1220.870 819.010 1221.010 ;
        RECT 816.200 1159.390 816.340 1220.870 ;
        RECT 818.450 1219.680 819.010 1220.870 ;
        RECT 815.220 1159.070 815.480 1159.390 ;
        RECT 816.140 1159.070 816.400 1159.390 ;
        RECT 815.280 1028.490 815.420 1159.070 ;
        RECT 814.300 1028.170 814.560 1028.490 ;
        RECT 815.220 1028.170 815.480 1028.490 ;
        RECT 814.360 1027.890 814.500 1028.170 ;
        RECT 814.360 1027.750 814.960 1027.890 ;
        RECT 814.820 980.290 814.960 1027.750 ;
        RECT 814.820 980.150 815.420 980.290 ;
        RECT 815.280 931.930 815.420 980.150 ;
        RECT 814.300 931.610 814.560 931.930 ;
        RECT 815.220 931.610 815.480 931.930 ;
        RECT 814.360 931.330 814.500 931.610 ;
        RECT 814.360 931.190 814.960 931.330 ;
        RECT 814.820 883.650 814.960 931.190 ;
        RECT 814.760 883.330 815.020 883.650 ;
        RECT 815.220 882.650 815.480 882.970 ;
        RECT 815.280 835.370 815.420 882.650 ;
        RECT 814.300 835.050 814.560 835.370 ;
        RECT 815.220 835.050 815.480 835.370 ;
        RECT 814.360 834.770 814.500 835.050 ;
        RECT 814.360 834.630 814.960 834.770 ;
        RECT 814.820 787.090 814.960 834.630 ;
        RECT 814.760 786.770 815.020 787.090 ;
        RECT 815.220 786.090 815.480 786.410 ;
        RECT 815.280 738.470 815.420 786.090 ;
        RECT 814.300 738.210 814.560 738.470 ;
        RECT 814.300 738.150 814.960 738.210 ;
        RECT 815.220 738.150 815.480 738.470 ;
        RECT 814.360 738.070 814.960 738.150 ;
        RECT 814.820 717.730 814.960 738.070 ;
        RECT 814.760 717.410 815.020 717.730 ;
        RECT 814.760 689.530 815.020 689.850 ;
        RECT 814.820 669.530 814.960 689.530 ;
        RECT 814.820 669.390 815.420 669.530 ;
        RECT 815.280 641.910 815.420 669.390 ;
        RECT 814.300 641.650 814.560 641.910 ;
        RECT 814.300 641.590 814.960 641.650 ;
        RECT 815.220 641.590 815.480 641.910 ;
        RECT 814.360 641.510 814.960 641.590 ;
        RECT 814.820 620.830 814.960 641.510 ;
        RECT 814.760 620.510 815.020 620.830 ;
        RECT 815.220 572.570 815.480 572.890 ;
        RECT 815.280 545.350 815.420 572.570 ;
        RECT 814.300 545.090 814.560 545.350 ;
        RECT 814.300 545.030 814.960 545.090 ;
        RECT 815.220 545.030 815.480 545.350 ;
        RECT 814.360 544.950 814.960 545.030 ;
        RECT 814.820 497.070 814.960 544.950 ;
        RECT 814.760 496.750 815.020 497.070 ;
        RECT 815.220 496.410 815.480 496.730 ;
        RECT 815.280 483.130 815.420 496.410 ;
        RECT 814.300 482.810 814.560 483.130 ;
        RECT 815.220 482.810 815.480 483.130 ;
        RECT 814.360 435.725 814.500 482.810 ;
        RECT 814.290 435.355 814.570 435.725 ;
        RECT 814.750 434.675 815.030 435.045 ;
        RECT 814.820 427.710 814.960 434.675 ;
        RECT 814.760 427.390 815.020 427.710 ;
        RECT 816.140 379.450 816.400 379.770 ;
        RECT 816.200 338.630 816.340 379.450 ;
        RECT 814.760 338.310 815.020 338.630 ;
        RECT 816.140 338.310 816.400 338.630 ;
        RECT 814.820 331.150 814.960 338.310 ;
        RECT 814.760 330.830 815.020 331.150 ;
        RECT 814.300 282.890 814.560 283.210 ;
        RECT 814.360 241.810 814.500 282.890 ;
        RECT 814.360 241.670 814.960 241.810 ;
        RECT 814.820 210.530 814.960 241.670 ;
        RECT 814.820 210.390 816.340 210.530 ;
        RECT 816.200 192.850 816.340 210.390 ;
        RECT 815.740 192.710 816.340 192.850 ;
        RECT 815.740 168.370 815.880 192.710 ;
        RECT 815.280 168.230 815.880 168.370 ;
        RECT 815.280 62.290 815.420 168.230 ;
        RECT 814.360 62.150 815.420 62.290 ;
        RECT 133.500 25.850 133.760 26.170 ;
        RECT 133.560 2.400 133.700 25.850 ;
        RECT 814.360 25.830 814.500 62.150 ;
        RECT 814.300 25.510 814.560 25.830 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 814.290 435.400 814.570 435.680 ;
        RECT 814.750 434.720 815.030 435.000 ;
      LAYER met3 ;
        RECT 814.265 435.690 814.595 435.705 ;
        RECT 814.265 435.375 814.810 435.690 ;
        RECT 814.510 435.025 814.810 435.375 ;
        RECT 814.510 434.710 815.055 435.025 ;
        RECT 814.725 434.695 815.055 434.710 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 760.525 26.605 761.615 26.775 ;
        RECT 760.525 26.265 760.695 26.605 ;
        RECT 804.225 25.245 804.395 26.435 ;
      LAYER mcon ;
        RECT 761.445 26.605 761.615 26.775 ;
        RECT 804.225 26.265 804.395 26.435 ;
      LAYER met1 ;
        RECT 821.630 1196.700 821.950 1196.760 ;
        RECT 826.230 1196.700 826.550 1196.760 ;
        RECT 821.630 1196.560 826.550 1196.700 ;
        RECT 821.630 1196.500 821.950 1196.560 ;
        RECT 826.230 1196.500 826.550 1196.560 ;
        RECT 761.385 26.760 761.675 26.805 ;
        RECT 761.385 26.620 762.980 26.760 ;
        RECT 761.385 26.575 761.675 26.620 ;
        RECT 151.410 26.420 151.730 26.480 ;
        RECT 760.465 26.420 760.755 26.465 ;
        RECT 151.410 26.280 760.755 26.420 ;
        RECT 762.840 26.420 762.980 26.620 ;
        RECT 804.165 26.420 804.455 26.465 ;
        RECT 762.840 26.280 804.455 26.420 ;
        RECT 151.410 26.220 151.730 26.280 ;
        RECT 760.465 26.235 760.755 26.280 ;
        RECT 804.165 26.235 804.455 26.280 ;
        RECT 821.630 25.740 821.950 25.800 ;
        RECT 814.820 25.600 821.950 25.740 ;
        RECT 804.165 25.400 804.455 25.445 ;
        RECT 814.820 25.400 814.960 25.600 ;
        RECT 821.630 25.540 821.950 25.600 ;
        RECT 804.165 25.260 814.960 25.400 ;
        RECT 804.165 25.215 804.455 25.260 ;
      LAYER via ;
        RECT 821.660 1196.500 821.920 1196.760 ;
        RECT 826.260 1196.500 826.520 1196.760 ;
        RECT 151.440 26.220 151.700 26.480 ;
        RECT 821.660 25.540 821.920 25.800 ;
      LAYER met2 ;
        RECT 827.650 1220.330 828.210 1228.680 ;
        RECT 826.320 1220.190 828.210 1220.330 ;
        RECT 826.320 1196.790 826.460 1220.190 ;
        RECT 827.650 1219.680 828.210 1220.190 ;
        RECT 821.660 1196.470 821.920 1196.790 ;
        RECT 826.260 1196.470 826.520 1196.790 ;
        RECT 151.440 26.190 151.700 26.510 ;
        RECT 151.500 2.400 151.640 26.190 ;
        RECT 821.720 25.830 821.860 1196.470 ;
        RECT 821.660 25.510 821.920 25.830 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 276.145 26.605 276.775 26.775 ;
        RECT 276.605 22.185 276.775 26.605 ;
        RECT 323.525 26.605 324.155 26.775 ;
        RECT 372.745 26.605 373.375 26.775 ;
        RECT 323.525 22.185 323.695 26.605 ;
        RECT 373.205 21.165 373.375 26.605 ;
        RECT 400.805 21.165 400.975 27.795 ;
        RECT 420.585 26.605 420.755 27.795 ;
        RECT 811.125 25.925 811.295 26.775 ;
      LAYER mcon ;
        RECT 400.805 27.625 400.975 27.795 ;
        RECT 323.985 26.605 324.155 26.775 ;
        RECT 420.585 27.625 420.755 27.795 ;
        RECT 811.125 26.605 811.295 26.775 ;
      LAYER met1 ;
        RECT 400.745 27.780 401.035 27.825 ;
        RECT 420.525 27.780 420.815 27.825 ;
        RECT 400.745 27.640 420.815 27.780 ;
        RECT 400.745 27.595 401.035 27.640 ;
        RECT 420.525 27.595 420.815 27.640 ;
        RECT 169.350 26.760 169.670 26.820 ;
        RECT 276.085 26.760 276.375 26.805 ;
        RECT 169.350 26.620 276.375 26.760 ;
        RECT 169.350 26.560 169.670 26.620 ;
        RECT 276.085 26.575 276.375 26.620 ;
        RECT 323.925 26.760 324.215 26.805 ;
        RECT 372.685 26.760 372.975 26.805 ;
        RECT 323.925 26.620 372.975 26.760 ;
        RECT 323.925 26.575 324.215 26.620 ;
        RECT 372.685 26.575 372.975 26.620 ;
        RECT 420.525 26.760 420.815 26.805 ;
        RECT 469.270 26.760 469.590 26.820 ;
        RECT 420.525 26.620 469.590 26.760 ;
        RECT 420.525 26.575 420.815 26.620 ;
        RECT 469.270 26.560 469.590 26.620 ;
        RECT 517.110 26.760 517.430 26.820 ;
        RECT 565.870 26.760 566.190 26.820 ;
        RECT 517.110 26.620 566.190 26.760 ;
        RECT 517.110 26.560 517.430 26.620 ;
        RECT 565.870 26.560 566.190 26.620 ;
        RECT 613.250 26.760 613.570 26.820 ;
        RECT 662.470 26.760 662.790 26.820 ;
        RECT 613.250 26.620 662.790 26.760 ;
        RECT 613.250 26.560 613.570 26.620 ;
        RECT 662.470 26.560 662.790 26.620 ;
        RECT 709.850 26.760 710.170 26.820 ;
        RECT 811.065 26.760 811.355 26.805 ;
        RECT 835.430 26.760 835.750 26.820 ;
        RECT 709.850 26.620 761.140 26.760 ;
        RECT 709.850 26.560 710.170 26.620 ;
        RECT 761.000 26.080 761.140 26.620 ;
        RECT 811.065 26.620 835.750 26.760 ;
        RECT 811.065 26.575 811.355 26.620 ;
        RECT 835.430 26.560 835.750 26.620 ;
        RECT 811.065 26.080 811.355 26.125 ;
        RECT 761.000 25.940 811.355 26.080 ;
        RECT 811.065 25.895 811.355 25.940 ;
        RECT 276.545 22.340 276.835 22.385 ;
        RECT 323.465 22.340 323.755 22.385 ;
        RECT 276.545 22.200 323.755 22.340 ;
        RECT 276.545 22.155 276.835 22.200 ;
        RECT 323.465 22.155 323.755 22.200 ;
        RECT 373.145 21.320 373.435 21.365 ;
        RECT 400.745 21.320 401.035 21.365 ;
        RECT 373.145 21.180 401.035 21.320 ;
        RECT 373.145 21.135 373.435 21.180 ;
        RECT 400.745 21.135 401.035 21.180 ;
      LAYER via ;
        RECT 169.380 26.560 169.640 26.820 ;
        RECT 469.300 26.560 469.560 26.820 ;
        RECT 517.140 26.560 517.400 26.820 ;
        RECT 565.900 26.560 566.160 26.820 ;
        RECT 613.280 26.560 613.540 26.820 ;
        RECT 662.500 26.560 662.760 26.820 ;
        RECT 709.880 26.560 710.140 26.820 ;
        RECT 835.460 26.560 835.720 26.820 ;
      LAYER met2 ;
        RECT 836.390 1220.330 836.950 1228.680 ;
        RECT 835.520 1220.190 836.950 1220.330 ;
        RECT 169.380 26.530 169.640 26.850 ;
        RECT 469.290 26.675 469.570 27.045 ;
        RECT 517.130 26.675 517.410 27.045 ;
        RECT 565.890 26.675 566.170 27.045 ;
        RECT 613.270 26.675 613.550 27.045 ;
        RECT 662.490 26.675 662.770 27.045 ;
        RECT 709.870 26.675 710.150 27.045 ;
        RECT 835.520 26.850 835.660 1220.190 ;
        RECT 836.390 1219.680 836.950 1220.190 ;
        RECT 469.300 26.530 469.560 26.675 ;
        RECT 517.140 26.530 517.400 26.675 ;
        RECT 565.900 26.530 566.160 26.675 ;
        RECT 613.280 26.530 613.540 26.675 ;
        RECT 662.500 26.530 662.760 26.675 ;
        RECT 709.880 26.530 710.140 26.675 ;
        RECT 835.460 26.530 835.720 26.850 ;
        RECT 169.440 2.400 169.580 26.530 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 469.290 26.720 469.570 27.000 ;
        RECT 517.130 26.720 517.410 27.000 ;
        RECT 565.890 26.720 566.170 27.000 ;
        RECT 613.270 26.720 613.550 27.000 ;
        RECT 662.490 26.720 662.770 27.000 ;
        RECT 709.870 26.720 710.150 27.000 ;
      LAYER met3 ;
        RECT 469.265 27.010 469.595 27.025 ;
        RECT 517.105 27.010 517.435 27.025 ;
        RECT 469.265 26.710 517.435 27.010 ;
        RECT 469.265 26.695 469.595 26.710 ;
        RECT 517.105 26.695 517.435 26.710 ;
        RECT 565.865 27.010 566.195 27.025 ;
        RECT 613.245 27.010 613.575 27.025 ;
        RECT 565.865 26.710 613.575 27.010 ;
        RECT 565.865 26.695 566.195 26.710 ;
        RECT 613.245 26.695 613.575 26.710 ;
        RECT 662.465 27.010 662.795 27.025 ;
        RECT 709.845 27.010 710.175 27.025 ;
        RECT 662.465 26.710 710.175 27.010 ;
        RECT 662.465 26.695 662.795 26.710 ;
        RECT 709.845 26.695 710.175 26.710 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 844.245 620.925 844.415 669.375 ;
        RECT 844.245 531.165 844.415 572.475 ;
        RECT 844.245 476.085 844.415 524.195 ;
        RECT 842.405 282.965 842.575 331.075 ;
        RECT 842.865 186.405 843.035 234.515 ;
      LAYER mcon ;
        RECT 844.245 669.205 844.415 669.375 ;
        RECT 844.245 572.305 844.415 572.475 ;
        RECT 844.245 524.025 844.415 524.195 ;
        RECT 842.405 330.905 842.575 331.075 ;
        RECT 842.865 234.345 843.035 234.515 ;
      LAYER met1 ;
        RECT 843.250 1125.300 843.570 1125.360 ;
        RECT 842.880 1125.160 843.570 1125.300 ;
        RECT 842.880 1124.680 843.020 1125.160 ;
        RECT 843.250 1125.100 843.570 1125.160 ;
        RECT 842.790 1124.420 843.110 1124.680 ;
        RECT 842.790 1110.480 843.110 1110.740 ;
        RECT 842.880 1110.000 843.020 1110.480 ;
        RECT 843.250 1110.000 843.570 1110.060 ;
        RECT 842.880 1109.860 843.570 1110.000 ;
        RECT 843.250 1109.800 843.570 1109.860 ;
        RECT 843.250 966.180 843.570 966.240 ;
        RECT 844.170 966.180 844.490 966.240 ;
        RECT 843.250 966.040 844.490 966.180 ;
        RECT 843.250 965.980 843.570 966.040 ;
        RECT 844.170 965.980 844.490 966.040 ;
        RECT 843.250 869.620 843.570 869.680 ;
        RECT 844.170 869.620 844.490 869.680 ;
        RECT 843.250 869.480 844.490 869.620 ;
        RECT 843.250 869.420 843.570 869.480 ;
        RECT 844.170 869.420 844.490 869.480 ;
        RECT 843.710 670.040 844.030 670.100 ;
        RECT 844.170 670.040 844.490 670.100 ;
        RECT 843.710 669.900 844.490 670.040 ;
        RECT 843.710 669.840 844.030 669.900 ;
        RECT 844.170 669.840 844.490 669.900 ;
        RECT 844.170 669.360 844.490 669.420 ;
        RECT 843.975 669.220 844.490 669.360 ;
        RECT 844.170 669.160 844.490 669.220 ;
        RECT 844.170 621.080 844.490 621.140 ;
        RECT 843.975 620.940 844.490 621.080 ;
        RECT 844.170 620.880 844.490 620.940 ;
        RECT 844.170 579.260 844.490 579.320 ;
        RECT 843.800 579.120 844.490 579.260 ;
        RECT 843.800 578.980 843.940 579.120 ;
        RECT 844.170 579.060 844.490 579.120 ;
        RECT 843.710 578.720 844.030 578.980 ;
        RECT 844.170 572.460 844.490 572.520 ;
        RECT 843.975 572.320 844.490 572.460 ;
        RECT 844.170 572.260 844.490 572.320 ;
        RECT 844.170 531.320 844.490 531.380 ;
        RECT 843.975 531.180 844.490 531.320 ;
        RECT 844.170 531.120 844.490 531.180 ;
        RECT 844.170 524.180 844.490 524.240 ;
        RECT 843.975 524.040 844.490 524.180 ;
        RECT 844.170 523.980 844.490 524.040 ;
        RECT 844.170 476.240 844.490 476.300 ;
        RECT 843.975 476.100 844.490 476.240 ;
        RECT 844.170 476.040 844.490 476.100 ;
        RECT 842.330 458.900 842.650 458.960 ;
        RECT 844.170 458.900 844.490 458.960 ;
        RECT 842.330 458.760 844.490 458.900 ;
        RECT 842.330 458.700 842.650 458.760 ;
        RECT 844.170 458.700 844.490 458.760 ;
        RECT 842.330 386.820 842.650 386.880 ;
        RECT 843.250 386.820 843.570 386.880 ;
        RECT 842.330 386.680 843.570 386.820 ;
        RECT 842.330 386.620 842.650 386.680 ;
        RECT 843.250 386.620 843.570 386.680 ;
        RECT 842.345 331.060 842.635 331.105 ;
        RECT 842.790 331.060 843.110 331.120 ;
        RECT 842.345 330.920 843.110 331.060 ;
        RECT 842.345 330.875 842.635 330.920 ;
        RECT 842.790 330.860 843.110 330.920 ;
        RECT 842.330 283.120 842.650 283.180 ;
        RECT 842.135 282.980 842.650 283.120 ;
        RECT 842.330 282.920 842.650 282.980 ;
        RECT 842.790 234.500 843.110 234.560 ;
        RECT 842.595 234.360 843.110 234.500 ;
        RECT 842.790 234.300 843.110 234.360 ;
        RECT 842.805 186.560 843.095 186.605 ;
        RECT 843.250 186.560 843.570 186.620 ;
        RECT 842.805 186.420 843.570 186.560 ;
        RECT 842.805 186.375 843.095 186.420 ;
        RECT 843.250 186.360 843.570 186.420 ;
        RECT 843.250 158.820 843.570 159.080 ;
        RECT 843.340 158.340 843.480 158.820 ;
        RECT 843.710 158.340 844.030 158.400 ;
        RECT 843.340 158.200 844.030 158.340 ;
        RECT 843.710 158.140 844.030 158.200 ;
        RECT 842.790 137.940 843.110 138.000 ;
        RECT 843.710 137.940 844.030 138.000 ;
        RECT 842.790 137.800 844.030 137.940 ;
        RECT 842.790 137.740 843.110 137.800 ;
        RECT 843.710 137.740 844.030 137.800 ;
        RECT 842.790 62.460 843.110 62.520 ;
        RECT 842.420 62.320 843.110 62.460 ;
        RECT 842.420 62.180 842.560 62.320 ;
        RECT 842.790 62.260 843.110 62.320 ;
        RECT 842.330 61.920 842.650 62.180 ;
      LAYER via ;
        RECT 843.280 1125.100 843.540 1125.360 ;
        RECT 842.820 1124.420 843.080 1124.680 ;
        RECT 842.820 1110.480 843.080 1110.740 ;
        RECT 843.280 1109.800 843.540 1110.060 ;
        RECT 843.280 965.980 843.540 966.240 ;
        RECT 844.200 965.980 844.460 966.240 ;
        RECT 843.280 869.420 843.540 869.680 ;
        RECT 844.200 869.420 844.460 869.680 ;
        RECT 843.740 669.840 844.000 670.100 ;
        RECT 844.200 669.840 844.460 670.100 ;
        RECT 844.200 669.160 844.460 669.420 ;
        RECT 844.200 620.880 844.460 621.140 ;
        RECT 844.200 579.060 844.460 579.320 ;
        RECT 843.740 578.720 844.000 578.980 ;
        RECT 844.200 572.260 844.460 572.520 ;
        RECT 844.200 531.120 844.460 531.380 ;
        RECT 844.200 523.980 844.460 524.240 ;
        RECT 844.200 476.040 844.460 476.300 ;
        RECT 842.360 458.700 842.620 458.960 ;
        RECT 844.200 458.700 844.460 458.960 ;
        RECT 842.360 386.620 842.620 386.880 ;
        RECT 843.280 386.620 843.540 386.880 ;
        RECT 842.820 330.860 843.080 331.120 ;
        RECT 842.360 282.920 842.620 283.180 ;
        RECT 842.820 234.300 843.080 234.560 ;
        RECT 843.280 186.360 843.540 186.620 ;
        RECT 843.280 158.820 843.540 159.080 ;
        RECT 843.740 158.140 844.000 158.400 ;
        RECT 842.820 137.740 843.080 138.000 ;
        RECT 843.740 137.740 844.000 138.000 ;
        RECT 842.820 62.260 843.080 62.520 ;
        RECT 842.360 61.920 842.620 62.180 ;
      LAYER met2 ;
        RECT 845.590 1220.330 846.150 1228.680 ;
        RECT 844.260 1220.190 846.150 1220.330 ;
        RECT 844.260 1196.530 844.400 1220.190 ;
        RECT 845.590 1219.680 846.150 1220.190 ;
        RECT 843.340 1196.390 844.400 1196.530 ;
        RECT 843.340 1125.390 843.480 1196.390 ;
        RECT 843.280 1125.070 843.540 1125.390 ;
        RECT 842.820 1124.390 843.080 1124.710 ;
        RECT 842.880 1110.770 843.020 1124.390 ;
        RECT 842.820 1110.450 843.080 1110.770 ;
        RECT 843.280 1109.770 843.540 1110.090 ;
        RECT 843.340 1027.890 843.480 1109.770 ;
        RECT 842.880 1027.750 843.480 1027.890 ;
        RECT 842.880 1014.405 843.020 1027.750 ;
        RECT 842.810 1014.035 843.090 1014.405 ;
        RECT 844.190 1014.035 844.470 1014.405 ;
        RECT 844.260 966.270 844.400 1014.035 ;
        RECT 843.280 965.950 843.540 966.270 ;
        RECT 844.200 965.950 844.460 966.270 ;
        RECT 843.340 931.330 843.480 965.950 ;
        RECT 842.880 931.190 843.480 931.330 ;
        RECT 842.880 917.845 843.020 931.190 ;
        RECT 842.810 917.475 843.090 917.845 ;
        RECT 844.190 917.475 844.470 917.845 ;
        RECT 844.260 869.710 844.400 917.475 ;
        RECT 843.280 869.390 843.540 869.710 ;
        RECT 844.200 869.390 844.460 869.710 ;
        RECT 843.340 834.770 843.480 869.390 ;
        RECT 842.880 834.630 843.480 834.770 ;
        RECT 842.880 796.690 843.020 834.630 ;
        RECT 842.880 796.550 843.940 796.690 ;
        RECT 843.800 772.890 843.940 796.550 ;
        RECT 843.340 772.750 843.940 772.890 ;
        RECT 843.340 741.610 843.480 772.750 ;
        RECT 842.420 741.470 843.480 741.610 ;
        RECT 842.420 717.925 842.560 741.470 ;
        RECT 842.350 717.555 842.630 717.925 ;
        RECT 844.190 717.555 844.470 717.925 ;
        RECT 844.260 674.290 844.400 717.555 ;
        RECT 843.800 674.150 844.400 674.290 ;
        RECT 843.800 670.130 843.940 674.150 ;
        RECT 843.740 669.810 844.000 670.130 ;
        RECT 844.200 669.810 844.460 670.130 ;
        RECT 844.260 669.450 844.400 669.810 ;
        RECT 844.200 669.130 844.460 669.450 ;
        RECT 844.200 620.850 844.460 621.170 ;
        RECT 844.260 579.350 844.400 620.850 ;
        RECT 844.200 579.030 844.460 579.350 ;
        RECT 843.740 578.690 844.000 579.010 ;
        RECT 843.800 572.970 843.940 578.690 ;
        RECT 843.800 572.830 844.400 572.970 ;
        RECT 844.260 572.550 844.400 572.830 ;
        RECT 844.200 572.230 844.460 572.550 ;
        RECT 844.200 531.090 844.460 531.410 ;
        RECT 844.260 524.270 844.400 531.090 ;
        RECT 844.200 523.950 844.460 524.270 ;
        RECT 844.200 476.010 844.460 476.330 ;
        RECT 844.260 458.990 844.400 476.010 ;
        RECT 842.360 458.670 842.620 458.990 ;
        RECT 844.200 458.670 844.460 458.990 ;
        RECT 842.420 386.910 842.560 458.670 ;
        RECT 842.360 386.590 842.620 386.910 ;
        RECT 843.280 386.590 843.540 386.910 ;
        RECT 843.340 339.165 843.480 386.590 ;
        RECT 843.270 338.795 843.550 339.165 ;
        RECT 842.810 337.945 843.090 338.315 ;
        RECT 842.880 331.150 843.020 337.945 ;
        RECT 842.820 330.830 843.080 331.150 ;
        RECT 842.360 282.890 842.620 283.210 ;
        RECT 842.420 254.730 842.560 282.890 ;
        RECT 842.420 254.590 843.020 254.730 ;
        RECT 842.880 234.590 843.020 254.590 ;
        RECT 842.820 234.270 843.080 234.590 ;
        RECT 843.280 186.330 843.540 186.650 ;
        RECT 843.340 159.110 843.480 186.330 ;
        RECT 843.280 158.790 843.540 159.110 ;
        RECT 843.740 158.110 844.000 158.430 ;
        RECT 843.800 138.030 843.940 158.110 ;
        RECT 842.820 137.710 843.080 138.030 ;
        RECT 843.740 137.710 844.000 138.030 ;
        RECT 842.880 62.550 843.020 137.710 ;
        RECT 842.820 62.230 843.080 62.550 ;
        RECT 842.360 61.890 842.620 62.210 ;
        RECT 842.420 31.125 842.560 61.890 ;
        RECT 186.850 30.755 187.130 31.125 ;
        RECT 842.350 30.755 842.630 31.125 ;
        RECT 186.920 2.400 187.060 30.755 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 842.810 1014.080 843.090 1014.360 ;
        RECT 844.190 1014.080 844.470 1014.360 ;
        RECT 842.810 917.520 843.090 917.800 ;
        RECT 844.190 917.520 844.470 917.800 ;
        RECT 842.350 717.600 842.630 717.880 ;
        RECT 844.190 717.600 844.470 717.880 ;
        RECT 843.270 338.840 843.550 339.120 ;
        RECT 842.810 337.990 843.090 338.270 ;
        RECT 186.850 30.800 187.130 31.080 ;
        RECT 842.350 30.800 842.630 31.080 ;
      LAYER met3 ;
        RECT 842.785 1014.370 843.115 1014.385 ;
        RECT 844.165 1014.370 844.495 1014.385 ;
        RECT 842.785 1014.070 844.495 1014.370 ;
        RECT 842.785 1014.055 843.115 1014.070 ;
        RECT 844.165 1014.055 844.495 1014.070 ;
        RECT 842.785 917.810 843.115 917.825 ;
        RECT 844.165 917.810 844.495 917.825 ;
        RECT 842.785 917.510 844.495 917.810 ;
        RECT 842.785 917.495 843.115 917.510 ;
        RECT 844.165 917.495 844.495 917.510 ;
        RECT 842.325 717.890 842.655 717.905 ;
        RECT 844.165 717.890 844.495 717.905 ;
        RECT 842.325 717.590 844.495 717.890 ;
        RECT 842.325 717.575 842.655 717.590 ;
        RECT 844.165 717.575 844.495 717.590 ;
        RECT 843.245 339.130 843.575 339.145 ;
        RECT 842.110 338.830 843.575 339.130 ;
        RECT 842.110 338.280 842.410 338.830 ;
        RECT 843.245 338.815 843.575 338.830 ;
        RECT 842.785 338.280 843.115 338.295 ;
        RECT 842.110 337.980 843.115 338.280 ;
        RECT 842.785 337.965 843.115 337.980 ;
        RECT 186.825 31.090 187.155 31.105 ;
        RECT 842.325 31.090 842.655 31.105 ;
        RECT 186.825 30.790 842.655 31.090 ;
        RECT 186.825 30.775 187.155 30.790 ;
        RECT 842.325 30.775 842.655 30.790 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 849.765 1110.865 849.935 1135.175 ;
        RECT 848.845 386.325 849.015 434.775 ;
        RECT 849.305 186.405 849.475 234.515 ;
      LAYER mcon ;
        RECT 849.765 1135.005 849.935 1135.175 ;
        RECT 848.845 434.605 849.015 434.775 ;
        RECT 849.305 234.345 849.475 234.515 ;
      LAYER met1 ;
        RECT 849.690 1135.160 850.010 1135.220 ;
        RECT 849.495 1135.020 850.010 1135.160 ;
        RECT 849.690 1134.960 850.010 1135.020 ;
        RECT 849.705 1111.020 849.995 1111.065 ;
        RECT 850.150 1111.020 850.470 1111.080 ;
        RECT 849.705 1110.880 850.470 1111.020 ;
        RECT 849.705 1110.835 849.995 1110.880 ;
        RECT 850.150 1110.820 850.470 1110.880 ;
        RECT 850.150 1062.740 850.470 1062.800 ;
        RECT 850.610 1062.740 850.930 1062.800 ;
        RECT 850.150 1062.600 850.930 1062.740 ;
        RECT 850.150 1062.540 850.470 1062.600 ;
        RECT 850.610 1062.540 850.930 1062.600 ;
        RECT 848.770 966.180 849.090 966.240 ;
        RECT 850.150 966.180 850.470 966.240 ;
        RECT 848.770 966.040 850.470 966.180 ;
        RECT 848.770 965.980 849.090 966.040 ;
        RECT 850.150 965.980 850.470 966.040 ;
        RECT 848.770 869.620 849.090 869.680 ;
        RECT 850.150 869.620 850.470 869.680 ;
        RECT 848.770 869.480 850.470 869.620 ;
        RECT 848.770 869.420 849.090 869.480 ;
        RECT 850.150 869.420 850.470 869.480 ;
        RECT 849.690 821.000 850.010 821.060 ;
        RECT 850.150 821.000 850.470 821.060 ;
        RECT 849.690 820.860 850.470 821.000 ;
        RECT 849.690 820.800 850.010 820.860 ;
        RECT 850.150 820.800 850.470 820.860 ;
        RECT 848.785 434.760 849.075 434.805 ;
        RECT 849.230 434.760 849.550 434.820 ;
        RECT 848.785 434.620 849.550 434.760 ;
        RECT 848.785 434.575 849.075 434.620 ;
        RECT 849.230 434.560 849.550 434.620 ;
        RECT 848.770 386.480 849.090 386.540 ;
        RECT 848.575 386.340 849.090 386.480 ;
        RECT 848.770 386.280 849.090 386.340 ;
        RECT 849.230 303.520 849.550 303.580 ;
        RECT 850.150 303.520 850.470 303.580 ;
        RECT 849.230 303.380 850.470 303.520 ;
        RECT 849.230 303.320 849.550 303.380 ;
        RECT 850.150 303.320 850.470 303.380 ;
        RECT 849.230 234.500 849.550 234.560 ;
        RECT 849.035 234.360 849.550 234.500 ;
        RECT 849.230 234.300 849.550 234.360 ;
        RECT 849.245 186.560 849.535 186.605 ;
        RECT 849.690 186.560 850.010 186.620 ;
        RECT 849.245 186.420 850.010 186.560 ;
        RECT 849.245 186.375 849.535 186.420 ;
        RECT 849.690 186.360 850.010 186.420 ;
        RECT 849.690 158.820 850.010 159.080 ;
        RECT 849.780 158.400 849.920 158.820 ;
        RECT 849.690 158.140 850.010 158.400 ;
        RECT 849.230 48.520 849.550 48.580 ;
        RECT 850.610 48.520 850.930 48.580 ;
        RECT 849.230 48.380 850.930 48.520 ;
        RECT 849.230 48.320 849.550 48.380 ;
        RECT 850.610 48.320 850.930 48.380 ;
        RECT 204.770 32.200 205.090 32.260 ;
        RECT 849.230 32.200 849.550 32.260 ;
        RECT 204.770 32.060 849.550 32.200 ;
        RECT 204.770 32.000 205.090 32.060 ;
        RECT 849.230 32.000 849.550 32.060 ;
      LAYER via ;
        RECT 849.720 1134.960 849.980 1135.220 ;
        RECT 850.180 1110.820 850.440 1111.080 ;
        RECT 850.180 1062.540 850.440 1062.800 ;
        RECT 850.640 1062.540 850.900 1062.800 ;
        RECT 848.800 965.980 849.060 966.240 ;
        RECT 850.180 965.980 850.440 966.240 ;
        RECT 848.800 869.420 849.060 869.680 ;
        RECT 850.180 869.420 850.440 869.680 ;
        RECT 849.720 820.800 849.980 821.060 ;
        RECT 850.180 820.800 850.440 821.060 ;
        RECT 849.260 434.560 849.520 434.820 ;
        RECT 848.800 386.280 849.060 386.540 ;
        RECT 849.260 303.320 849.520 303.580 ;
        RECT 850.180 303.320 850.440 303.580 ;
        RECT 849.260 234.300 849.520 234.560 ;
        RECT 849.720 186.360 849.980 186.620 ;
        RECT 849.720 158.820 849.980 159.080 ;
        RECT 849.720 158.140 849.980 158.400 ;
        RECT 849.260 48.320 849.520 48.580 ;
        RECT 850.640 48.320 850.900 48.580 ;
        RECT 204.800 32.000 205.060 32.260 ;
        RECT 849.260 32.000 849.520 32.260 ;
      LAYER met2 ;
        RECT 854.790 1220.330 855.350 1228.680 ;
        RECT 853.460 1220.190 855.350 1220.330 ;
        RECT 853.460 1196.530 853.600 1220.190 ;
        RECT 854.790 1219.680 855.350 1220.190 ;
        RECT 849.780 1196.390 853.600 1196.530 ;
        RECT 849.780 1135.250 849.920 1196.390 ;
        RECT 849.720 1134.930 849.980 1135.250 ;
        RECT 850.240 1111.110 850.380 1111.265 ;
        RECT 850.180 1110.850 850.440 1111.110 ;
        RECT 850.180 1110.790 850.840 1110.850 ;
        RECT 850.240 1110.710 850.840 1110.790 ;
        RECT 850.700 1062.830 850.840 1110.710 ;
        RECT 850.180 1062.510 850.440 1062.830 ;
        RECT 850.640 1062.510 850.900 1062.830 ;
        RECT 850.240 1027.890 850.380 1062.510 ;
        RECT 849.780 1027.750 850.380 1027.890 ;
        RECT 849.780 1014.405 849.920 1027.750 ;
        RECT 848.790 1014.035 849.070 1014.405 ;
        RECT 849.710 1014.035 849.990 1014.405 ;
        RECT 848.860 966.270 849.000 1014.035 ;
        RECT 848.800 965.950 849.060 966.270 ;
        RECT 850.180 965.950 850.440 966.270 ;
        RECT 850.240 931.330 850.380 965.950 ;
        RECT 849.780 931.190 850.380 931.330 ;
        RECT 849.780 917.845 849.920 931.190 ;
        RECT 848.790 917.475 849.070 917.845 ;
        RECT 849.710 917.475 849.990 917.845 ;
        RECT 848.860 869.710 849.000 917.475 ;
        RECT 848.800 869.390 849.060 869.710 ;
        RECT 850.180 869.390 850.440 869.710 ;
        RECT 850.240 834.770 850.380 869.390 ;
        RECT 849.780 834.630 850.380 834.770 ;
        RECT 849.780 821.090 849.920 834.630 ;
        RECT 849.720 820.770 849.980 821.090 ;
        RECT 850.180 820.770 850.440 821.090 ;
        RECT 850.240 738.210 850.380 820.770 ;
        RECT 849.780 738.070 850.380 738.210 ;
        RECT 849.780 724.440 849.920 738.070 ;
        RECT 848.860 724.300 849.920 724.440 ;
        RECT 848.860 676.445 849.000 724.300 ;
        RECT 848.790 676.075 849.070 676.445 ;
        RECT 850.170 676.075 850.450 676.445 ;
        RECT 850.240 641.650 850.380 676.075 ;
        RECT 849.780 641.510 850.380 641.650 ;
        RECT 849.780 627.880 849.920 641.510 ;
        RECT 848.860 627.740 849.920 627.880 ;
        RECT 848.860 579.885 849.000 627.740 ;
        RECT 848.790 579.515 849.070 579.885 ;
        RECT 850.170 579.515 850.450 579.885 ;
        RECT 850.240 545.090 850.380 579.515 ;
        RECT 849.780 544.950 850.380 545.090 ;
        RECT 849.780 531.320 849.920 544.950 ;
        RECT 848.860 531.180 849.920 531.320 ;
        RECT 848.860 483.325 849.000 531.180 ;
        RECT 848.790 482.955 849.070 483.325 ;
        RECT 850.170 482.955 850.450 483.325 ;
        RECT 850.240 448.530 850.380 482.955 ;
        RECT 849.320 448.390 850.380 448.530 ;
        RECT 849.320 434.850 849.460 448.390 ;
        RECT 849.260 434.530 849.520 434.850 ;
        RECT 848.800 386.250 849.060 386.570 ;
        RECT 848.860 351.290 849.000 386.250 ;
        RECT 848.860 351.150 849.460 351.290 ;
        RECT 849.320 303.610 849.460 351.150 ;
        RECT 849.260 303.290 849.520 303.610 ;
        RECT 850.180 303.290 850.440 303.610 ;
        RECT 850.240 241.640 850.380 303.290 ;
        RECT 849.320 241.500 850.380 241.640 ;
        RECT 849.320 234.590 849.460 241.500 ;
        RECT 849.260 234.270 849.520 234.590 ;
        RECT 849.720 186.330 849.980 186.650 ;
        RECT 849.780 159.110 849.920 186.330 ;
        RECT 849.720 158.790 849.980 159.110 ;
        RECT 849.720 158.110 849.980 158.430 ;
        RECT 849.780 137.770 849.920 158.110 ;
        RECT 849.780 137.630 850.840 137.770 ;
        RECT 850.700 48.610 850.840 137.630 ;
        RECT 849.260 48.290 849.520 48.610 ;
        RECT 850.640 48.290 850.900 48.610 ;
        RECT 849.320 32.290 849.460 48.290 ;
        RECT 204.800 31.970 205.060 32.290 ;
        RECT 849.260 31.970 849.520 32.290 ;
        RECT 204.860 2.400 205.000 31.970 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 848.790 1014.080 849.070 1014.360 ;
        RECT 849.710 1014.080 849.990 1014.360 ;
        RECT 848.790 917.520 849.070 917.800 ;
        RECT 849.710 917.520 849.990 917.800 ;
        RECT 848.790 676.120 849.070 676.400 ;
        RECT 850.170 676.120 850.450 676.400 ;
        RECT 848.790 579.560 849.070 579.840 ;
        RECT 850.170 579.560 850.450 579.840 ;
        RECT 848.790 483.000 849.070 483.280 ;
        RECT 850.170 483.000 850.450 483.280 ;
      LAYER met3 ;
        RECT 848.765 1014.370 849.095 1014.385 ;
        RECT 849.685 1014.370 850.015 1014.385 ;
        RECT 848.765 1014.070 850.015 1014.370 ;
        RECT 848.765 1014.055 849.095 1014.070 ;
        RECT 849.685 1014.055 850.015 1014.070 ;
        RECT 848.765 917.810 849.095 917.825 ;
        RECT 849.685 917.810 850.015 917.825 ;
        RECT 848.765 917.510 850.015 917.810 ;
        RECT 848.765 917.495 849.095 917.510 ;
        RECT 849.685 917.495 850.015 917.510 ;
        RECT 848.765 676.410 849.095 676.425 ;
        RECT 850.145 676.410 850.475 676.425 ;
        RECT 848.765 676.110 850.475 676.410 ;
        RECT 848.765 676.095 849.095 676.110 ;
        RECT 850.145 676.095 850.475 676.110 ;
        RECT 848.765 579.850 849.095 579.865 ;
        RECT 850.145 579.850 850.475 579.865 ;
        RECT 848.765 579.550 850.475 579.850 ;
        RECT 848.765 579.535 849.095 579.550 ;
        RECT 850.145 579.535 850.475 579.550 ;
        RECT 848.765 483.290 849.095 483.305 ;
        RECT 850.145 483.290 850.475 483.305 ;
        RECT 848.765 482.990 850.475 483.290 ;
        RECT 848.765 482.975 849.095 482.990 ;
        RECT 850.145 482.975 850.475 482.990 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.990 1220.330 864.550 1228.680 ;
        RECT 863.120 1220.190 864.550 1220.330 ;
        RECT 863.120 31.805 863.260 1220.190 ;
        RECT 863.990 1219.680 864.550 1220.190 ;
        RECT 222.730 31.435 223.010 31.805 ;
        RECT 863.050 31.435 863.330 31.805 ;
        RECT 222.800 2.400 222.940 31.435 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 222.730 31.480 223.010 31.760 ;
        RECT 863.050 31.480 863.330 31.760 ;
      LAYER met3 ;
        RECT 222.705 31.770 223.035 31.785 ;
        RECT 863.025 31.770 863.355 31.785 ;
        RECT 222.705 31.470 863.355 31.770 ;
        RECT 222.705 31.455 223.035 31.470 ;
        RECT 863.025 31.455 863.355 31.470 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 30.840 20.630 30.900 ;
        RECT 759.530 30.840 759.850 30.900 ;
        RECT 20.310 30.700 759.850 30.840 ;
        RECT 20.310 30.640 20.630 30.700 ;
        RECT 759.530 30.640 759.850 30.700 ;
      LAYER via ;
        RECT 20.340 30.640 20.600 30.900 ;
        RECT 759.560 30.640 759.820 30.900 ;
      LAYER met2 ;
        RECT 760.030 1220.330 760.590 1228.680 ;
        RECT 759.620 1220.190 760.590 1220.330 ;
        RECT 759.620 30.930 759.760 1220.190 ;
        RECT 760.030 1219.680 760.590 1220.190 ;
        RECT 20.340 30.610 20.600 30.930 ;
        RECT 759.560 30.610 759.820 30.930 ;
        RECT 20.400 2.400 20.540 30.610 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 766.965 620.925 767.135 669.375 ;
        RECT 766.505 524.365 766.675 572.135 ;
      LAYER mcon ;
        RECT 766.965 669.205 767.135 669.375 ;
        RECT 766.505 571.965 766.675 572.135 ;
      LAYER met1 ;
        RECT 766.890 669.360 767.210 669.420 ;
        RECT 766.695 669.220 767.210 669.360 ;
        RECT 766.890 669.160 767.210 669.220 ;
        RECT 766.890 621.080 767.210 621.140 ;
        RECT 766.695 620.940 767.210 621.080 ;
        RECT 766.890 620.880 767.210 620.940 ;
        RECT 767.350 572.940 767.670 573.200 ;
        RECT 766.430 572.800 766.750 572.860 ;
        RECT 767.440 572.800 767.580 572.940 ;
        RECT 766.430 572.660 767.580 572.800 ;
        RECT 766.430 572.600 766.750 572.660 ;
        RECT 766.430 572.120 766.750 572.180 ;
        RECT 766.235 571.980 766.750 572.120 ;
        RECT 766.430 571.920 766.750 571.980 ;
        RECT 766.445 524.520 766.735 524.565 ;
        RECT 766.890 524.520 767.210 524.580 ;
        RECT 766.445 524.380 767.210 524.520 ;
        RECT 766.445 524.335 766.735 524.380 ;
        RECT 766.890 524.320 767.210 524.380 ;
        RECT 766.890 497.120 767.210 497.380 ;
        RECT 766.980 496.700 767.120 497.120 ;
        RECT 766.890 496.440 767.210 496.700 ;
        RECT 44.230 31.180 44.550 31.240 ;
        RECT 766.890 31.180 767.210 31.240 ;
        RECT 44.230 31.040 767.210 31.180 ;
        RECT 44.230 30.980 44.550 31.040 ;
        RECT 766.890 30.980 767.210 31.040 ;
      LAYER via ;
        RECT 766.920 669.160 767.180 669.420 ;
        RECT 766.920 620.880 767.180 621.140 ;
        RECT 767.380 572.940 767.640 573.200 ;
        RECT 766.460 572.600 766.720 572.860 ;
        RECT 766.460 571.920 766.720 572.180 ;
        RECT 766.920 524.320 767.180 524.580 ;
        RECT 766.920 497.120 767.180 497.380 ;
        RECT 766.920 496.440 767.180 496.700 ;
        RECT 44.260 30.980 44.520 31.240 ;
        RECT 766.920 30.980 767.180 31.240 ;
      LAYER met2 ;
        RECT 772.450 1220.330 773.010 1228.680 ;
        RECT 770.200 1220.190 773.010 1220.330 ;
        RECT 770.200 1184.970 770.340 1220.190 ;
        RECT 772.450 1219.680 773.010 1220.190 ;
        RECT 766.980 1184.830 770.340 1184.970 ;
        RECT 766.980 1104.165 767.120 1184.830 ;
        RECT 766.910 1103.795 767.190 1104.165 ;
        RECT 767.830 1103.795 768.110 1104.165 ;
        RECT 767.900 1061.210 768.040 1103.795 ;
        RECT 766.980 1061.070 768.040 1061.210 ;
        RECT 766.980 1038.770 767.120 1061.070 ;
        RECT 766.520 1038.630 767.120 1038.770 ;
        RECT 766.520 979.610 766.660 1038.630 ;
        RECT 766.520 979.470 767.120 979.610 ;
        RECT 766.980 883.730 767.120 979.470 ;
        RECT 766.520 883.590 767.120 883.730 ;
        RECT 766.520 883.050 766.660 883.590 ;
        RECT 766.520 882.910 767.120 883.050 ;
        RECT 766.980 787.170 767.120 882.910 ;
        RECT 766.520 787.030 767.120 787.170 ;
        RECT 766.520 786.490 766.660 787.030 ;
        RECT 766.520 786.350 767.120 786.490 ;
        RECT 766.980 689.930 767.120 786.350 ;
        RECT 766.980 689.790 768.040 689.930 ;
        RECT 767.900 669.645 768.040 689.790 ;
        RECT 766.910 669.275 767.190 669.645 ;
        RECT 767.830 669.275 768.110 669.645 ;
        RECT 766.920 669.130 767.180 669.275 ;
        RECT 766.920 620.850 767.180 621.170 ;
        RECT 766.980 594.050 767.120 620.850 ;
        RECT 766.980 593.910 767.580 594.050 ;
        RECT 767.440 573.230 767.580 593.910 ;
        RECT 767.380 572.910 767.640 573.230 ;
        RECT 766.460 572.570 766.720 572.890 ;
        RECT 766.520 572.210 766.660 572.570 ;
        RECT 766.460 571.890 766.720 572.210 ;
        RECT 766.920 524.290 767.180 524.610 ;
        RECT 766.980 497.410 767.120 524.290 ;
        RECT 766.920 497.090 767.180 497.410 ;
        RECT 766.920 496.410 767.180 496.730 ;
        RECT 766.980 31.270 767.120 496.410 ;
        RECT 44.260 30.950 44.520 31.270 ;
        RECT 766.920 30.950 767.180 31.270 ;
        RECT 44.320 2.400 44.460 30.950 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 766.910 1103.840 767.190 1104.120 ;
        RECT 767.830 1103.840 768.110 1104.120 ;
        RECT 766.910 669.320 767.190 669.600 ;
        RECT 767.830 669.320 768.110 669.600 ;
      LAYER met3 ;
        RECT 766.885 1104.130 767.215 1104.145 ;
        RECT 767.805 1104.130 768.135 1104.145 ;
        RECT 766.885 1103.830 768.135 1104.130 ;
        RECT 766.885 1103.815 767.215 1103.830 ;
        RECT 767.805 1103.815 768.135 1103.830 ;
        RECT 766.885 669.610 767.215 669.625 ;
        RECT 767.805 669.610 768.135 669.625 ;
        RECT 766.885 669.310 768.135 669.610 ;
        RECT 766.885 669.295 767.215 669.310 ;
        RECT 767.805 669.295 768.135 669.310 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 32.540 246.950 32.600 ;
        RECT 876.370 32.540 876.690 32.600 ;
        RECT 246.630 32.400 876.690 32.540 ;
        RECT 246.630 32.340 246.950 32.400 ;
        RECT 876.370 32.340 876.690 32.400 ;
      LAYER via ;
        RECT 246.660 32.340 246.920 32.600 ;
        RECT 876.400 32.340 876.660 32.600 ;
      LAYER met2 ;
        RECT 876.410 1220.330 876.970 1228.680 ;
        RECT 876.410 1219.680 877.060 1220.330 ;
        RECT 876.920 33.050 877.060 1219.680 ;
        RECT 876.460 32.910 877.060 33.050 ;
        RECT 876.460 32.630 876.600 32.910 ;
        RECT 246.660 32.310 246.920 32.630 ;
        RECT 876.400 32.310 876.660 32.630 ;
        RECT 246.720 2.400 246.860 32.310 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 32.880 264.430 32.940 ;
        RECT 883.730 32.880 884.050 32.940 ;
        RECT 264.110 32.740 884.050 32.880 ;
        RECT 264.110 32.680 264.430 32.740 ;
        RECT 883.730 32.680 884.050 32.740 ;
      LAYER via ;
        RECT 264.140 32.680 264.400 32.940 ;
        RECT 883.760 32.680 884.020 32.940 ;
      LAYER met2 ;
        RECT 885.610 1220.330 886.170 1228.680 ;
        RECT 883.820 1220.190 886.170 1220.330 ;
        RECT 883.820 32.970 883.960 1220.190 ;
        RECT 885.610 1219.680 886.170 1220.190 ;
        RECT 264.140 32.650 264.400 32.970 ;
        RECT 883.760 32.650 884.020 32.970 ;
        RECT 264.200 2.400 264.340 32.650 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 891.165 1062.585 891.335 1076.355 ;
        RECT 891.165 579.785 891.335 627.895 ;
        RECT 891.165 483.225 891.335 531.335 ;
        RECT 891.165 386.325 891.335 434.775 ;
        RECT 891.165 241.485 891.335 289.595 ;
      LAYER mcon ;
        RECT 891.165 1076.185 891.335 1076.355 ;
        RECT 891.165 627.725 891.335 627.895 ;
        RECT 891.165 531.165 891.335 531.335 ;
        RECT 891.165 434.605 891.335 434.775 ;
        RECT 891.165 289.425 891.335 289.595 ;
      LAYER met1 ;
        RECT 891.090 1076.340 891.410 1076.400 ;
        RECT 890.895 1076.200 891.410 1076.340 ;
        RECT 891.090 1076.140 891.410 1076.200 ;
        RECT 891.090 1062.740 891.410 1062.800 ;
        RECT 890.895 1062.600 891.410 1062.740 ;
        RECT 891.090 1062.540 891.410 1062.600 ;
        RECT 891.090 966.180 891.410 966.240 ;
        RECT 892.010 966.180 892.330 966.240 ;
        RECT 891.090 966.040 892.330 966.180 ;
        RECT 891.090 965.980 891.410 966.040 ;
        RECT 892.010 965.980 892.330 966.040 ;
        RECT 891.090 869.620 891.410 869.680 ;
        RECT 892.010 869.620 892.330 869.680 ;
        RECT 891.090 869.480 892.330 869.620 ;
        RECT 891.090 869.420 891.410 869.480 ;
        RECT 892.010 869.420 892.330 869.480 ;
        RECT 891.090 821.000 891.410 821.060 ;
        RECT 892.010 821.000 892.330 821.060 ;
        RECT 891.090 820.860 892.330 821.000 ;
        RECT 891.090 820.800 891.410 820.860 ;
        RECT 892.010 820.800 892.330 820.860 ;
        RECT 891.090 724.440 891.410 724.500 ;
        RECT 892.010 724.440 892.330 724.500 ;
        RECT 891.090 724.300 892.330 724.440 ;
        RECT 891.090 724.240 891.410 724.300 ;
        RECT 892.010 724.240 892.330 724.300 ;
        RECT 891.090 627.880 891.410 627.940 ;
        RECT 890.895 627.740 891.410 627.880 ;
        RECT 891.090 627.680 891.410 627.740 ;
        RECT 891.090 579.940 891.410 580.000 ;
        RECT 890.895 579.800 891.410 579.940 ;
        RECT 891.090 579.740 891.410 579.800 ;
        RECT 891.090 531.320 891.410 531.380 ;
        RECT 890.895 531.180 891.410 531.320 ;
        RECT 891.090 531.120 891.410 531.180 ;
        RECT 891.090 483.380 891.410 483.440 ;
        RECT 890.895 483.240 891.410 483.380 ;
        RECT 891.090 483.180 891.410 483.240 ;
        RECT 891.090 434.760 891.410 434.820 ;
        RECT 890.895 434.620 891.410 434.760 ;
        RECT 891.090 434.560 891.410 434.620 ;
        RECT 891.090 386.480 891.410 386.540 ;
        RECT 890.895 386.340 891.410 386.480 ;
        RECT 891.090 386.280 891.410 386.340 ;
        RECT 889.710 314.060 890.030 314.120 ;
        RECT 891.090 314.060 891.410 314.120 ;
        RECT 889.710 313.920 891.410 314.060 ;
        RECT 889.710 313.860 890.030 313.920 ;
        RECT 891.090 313.860 891.410 313.920 ;
        RECT 891.090 289.580 891.410 289.640 ;
        RECT 890.895 289.440 891.410 289.580 ;
        RECT 891.090 289.380 891.410 289.440 ;
        RECT 891.105 241.640 891.395 241.685 ;
        RECT 891.550 241.640 891.870 241.700 ;
        RECT 891.105 241.500 891.870 241.640 ;
        RECT 891.105 241.455 891.395 241.500 ;
        RECT 891.550 241.440 891.870 241.500 ;
        RECT 890.630 206.960 890.950 207.020 ;
        RECT 891.550 206.960 891.870 207.020 ;
        RECT 890.630 206.820 891.870 206.960 ;
        RECT 890.630 206.760 890.950 206.820 ;
        RECT 891.550 206.760 891.870 206.820 ;
        RECT 891.550 156.100 891.870 156.360 ;
        RECT 891.640 155.680 891.780 156.100 ;
        RECT 891.550 155.420 891.870 155.680 ;
        RECT 282.050 33.220 282.370 33.280 ;
        RECT 891.090 33.220 891.410 33.280 ;
        RECT 282.050 33.080 891.410 33.220 ;
        RECT 282.050 33.020 282.370 33.080 ;
        RECT 891.090 33.020 891.410 33.080 ;
      LAYER via ;
        RECT 891.120 1076.140 891.380 1076.400 ;
        RECT 891.120 1062.540 891.380 1062.800 ;
        RECT 891.120 965.980 891.380 966.240 ;
        RECT 892.040 965.980 892.300 966.240 ;
        RECT 891.120 869.420 891.380 869.680 ;
        RECT 892.040 869.420 892.300 869.680 ;
        RECT 891.120 820.800 891.380 821.060 ;
        RECT 892.040 820.800 892.300 821.060 ;
        RECT 891.120 724.240 891.380 724.500 ;
        RECT 892.040 724.240 892.300 724.500 ;
        RECT 891.120 627.680 891.380 627.940 ;
        RECT 891.120 579.740 891.380 580.000 ;
        RECT 891.120 531.120 891.380 531.380 ;
        RECT 891.120 483.180 891.380 483.440 ;
        RECT 891.120 434.560 891.380 434.820 ;
        RECT 891.120 386.280 891.380 386.540 ;
        RECT 889.740 313.860 890.000 314.120 ;
        RECT 891.120 313.860 891.380 314.120 ;
        RECT 891.120 289.380 891.380 289.640 ;
        RECT 891.580 241.440 891.840 241.700 ;
        RECT 890.660 206.760 890.920 207.020 ;
        RECT 891.580 206.760 891.840 207.020 ;
        RECT 891.580 156.100 891.840 156.360 ;
        RECT 891.580 155.420 891.840 155.680 ;
        RECT 282.080 33.020 282.340 33.280 ;
        RECT 891.120 33.020 891.380 33.280 ;
      LAYER met2 ;
        RECT 894.810 1221.010 895.370 1228.680 ;
        RECT 892.560 1220.870 895.370 1221.010 ;
        RECT 892.560 1196.530 892.700 1220.870 ;
        RECT 894.810 1219.680 895.370 1220.870 ;
        RECT 891.180 1196.390 892.700 1196.530 ;
        RECT 891.180 1076.430 891.320 1196.390 ;
        RECT 891.120 1076.110 891.380 1076.430 ;
        RECT 891.120 1062.510 891.380 1062.830 ;
        RECT 891.180 1014.405 891.320 1062.510 ;
        RECT 891.110 1014.035 891.390 1014.405 ;
        RECT 892.030 1014.035 892.310 1014.405 ;
        RECT 892.100 966.270 892.240 1014.035 ;
        RECT 891.120 965.950 891.380 966.270 ;
        RECT 892.040 965.950 892.300 966.270 ;
        RECT 891.180 917.845 891.320 965.950 ;
        RECT 891.110 917.475 891.390 917.845 ;
        RECT 892.030 917.475 892.310 917.845 ;
        RECT 892.100 869.710 892.240 917.475 ;
        RECT 891.120 869.390 891.380 869.710 ;
        RECT 892.040 869.390 892.300 869.710 ;
        RECT 891.180 821.090 891.320 869.390 ;
        RECT 891.120 820.770 891.380 821.090 ;
        RECT 892.040 820.770 892.300 821.090 ;
        RECT 892.100 773.005 892.240 820.770 ;
        RECT 891.110 772.635 891.390 773.005 ;
        RECT 892.030 772.635 892.310 773.005 ;
        RECT 891.180 724.530 891.320 772.635 ;
        RECT 891.120 724.210 891.380 724.530 ;
        RECT 892.040 724.210 892.300 724.530 ;
        RECT 892.100 676.445 892.240 724.210 ;
        RECT 891.110 676.075 891.390 676.445 ;
        RECT 892.030 676.075 892.310 676.445 ;
        RECT 891.180 627.970 891.320 676.075 ;
        RECT 891.120 627.650 891.380 627.970 ;
        RECT 891.120 579.710 891.380 580.030 ;
        RECT 891.180 531.410 891.320 579.710 ;
        RECT 891.120 531.090 891.380 531.410 ;
        RECT 891.120 483.150 891.380 483.470 ;
        RECT 891.180 434.850 891.320 483.150 ;
        RECT 891.120 434.530 891.380 434.850 ;
        RECT 891.120 386.250 891.380 386.570 ;
        RECT 891.180 314.150 891.320 386.250 ;
        RECT 889.740 313.830 890.000 314.150 ;
        RECT 891.120 313.830 891.380 314.150 ;
        RECT 889.800 290.205 889.940 313.830 ;
        RECT 889.730 289.835 890.010 290.205 ;
        RECT 890.650 290.090 890.930 290.205 ;
        RECT 890.650 289.950 891.320 290.090 ;
        RECT 890.650 289.835 890.930 289.950 ;
        RECT 891.180 289.670 891.320 289.950 ;
        RECT 891.120 289.350 891.380 289.670 ;
        RECT 891.580 241.410 891.840 241.730 ;
        RECT 891.640 207.130 891.780 241.410 ;
        RECT 890.720 207.050 891.780 207.130 ;
        RECT 890.660 206.990 891.840 207.050 ;
        RECT 890.660 206.730 890.920 206.990 ;
        RECT 891.580 206.730 891.840 206.990 ;
        RECT 891.640 156.390 891.780 206.730 ;
        RECT 891.580 156.070 891.840 156.390 ;
        RECT 891.580 155.390 891.840 155.710 ;
        RECT 891.640 111.250 891.780 155.390 ;
        RECT 891.180 111.110 891.780 111.250 ;
        RECT 891.180 110.570 891.320 111.110 ;
        RECT 890.720 110.430 891.320 110.570 ;
        RECT 890.720 109.890 890.860 110.430 ;
        RECT 890.720 109.750 891.320 109.890 ;
        RECT 891.180 33.310 891.320 109.750 ;
        RECT 282.080 32.990 282.340 33.310 ;
        RECT 891.120 32.990 891.380 33.310 ;
        RECT 282.140 2.400 282.280 32.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 891.110 1014.080 891.390 1014.360 ;
        RECT 892.030 1014.080 892.310 1014.360 ;
        RECT 891.110 917.520 891.390 917.800 ;
        RECT 892.030 917.520 892.310 917.800 ;
        RECT 891.110 772.680 891.390 772.960 ;
        RECT 892.030 772.680 892.310 772.960 ;
        RECT 891.110 676.120 891.390 676.400 ;
        RECT 892.030 676.120 892.310 676.400 ;
        RECT 889.730 289.880 890.010 290.160 ;
        RECT 890.650 289.880 890.930 290.160 ;
      LAYER met3 ;
        RECT 891.085 1014.370 891.415 1014.385 ;
        RECT 892.005 1014.370 892.335 1014.385 ;
        RECT 891.085 1014.070 892.335 1014.370 ;
        RECT 891.085 1014.055 891.415 1014.070 ;
        RECT 892.005 1014.055 892.335 1014.070 ;
        RECT 891.085 917.810 891.415 917.825 ;
        RECT 892.005 917.810 892.335 917.825 ;
        RECT 891.085 917.510 892.335 917.810 ;
        RECT 891.085 917.495 891.415 917.510 ;
        RECT 892.005 917.495 892.335 917.510 ;
        RECT 891.085 772.970 891.415 772.985 ;
        RECT 892.005 772.970 892.335 772.985 ;
        RECT 891.085 772.670 892.335 772.970 ;
        RECT 891.085 772.655 891.415 772.670 ;
        RECT 892.005 772.655 892.335 772.670 ;
        RECT 891.085 676.410 891.415 676.425 ;
        RECT 892.005 676.410 892.335 676.425 ;
        RECT 891.085 676.110 892.335 676.410 ;
        RECT 891.085 676.095 891.415 676.110 ;
        RECT 892.005 676.095 892.335 676.110 ;
        RECT 889.705 290.170 890.035 290.185 ;
        RECT 890.625 290.170 890.955 290.185 ;
        RECT 889.705 289.870 890.955 290.170 ;
        RECT 889.705 289.855 890.035 289.870 ;
        RECT 890.625 289.855 890.955 289.870 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 33.560 300.310 33.620 ;
        RECT 904.430 33.560 904.750 33.620 ;
        RECT 299.990 33.420 904.750 33.560 ;
        RECT 299.990 33.360 300.310 33.420 ;
        RECT 904.430 33.360 904.750 33.420 ;
      LAYER via ;
        RECT 300.020 33.360 300.280 33.620 ;
        RECT 904.460 33.360 904.720 33.620 ;
      LAYER met2 ;
        RECT 904.010 1220.330 904.570 1228.680 ;
        RECT 904.010 1219.680 904.660 1220.330 ;
        RECT 904.520 33.650 904.660 1219.680 ;
        RECT 300.020 33.330 300.280 33.650 ;
        RECT 904.460 33.330 904.720 33.650 ;
        RECT 300.080 2.400 300.220 33.330 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 33.900 318.250 33.960 ;
        RECT 911.330 33.900 911.650 33.960 ;
        RECT 317.930 33.760 911.650 33.900 ;
        RECT 317.930 33.700 318.250 33.760 ;
        RECT 911.330 33.700 911.650 33.760 ;
      LAYER via ;
        RECT 317.960 33.700 318.220 33.960 ;
        RECT 911.360 33.700 911.620 33.960 ;
      LAYER met2 ;
        RECT 913.210 1220.330 913.770 1228.680 ;
        RECT 911.420 1220.190 913.770 1220.330 ;
        RECT 911.420 33.990 911.560 1220.190 ;
        RECT 913.210 1219.680 913.770 1220.190 ;
        RECT 317.960 33.670 318.220 33.990 ;
        RECT 911.360 33.670 911.620 33.990 ;
        RECT 318.020 2.400 318.160 33.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 34.240 336.190 34.300 ;
        RECT 918.690 34.240 919.010 34.300 ;
        RECT 335.870 34.100 919.010 34.240 ;
        RECT 335.870 34.040 336.190 34.100 ;
        RECT 918.690 34.040 919.010 34.100 ;
      LAYER via ;
        RECT 335.900 34.040 336.160 34.300 ;
        RECT 918.720 34.040 918.980 34.300 ;
      LAYER met2 ;
        RECT 921.950 1220.330 922.510 1228.680 ;
        RECT 920.620 1220.190 922.510 1220.330 ;
        RECT 920.620 1196.530 920.760 1220.190 ;
        RECT 921.950 1219.680 922.510 1220.190 ;
        RECT 918.780 1196.390 920.760 1196.530 ;
        RECT 918.780 883.050 918.920 1196.390 ;
        RECT 918.320 882.910 918.920 883.050 ;
        RECT 918.320 881.690 918.460 882.910 ;
        RECT 918.320 881.550 918.920 881.690 ;
        RECT 918.780 787.170 918.920 881.550 ;
        RECT 918.320 787.030 918.920 787.170 ;
        RECT 918.320 786.490 918.460 787.030 ;
        RECT 918.320 786.350 918.920 786.490 ;
        RECT 918.780 690.610 918.920 786.350 ;
        RECT 918.320 690.470 918.920 690.610 ;
        RECT 918.320 688.570 918.460 690.470 ;
        RECT 918.320 688.430 918.920 688.570 ;
        RECT 918.780 594.050 918.920 688.430 ;
        RECT 918.320 593.910 918.920 594.050 ;
        RECT 918.320 593.370 918.460 593.910 ;
        RECT 918.320 593.230 918.920 593.370 ;
        RECT 918.780 303.690 918.920 593.230 ;
        RECT 918.320 303.550 918.920 303.690 ;
        RECT 918.320 303.010 918.460 303.550 ;
        RECT 918.320 302.870 918.920 303.010 ;
        RECT 918.780 110.570 918.920 302.870 ;
        RECT 918.320 110.430 918.920 110.570 ;
        RECT 918.320 109.890 918.460 110.430 ;
        RECT 918.320 109.750 918.920 109.890 ;
        RECT 918.780 34.330 918.920 109.750 ;
        RECT 335.900 34.010 336.160 34.330 ;
        RECT 918.720 34.010 918.980 34.330 ;
        RECT 335.960 2.400 336.100 34.010 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 925.130 1159.640 925.450 1159.700 ;
        RECT 929.270 1159.640 929.590 1159.700 ;
        RECT 925.130 1159.500 929.590 1159.640 ;
        RECT 925.130 1159.440 925.450 1159.500 ;
        RECT 929.270 1159.440 929.590 1159.500 ;
      LAYER via ;
        RECT 925.160 1159.440 925.420 1159.700 ;
        RECT 929.300 1159.440 929.560 1159.700 ;
      LAYER met2 ;
        RECT 931.150 1220.330 931.710 1228.680 ;
        RECT 929.360 1220.190 931.710 1220.330 ;
        RECT 929.360 1159.730 929.500 1220.190 ;
        RECT 931.150 1219.680 931.710 1220.190 ;
        RECT 925.160 1159.410 925.420 1159.730 ;
        RECT 929.300 1159.410 929.560 1159.730 ;
        RECT 925.220 37.925 925.360 1159.410 ;
        RECT 353.370 37.555 353.650 37.925 ;
        RECT 925.150 37.555 925.430 37.925 ;
        RECT 353.440 2.400 353.580 37.555 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 353.370 37.600 353.650 37.880 ;
        RECT 925.150 37.600 925.430 37.880 ;
      LAYER met3 ;
        RECT 353.345 37.890 353.675 37.905 ;
        RECT 925.125 37.890 925.455 37.905 ;
        RECT 353.345 37.590 925.455 37.890 ;
        RECT 353.345 37.575 353.675 37.590 ;
        RECT 925.125 37.575 925.455 37.590 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 371.290 45.120 371.610 45.180 ;
        RECT 938.930 45.120 939.250 45.180 ;
        RECT 371.290 44.980 939.250 45.120 ;
        RECT 371.290 44.920 371.610 44.980 ;
        RECT 938.930 44.920 939.250 44.980 ;
      LAYER via ;
        RECT 371.320 44.920 371.580 45.180 ;
        RECT 938.960 44.920 939.220 45.180 ;
      LAYER met2 ;
        RECT 940.350 1220.330 940.910 1228.680 ;
        RECT 939.020 1220.190 940.910 1220.330 ;
        RECT 939.020 45.210 939.160 1220.190 ;
        RECT 940.350 1219.680 940.910 1220.190 ;
        RECT 371.320 44.890 371.580 45.210 ;
        RECT 938.960 44.890 939.220 45.210 ;
        RECT 371.380 2.400 371.520 44.890 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 946.365 669.545 946.535 717.655 ;
        RECT 946.365 572.645 946.535 620.755 ;
        RECT 944.985 427.805 945.155 475.915 ;
        RECT 945.905 234.685 946.075 324.275 ;
        RECT 945.905 83.045 946.075 131.155 ;
      LAYER mcon ;
        RECT 946.365 717.485 946.535 717.655 ;
        RECT 946.365 620.585 946.535 620.755 ;
        RECT 944.985 475.745 945.155 475.915 ;
        RECT 945.905 324.105 946.075 324.275 ;
        RECT 945.905 130.985 946.075 131.155 ;
      LAYER met1 ;
        RECT 946.290 717.640 946.610 717.700 ;
        RECT 946.095 717.500 946.610 717.640 ;
        RECT 946.290 717.440 946.610 717.500 ;
        RECT 946.290 669.700 946.610 669.760 ;
        RECT 946.095 669.560 946.610 669.700 ;
        RECT 946.290 669.500 946.610 669.560 ;
        RECT 946.290 620.740 946.610 620.800 ;
        RECT 946.095 620.600 946.610 620.740 ;
        RECT 946.290 620.540 946.610 620.600 ;
        RECT 946.290 572.800 946.610 572.860 ;
        RECT 946.095 572.660 946.610 572.800 ;
        RECT 946.290 572.600 946.610 572.660 ;
        RECT 945.830 524.520 946.150 524.580 ;
        RECT 946.290 524.520 946.610 524.580 ;
        RECT 945.830 524.380 946.610 524.520 ;
        RECT 945.830 524.320 946.150 524.380 ;
        RECT 946.290 524.320 946.610 524.380 ;
        RECT 944.910 475.900 945.230 475.960 ;
        RECT 944.715 475.760 945.230 475.900 ;
        RECT 944.910 475.700 945.230 475.760 ;
        RECT 944.925 427.960 945.215 428.005 ;
        RECT 945.830 427.960 946.150 428.020 ;
        RECT 944.925 427.820 946.150 427.960 ;
        RECT 944.925 427.775 945.215 427.820 ;
        RECT 945.830 427.760 946.150 427.820 ;
        RECT 945.830 324.260 946.150 324.320 ;
        RECT 945.635 324.120 946.150 324.260 ;
        RECT 945.830 324.060 946.150 324.120 ;
        RECT 945.845 234.840 946.135 234.885 ;
        RECT 946.750 234.840 947.070 234.900 ;
        RECT 945.845 234.700 947.070 234.840 ;
        RECT 945.845 234.655 946.135 234.700 ;
        RECT 946.750 234.640 947.070 234.700 ;
        RECT 946.290 193.360 946.610 193.420 ;
        RECT 946.750 193.360 947.070 193.420 ;
        RECT 946.290 193.220 947.070 193.360 ;
        RECT 946.290 193.160 946.610 193.220 ;
        RECT 946.750 193.160 947.070 193.220 ;
        RECT 945.830 131.140 946.150 131.200 ;
        RECT 945.635 131.000 946.150 131.140 ;
        RECT 945.830 130.940 946.150 131.000 ;
        RECT 945.830 83.200 946.150 83.260 ;
        RECT 945.635 83.060 946.150 83.200 ;
        RECT 945.830 83.000 946.150 83.060 ;
        RECT 389.230 45.460 389.550 45.520 ;
        RECT 945.830 45.460 946.150 45.520 ;
        RECT 389.230 45.320 946.150 45.460 ;
        RECT 389.230 45.260 389.550 45.320 ;
        RECT 945.830 45.260 946.150 45.320 ;
      LAYER via ;
        RECT 946.320 717.440 946.580 717.700 ;
        RECT 946.320 669.500 946.580 669.760 ;
        RECT 946.320 620.540 946.580 620.800 ;
        RECT 946.320 572.600 946.580 572.860 ;
        RECT 945.860 524.320 946.120 524.580 ;
        RECT 946.320 524.320 946.580 524.580 ;
        RECT 944.940 475.700 945.200 475.960 ;
        RECT 945.860 427.760 946.120 428.020 ;
        RECT 945.860 324.060 946.120 324.320 ;
        RECT 946.780 234.640 947.040 234.900 ;
        RECT 946.320 193.160 946.580 193.420 ;
        RECT 946.780 193.160 947.040 193.420 ;
        RECT 945.860 130.940 946.120 131.200 ;
        RECT 945.860 83.000 946.120 83.260 ;
        RECT 389.260 45.260 389.520 45.520 ;
        RECT 945.860 45.260 946.120 45.520 ;
      LAYER met2 ;
        RECT 949.550 1220.330 950.110 1228.680 ;
        RECT 948.220 1220.190 950.110 1220.330 ;
        RECT 948.220 1196.530 948.360 1220.190 ;
        RECT 949.550 1219.680 950.110 1220.190 ;
        RECT 946.380 1196.390 948.360 1196.530 ;
        RECT 946.380 787.170 946.520 1196.390 ;
        RECT 945.920 787.030 946.520 787.170 ;
        RECT 945.920 786.490 946.060 787.030 ;
        RECT 945.920 786.350 946.520 786.490 ;
        RECT 946.380 725.405 946.520 786.350 ;
        RECT 946.310 725.035 946.590 725.405 ;
        RECT 946.310 724.355 946.590 724.725 ;
        RECT 946.380 717.730 946.520 724.355 ;
        RECT 946.320 717.410 946.580 717.730 ;
        RECT 946.320 669.470 946.580 669.790 ;
        RECT 946.380 628.845 946.520 669.470 ;
        RECT 946.310 628.475 946.590 628.845 ;
        RECT 946.310 627.795 946.590 628.165 ;
        RECT 946.380 620.830 946.520 627.795 ;
        RECT 946.320 620.510 946.580 620.830 ;
        RECT 946.320 572.570 946.580 572.890 ;
        RECT 946.380 524.610 946.520 572.570 ;
        RECT 945.860 524.290 946.120 524.610 ;
        RECT 946.320 524.290 946.580 524.610 ;
        RECT 945.920 524.125 946.060 524.290 ;
        RECT 945.850 523.755 946.130 524.125 ;
        RECT 944.930 476.155 945.210 476.525 ;
        RECT 945.000 475.990 945.140 476.155 ;
        RECT 944.940 475.670 945.200 475.990 ;
        RECT 945.860 427.730 946.120 428.050 ;
        RECT 945.920 427.565 946.060 427.730 ;
        RECT 945.850 427.195 946.130 427.565 ;
        RECT 946.310 426.515 946.590 426.885 ;
        RECT 946.380 331.060 946.520 426.515 ;
        RECT 945.920 330.920 946.520 331.060 ;
        RECT 945.920 324.350 946.060 330.920 ;
        RECT 945.860 324.030 946.120 324.350 ;
        RECT 946.780 234.610 947.040 234.930 ;
        RECT 946.840 193.450 946.980 234.610 ;
        RECT 946.320 193.130 946.580 193.450 ;
        RECT 946.780 193.130 947.040 193.450 ;
        RECT 946.380 139.245 946.520 193.130 ;
        RECT 946.310 138.875 946.590 139.245 ;
        RECT 945.850 138.195 946.130 138.565 ;
        RECT 945.920 131.230 946.060 138.195 ;
        RECT 945.860 130.910 946.120 131.230 ;
        RECT 945.860 82.970 946.120 83.290 ;
        RECT 945.920 45.550 946.060 82.970 ;
        RECT 389.260 45.230 389.520 45.550 ;
        RECT 945.860 45.230 946.120 45.550 ;
        RECT 389.320 2.400 389.460 45.230 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 946.310 725.080 946.590 725.360 ;
        RECT 946.310 724.400 946.590 724.680 ;
        RECT 946.310 628.520 946.590 628.800 ;
        RECT 946.310 627.840 946.590 628.120 ;
        RECT 945.850 523.800 946.130 524.080 ;
        RECT 944.930 476.200 945.210 476.480 ;
        RECT 945.850 427.240 946.130 427.520 ;
        RECT 946.310 426.560 946.590 426.840 ;
        RECT 946.310 138.920 946.590 139.200 ;
        RECT 945.850 138.240 946.130 138.520 ;
      LAYER met3 ;
        RECT 946.285 725.370 946.615 725.385 ;
        RECT 946.285 725.070 947.290 725.370 ;
        RECT 946.285 725.055 946.615 725.070 ;
        RECT 946.285 724.690 946.615 724.705 ;
        RECT 946.990 724.690 947.290 725.070 ;
        RECT 946.285 724.390 947.290 724.690 ;
        RECT 946.285 724.375 946.615 724.390 ;
        RECT 946.285 628.810 946.615 628.825 ;
        RECT 946.285 628.510 947.290 628.810 ;
        RECT 946.285 628.495 946.615 628.510 ;
        RECT 946.285 628.130 946.615 628.145 ;
        RECT 946.990 628.130 947.290 628.510 ;
        RECT 946.285 627.830 947.290 628.130 ;
        RECT 946.285 627.815 946.615 627.830 ;
        RECT 945.110 524.090 945.490 524.100 ;
        RECT 945.825 524.090 946.155 524.105 ;
        RECT 945.110 523.790 946.155 524.090 ;
        RECT 945.110 523.780 945.490 523.790 ;
        RECT 945.825 523.775 946.155 523.790 ;
        RECT 944.905 476.500 945.235 476.505 ;
        RECT 944.905 476.490 945.490 476.500 ;
        RECT 944.905 476.190 945.690 476.490 ;
        RECT 944.905 476.180 945.490 476.190 ;
        RECT 944.905 476.175 945.235 476.180 ;
        RECT 945.825 427.530 946.155 427.545 ;
        RECT 945.150 427.230 946.155 427.530 ;
        RECT 945.150 426.850 945.450 427.230 ;
        RECT 945.825 427.215 946.155 427.230 ;
        RECT 946.285 426.850 946.615 426.865 ;
        RECT 945.150 426.550 946.615 426.850 ;
        RECT 946.285 426.535 946.615 426.550 ;
        RECT 946.285 139.210 946.615 139.225 ;
        RECT 945.150 138.910 946.615 139.210 ;
        RECT 945.150 138.530 945.450 138.910 ;
        RECT 946.285 138.895 946.615 138.910 ;
        RECT 945.825 138.530 946.155 138.545 ;
        RECT 945.150 138.230 946.155 138.530 ;
        RECT 945.825 138.215 946.155 138.230 ;
      LAYER via3 ;
        RECT 945.140 523.780 945.460 524.100 ;
        RECT 945.140 476.180 945.460 476.500 ;
      LAYER met4 ;
        RECT 945.135 523.775 945.465 524.105 ;
        RECT 945.150 476.505 945.450 523.775 ;
        RECT 945.135 476.175 945.465 476.505 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 952.730 1196.700 953.050 1196.760 ;
        RECT 956.870 1196.700 957.190 1196.760 ;
        RECT 952.730 1196.560 957.190 1196.700 ;
        RECT 952.730 1196.500 953.050 1196.560 ;
        RECT 956.870 1196.500 957.190 1196.560 ;
        RECT 407.170 45.800 407.490 45.860 ;
        RECT 952.730 45.800 953.050 45.860 ;
        RECT 407.170 45.660 953.050 45.800 ;
        RECT 407.170 45.600 407.490 45.660 ;
        RECT 952.730 45.600 953.050 45.660 ;
      LAYER via ;
        RECT 952.760 1196.500 953.020 1196.760 ;
        RECT 956.900 1196.500 957.160 1196.760 ;
        RECT 407.200 45.600 407.460 45.860 ;
        RECT 952.760 45.600 953.020 45.860 ;
      LAYER met2 ;
        RECT 958.750 1220.330 959.310 1228.680 ;
        RECT 956.960 1220.190 959.310 1220.330 ;
        RECT 956.960 1196.790 957.100 1220.190 ;
        RECT 958.750 1219.680 959.310 1220.190 ;
        RECT 952.760 1196.470 953.020 1196.790 ;
        RECT 956.900 1196.470 957.160 1196.790 ;
        RECT 952.820 45.890 952.960 1196.470 ;
        RECT 407.200 45.570 407.460 45.890 ;
        RECT 952.760 45.570 953.020 45.890 ;
        RECT 407.260 2.400 407.400 45.570 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 780.765 1110.865 780.935 1124.975 ;
        RECT 780.765 772.905 780.935 821.015 ;
        RECT 780.765 620.925 780.935 669.375 ;
      LAYER mcon ;
        RECT 780.765 1124.805 780.935 1124.975 ;
        RECT 780.765 820.845 780.935 821.015 ;
        RECT 780.765 669.205 780.935 669.375 ;
      LAYER met1 ;
        RECT 780.690 1124.960 781.010 1125.020 ;
        RECT 780.495 1124.820 781.010 1124.960 ;
        RECT 780.690 1124.760 781.010 1124.820 ;
        RECT 780.690 1111.020 781.010 1111.080 ;
        RECT 780.495 1110.880 781.010 1111.020 ;
        RECT 780.690 1110.820 781.010 1110.880 ;
        RECT 780.690 883.020 781.010 883.280 ;
        RECT 780.780 882.600 780.920 883.020 ;
        RECT 780.690 882.340 781.010 882.600 ;
        RECT 780.690 821.000 781.010 821.060 ;
        RECT 780.495 820.860 781.010 821.000 ;
        RECT 780.690 820.800 781.010 820.860 ;
        RECT 780.690 773.060 781.010 773.120 ;
        RECT 780.495 772.920 781.010 773.060 ;
        RECT 780.690 772.860 781.010 772.920 ;
        RECT 780.690 669.360 781.010 669.420 ;
        RECT 780.495 669.220 781.010 669.360 ;
        RECT 780.690 669.160 781.010 669.220 ;
        RECT 780.690 621.080 781.010 621.140 ;
        RECT 780.495 620.940 781.010 621.080 ;
        RECT 780.690 620.880 781.010 620.940 ;
        RECT 780.690 593.680 781.010 593.940 ;
        RECT 780.780 593.260 780.920 593.680 ;
        RECT 780.690 593.000 781.010 593.260 ;
        RECT 780.690 497.120 781.010 497.380 ;
        RECT 780.780 496.700 780.920 497.120 ;
        RECT 780.690 496.440 781.010 496.700 ;
        RECT 68.150 31.520 68.470 31.580 ;
        RECT 780.690 31.520 781.010 31.580 ;
        RECT 68.150 31.380 781.010 31.520 ;
        RECT 68.150 31.320 68.470 31.380 ;
        RECT 780.690 31.320 781.010 31.380 ;
      LAYER via ;
        RECT 780.720 1124.760 780.980 1125.020 ;
        RECT 780.720 1110.820 780.980 1111.080 ;
        RECT 780.720 883.020 780.980 883.280 ;
        RECT 780.720 882.340 780.980 882.600 ;
        RECT 780.720 820.800 780.980 821.060 ;
        RECT 780.720 772.860 780.980 773.120 ;
        RECT 780.720 669.160 780.980 669.420 ;
        RECT 780.720 620.880 780.980 621.140 ;
        RECT 780.720 593.680 780.980 593.940 ;
        RECT 780.720 593.000 780.980 593.260 ;
        RECT 780.720 497.120 780.980 497.380 ;
        RECT 780.720 496.440 780.980 496.700 ;
        RECT 68.180 31.320 68.440 31.580 ;
        RECT 780.720 31.320 780.980 31.580 ;
      LAYER met2 ;
        RECT 784.870 1220.330 785.430 1228.680 ;
        RECT 782.620 1220.190 785.430 1220.330 ;
        RECT 782.620 1196.530 782.760 1220.190 ;
        RECT 784.870 1219.680 785.430 1220.190 ;
        RECT 780.780 1196.390 782.760 1196.530 ;
        RECT 780.780 1125.050 780.920 1196.390 ;
        RECT 780.720 1124.730 780.980 1125.050 ;
        RECT 780.720 1110.790 780.980 1111.110 ;
        RECT 780.780 1087.050 780.920 1110.790 ;
        RECT 780.320 1086.910 780.920 1087.050 ;
        RECT 780.320 979.610 780.460 1086.910 ;
        RECT 780.320 979.470 780.920 979.610 ;
        RECT 780.780 883.310 780.920 979.470 ;
        RECT 780.720 882.990 780.980 883.310 ;
        RECT 780.720 882.310 780.980 882.630 ;
        RECT 780.780 821.090 780.920 882.310 ;
        RECT 780.720 820.770 780.980 821.090 ;
        RECT 780.720 772.830 780.980 773.150 ;
        RECT 780.780 681.090 780.920 772.830 ;
        RECT 780.780 680.950 781.840 681.090 ;
        RECT 781.700 669.645 781.840 680.950 ;
        RECT 780.710 669.275 780.990 669.645 ;
        RECT 781.630 669.275 781.910 669.645 ;
        RECT 780.720 669.130 780.980 669.275 ;
        RECT 780.720 620.850 780.980 621.170 ;
        RECT 780.780 593.970 780.920 620.850 ;
        RECT 780.720 593.650 780.980 593.970 ;
        RECT 780.720 592.970 780.980 593.290 ;
        RECT 780.780 497.410 780.920 592.970 ;
        RECT 780.720 497.090 780.980 497.410 ;
        RECT 780.720 496.410 780.980 496.730 ;
        RECT 780.780 31.610 780.920 496.410 ;
        RECT 68.180 31.290 68.440 31.610 ;
        RECT 780.720 31.290 780.980 31.610 ;
        RECT 68.240 2.400 68.380 31.290 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 780.710 669.320 780.990 669.600 ;
        RECT 781.630 669.320 781.910 669.600 ;
      LAYER met3 ;
        RECT 780.685 669.610 781.015 669.625 ;
        RECT 781.605 669.610 781.935 669.625 ;
        RECT 780.685 669.310 781.935 669.610 ;
        RECT 780.685 669.295 781.015 669.310 ;
        RECT 781.605 669.295 781.935 669.310 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 46.140 424.970 46.200 ;
        RECT 966.530 46.140 966.850 46.200 ;
        RECT 424.650 46.000 966.850 46.140 ;
        RECT 424.650 45.940 424.970 46.000 ;
        RECT 966.530 45.940 966.850 46.000 ;
      LAYER via ;
        RECT 424.680 45.940 424.940 46.200 ;
        RECT 966.560 45.940 966.820 46.200 ;
      LAYER met2 ;
        RECT 967.950 1220.330 968.510 1228.680 ;
        RECT 966.620 1220.190 968.510 1220.330 ;
        RECT 966.620 46.230 966.760 1220.190 ;
        RECT 967.950 1219.680 968.510 1220.190 ;
        RECT 424.680 45.910 424.940 46.230 ;
        RECT 966.560 45.910 966.820 46.230 ;
        RECT 424.740 2.400 424.880 45.910 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 974.885 1131.605 975.055 1179.715 ;
        RECT 973.965 848.725 974.135 896.835 ;
        RECT 973.965 793.645 974.135 841.755 ;
        RECT 973.505 703.885 973.675 751.995 ;
        RECT 974.425 372.725 974.595 420.835 ;
        RECT 973.505 269.025 973.675 276.335 ;
        RECT 973.505 83.045 973.675 131.155 ;
      LAYER mcon ;
        RECT 974.885 1179.545 975.055 1179.715 ;
        RECT 973.965 896.665 974.135 896.835 ;
        RECT 973.965 841.585 974.135 841.755 ;
        RECT 973.505 751.825 973.675 751.995 ;
        RECT 974.425 420.665 974.595 420.835 ;
        RECT 973.505 276.165 973.675 276.335 ;
        RECT 973.505 130.985 973.675 131.155 ;
      LAYER met1 ;
        RECT 974.810 1179.700 975.130 1179.760 ;
        RECT 974.615 1179.560 975.130 1179.700 ;
        RECT 974.810 1179.500 975.130 1179.560 ;
        RECT 974.810 1131.760 975.130 1131.820 ;
        RECT 974.615 1131.620 975.130 1131.760 ;
        RECT 974.810 1131.560 975.130 1131.620 ;
        RECT 972.510 1083.140 972.830 1083.200 ;
        RECT 974.810 1083.140 975.130 1083.200 ;
        RECT 972.510 1083.000 975.130 1083.140 ;
        RECT 972.510 1082.940 972.830 1083.000 ;
        RECT 974.810 1082.940 975.130 1083.000 ;
        RECT 973.890 896.820 974.210 896.880 ;
        RECT 973.695 896.680 974.210 896.820 ;
        RECT 973.890 896.620 974.210 896.680 ;
        RECT 973.890 848.880 974.210 848.940 ;
        RECT 973.695 848.740 974.210 848.880 ;
        RECT 973.890 848.680 974.210 848.740 ;
        RECT 973.890 841.740 974.210 841.800 ;
        RECT 973.695 841.600 974.210 841.740 ;
        RECT 973.890 841.540 974.210 841.600 ;
        RECT 973.905 793.800 974.195 793.845 ;
        RECT 974.350 793.800 974.670 793.860 ;
        RECT 973.905 793.660 974.670 793.800 ;
        RECT 973.905 793.615 974.195 793.660 ;
        RECT 974.350 793.600 974.670 793.660 ;
        RECT 973.445 751.980 973.735 752.025 ;
        RECT 973.890 751.980 974.210 752.040 ;
        RECT 973.445 751.840 974.210 751.980 ;
        RECT 973.445 751.795 973.735 751.840 ;
        RECT 973.890 751.780 974.210 751.840 ;
        RECT 973.430 704.040 973.750 704.100 ;
        RECT 973.235 703.900 973.750 704.040 ;
        RECT 973.430 703.840 973.750 703.900 ;
        RECT 973.430 566.000 973.750 566.060 ;
        RECT 973.890 566.000 974.210 566.060 ;
        RECT 973.430 565.860 974.210 566.000 ;
        RECT 973.430 565.800 973.750 565.860 ;
        RECT 973.890 565.800 974.210 565.860 ;
        RECT 973.430 427.960 973.750 428.020 ;
        RECT 973.890 427.960 974.210 428.020 ;
        RECT 973.430 427.820 974.210 427.960 ;
        RECT 973.430 427.760 973.750 427.820 ;
        RECT 973.890 427.760 974.210 427.820 ;
        RECT 973.890 420.820 974.210 420.880 ;
        RECT 974.365 420.820 974.655 420.865 ;
        RECT 973.890 420.680 974.655 420.820 ;
        RECT 973.890 420.620 974.210 420.680 ;
        RECT 974.365 420.635 974.655 420.680 ;
        RECT 973.890 372.880 974.210 372.940 ;
        RECT 974.365 372.880 974.655 372.925 ;
        RECT 973.890 372.740 974.655 372.880 ;
        RECT 973.890 372.680 974.210 372.740 ;
        RECT 974.365 372.695 974.655 372.740 ;
        RECT 973.890 352.480 974.210 352.540 ;
        RECT 973.520 352.340 974.210 352.480 ;
        RECT 973.520 351.860 973.660 352.340 ;
        RECT 973.890 352.280 974.210 352.340 ;
        RECT 973.430 351.600 973.750 351.860 ;
        RECT 973.430 276.320 973.750 276.380 ;
        RECT 973.235 276.180 973.750 276.320 ;
        RECT 973.430 276.120 973.750 276.180 ;
        RECT 973.430 269.180 973.750 269.240 ;
        RECT 973.235 269.040 973.750 269.180 ;
        RECT 973.430 268.980 973.750 269.040 ;
        RECT 973.430 229.060 973.750 229.120 ;
        RECT 973.430 228.920 974.120 229.060 ;
        RECT 973.430 228.860 973.750 228.920 ;
        RECT 973.980 228.100 974.120 228.920 ;
        RECT 973.890 227.840 974.210 228.100 ;
        RECT 972.510 172.620 972.830 172.680 ;
        RECT 973.430 172.620 973.750 172.680 ;
        RECT 972.510 172.480 973.750 172.620 ;
        RECT 972.510 172.420 972.830 172.480 ;
        RECT 973.430 172.420 973.750 172.480 ;
        RECT 973.430 131.140 973.750 131.200 ;
        RECT 973.235 131.000 973.750 131.140 ;
        RECT 973.430 130.940 973.750 131.000 ;
        RECT 973.430 83.200 973.750 83.260 ;
        RECT 973.235 83.060 973.750 83.200 ;
        RECT 973.430 83.000 973.750 83.060 ;
        RECT 442.590 46.480 442.910 46.540 ;
        RECT 973.890 46.480 974.210 46.540 ;
        RECT 442.590 46.340 974.210 46.480 ;
        RECT 442.590 46.280 442.910 46.340 ;
        RECT 973.890 46.280 974.210 46.340 ;
      LAYER via ;
        RECT 974.840 1179.500 975.100 1179.760 ;
        RECT 974.840 1131.560 975.100 1131.820 ;
        RECT 972.540 1082.940 972.800 1083.200 ;
        RECT 974.840 1082.940 975.100 1083.200 ;
        RECT 973.920 896.620 974.180 896.880 ;
        RECT 973.920 848.680 974.180 848.940 ;
        RECT 973.920 841.540 974.180 841.800 ;
        RECT 974.380 793.600 974.640 793.860 ;
        RECT 973.920 751.780 974.180 752.040 ;
        RECT 973.460 703.840 973.720 704.100 ;
        RECT 973.460 565.800 973.720 566.060 ;
        RECT 973.920 565.800 974.180 566.060 ;
        RECT 973.460 427.760 973.720 428.020 ;
        RECT 973.920 427.760 974.180 428.020 ;
        RECT 973.920 420.620 974.180 420.880 ;
        RECT 973.920 372.680 974.180 372.940 ;
        RECT 973.920 352.280 974.180 352.540 ;
        RECT 973.460 351.600 973.720 351.860 ;
        RECT 973.460 276.120 973.720 276.380 ;
        RECT 973.460 268.980 973.720 269.240 ;
        RECT 973.460 228.860 973.720 229.120 ;
        RECT 973.920 227.840 974.180 228.100 ;
        RECT 972.540 172.420 972.800 172.680 ;
        RECT 973.460 172.420 973.720 172.680 ;
        RECT 973.460 130.940 973.720 131.200 ;
        RECT 973.460 83.000 973.720 83.260 ;
        RECT 442.620 46.280 442.880 46.540 ;
        RECT 973.920 46.280 974.180 46.540 ;
      LAYER met2 ;
        RECT 977.150 1221.010 977.710 1228.680 ;
        RECT 974.900 1220.870 977.710 1221.010 ;
        RECT 974.900 1179.790 975.040 1220.870 ;
        RECT 977.150 1219.680 977.710 1220.870 ;
        RECT 974.840 1179.470 975.100 1179.790 ;
        RECT 974.840 1131.530 975.100 1131.850 ;
        RECT 974.900 1083.230 975.040 1131.530 ;
        RECT 972.540 1082.910 972.800 1083.230 ;
        RECT 974.840 1082.910 975.100 1083.230 ;
        RECT 972.600 994.005 972.740 1082.910 ;
        RECT 972.530 993.635 972.810 994.005 ;
        RECT 973.910 992.275 974.190 992.645 ;
        RECT 973.980 896.910 974.120 992.275 ;
        RECT 973.920 896.590 974.180 896.910 ;
        RECT 973.920 848.650 974.180 848.970 ;
        RECT 973.980 841.830 974.120 848.650 ;
        RECT 973.920 841.510 974.180 841.830 ;
        RECT 974.380 793.570 974.640 793.890 ;
        RECT 974.440 785.810 974.580 793.570 ;
        RECT 973.980 785.670 974.580 785.810 ;
        RECT 973.980 752.070 974.120 785.670 ;
        RECT 973.920 751.750 974.180 752.070 ;
        RECT 973.460 703.810 973.720 704.130 ;
        RECT 973.520 566.090 973.660 703.810 ;
        RECT 973.460 565.770 973.720 566.090 ;
        RECT 973.920 565.770 974.180 566.090 ;
        RECT 973.980 545.770 974.120 565.770 ;
        RECT 973.980 545.630 974.580 545.770 ;
        RECT 974.440 542.370 974.580 545.630 ;
        RECT 973.980 542.230 974.580 542.370 ;
        RECT 973.980 428.050 974.120 542.230 ;
        RECT 973.460 427.730 973.720 428.050 ;
        RECT 973.920 427.730 974.180 428.050 ;
        RECT 973.520 427.450 973.660 427.730 ;
        RECT 973.520 427.310 974.120 427.450 ;
        RECT 973.980 420.910 974.120 427.310 ;
        RECT 973.920 420.590 974.180 420.910 ;
        RECT 973.920 372.650 974.180 372.970 ;
        RECT 973.980 352.570 974.120 372.650 ;
        RECT 973.920 352.250 974.180 352.570 ;
        RECT 973.460 351.570 973.720 351.890 ;
        RECT 973.520 276.410 973.660 351.570 ;
        RECT 973.460 276.090 973.720 276.410 ;
        RECT 973.460 268.950 973.720 269.270 ;
        RECT 973.520 229.150 973.660 268.950 ;
        RECT 973.460 228.830 973.720 229.150 ;
        RECT 973.920 227.810 974.180 228.130 ;
        RECT 973.980 220.845 974.120 227.810 ;
        RECT 972.530 220.475 972.810 220.845 ;
        RECT 973.910 220.475 974.190 220.845 ;
        RECT 972.600 172.710 972.740 220.475 ;
        RECT 972.540 172.390 972.800 172.710 ;
        RECT 973.460 172.390 973.720 172.710 ;
        RECT 973.520 131.230 973.660 172.390 ;
        RECT 973.460 130.910 973.720 131.230 ;
        RECT 973.460 82.970 973.720 83.290 ;
        RECT 973.520 48.010 973.660 82.970 ;
        RECT 973.520 47.870 974.120 48.010 ;
        RECT 973.980 46.570 974.120 47.870 ;
        RECT 442.620 46.250 442.880 46.570 ;
        RECT 973.920 46.250 974.180 46.570 ;
        RECT 442.680 2.400 442.820 46.250 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 972.530 993.680 972.810 993.960 ;
        RECT 973.910 992.320 974.190 992.600 ;
        RECT 972.530 220.520 972.810 220.800 ;
        RECT 973.910 220.520 974.190 220.800 ;
      LAYER met3 ;
        RECT 972.505 993.970 972.835 993.985 ;
        RECT 972.505 993.655 973.050 993.970 ;
        RECT 972.750 992.610 973.050 993.655 ;
        RECT 973.885 992.610 974.215 992.625 ;
        RECT 972.750 992.310 974.215 992.610 ;
        RECT 973.885 992.295 974.215 992.310 ;
        RECT 972.505 220.810 972.835 220.825 ;
        RECT 973.885 220.810 974.215 220.825 ;
        RECT 972.505 220.510 974.215 220.810 ;
        RECT 972.505 220.495 972.835 220.510 ;
        RECT 973.885 220.495 974.215 220.510 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 980.330 1196.700 980.650 1196.760 ;
        RECT 984.470 1196.700 984.790 1196.760 ;
        RECT 980.330 1196.560 984.790 1196.700 ;
        RECT 980.330 1196.500 980.650 1196.560 ;
        RECT 984.470 1196.500 984.790 1196.560 ;
        RECT 460.530 46.820 460.850 46.880 ;
        RECT 980.330 46.820 980.650 46.880 ;
        RECT 460.530 46.680 980.650 46.820 ;
        RECT 460.530 46.620 460.850 46.680 ;
        RECT 980.330 46.620 980.650 46.680 ;
      LAYER via ;
        RECT 980.360 1196.500 980.620 1196.760 ;
        RECT 984.500 1196.500 984.760 1196.760 ;
        RECT 460.560 46.620 460.820 46.880 ;
        RECT 980.360 46.620 980.620 46.880 ;
      LAYER met2 ;
        RECT 986.350 1220.330 986.910 1228.680 ;
        RECT 984.560 1220.190 986.910 1220.330 ;
        RECT 984.560 1196.790 984.700 1220.190 ;
        RECT 986.350 1219.680 986.910 1220.190 ;
        RECT 980.360 1196.470 980.620 1196.790 ;
        RECT 984.500 1196.470 984.760 1196.790 ;
        RECT 980.420 46.910 980.560 1196.470 ;
        RECT 460.560 46.590 460.820 46.910 ;
        RECT 980.360 46.590 980.620 46.910 ;
        RECT 460.620 2.400 460.760 46.590 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 478.470 47.160 478.790 47.220 ;
        RECT 994.130 47.160 994.450 47.220 ;
        RECT 478.470 47.020 994.450 47.160 ;
        RECT 478.470 46.960 478.790 47.020 ;
        RECT 994.130 46.960 994.450 47.020 ;
      LAYER via ;
        RECT 478.500 46.960 478.760 47.220 ;
        RECT 994.160 46.960 994.420 47.220 ;
      LAYER met2 ;
        RECT 995.550 1220.330 996.110 1228.680 ;
        RECT 994.220 1220.190 996.110 1220.330 ;
        RECT 994.220 47.250 994.360 1220.190 ;
        RECT 995.550 1219.680 996.110 1220.190 ;
        RECT 478.500 46.930 478.760 47.250 ;
        RECT 994.160 46.930 994.420 47.250 ;
        RECT 478.560 2.400 478.700 46.930 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 817.490 1211.320 817.810 1211.380 ;
        RECT 1004.710 1211.320 1005.030 1211.380 ;
        RECT 817.490 1211.180 1005.030 1211.320 ;
        RECT 817.490 1211.120 817.810 1211.180 ;
        RECT 1004.710 1211.120 1005.030 1211.180 ;
        RECT 496.410 28.120 496.730 28.180 ;
        RECT 817.490 28.120 817.810 28.180 ;
        RECT 496.410 27.980 817.810 28.120 ;
        RECT 496.410 27.920 496.730 27.980 ;
        RECT 817.490 27.920 817.810 27.980 ;
      LAYER via ;
        RECT 817.520 1211.120 817.780 1211.380 ;
        RECT 1004.740 1211.120 1005.000 1211.380 ;
        RECT 496.440 27.920 496.700 28.180 ;
        RECT 817.520 27.920 817.780 28.180 ;
      LAYER met2 ;
        RECT 1004.750 1219.680 1005.310 1228.680 ;
        RECT 1004.800 1211.410 1004.940 1219.680 ;
        RECT 817.520 1211.090 817.780 1211.410 ;
        RECT 1004.740 1211.090 1005.000 1211.410 ;
        RECT 817.580 28.210 817.720 1211.090 ;
        RECT 496.440 27.890 496.700 28.210 ;
        RECT 817.520 27.890 817.780 28.210 ;
        RECT 496.500 2.400 496.640 27.890 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.930 1196.700 1008.250 1196.760 ;
        RECT 1012.070 1196.700 1012.390 1196.760 ;
        RECT 1007.930 1196.560 1012.390 1196.700 ;
        RECT 1007.930 1196.500 1008.250 1196.560 ;
        RECT 1012.070 1196.500 1012.390 1196.560 ;
        RECT 513.890 47.500 514.210 47.560 ;
        RECT 1007.930 47.500 1008.250 47.560 ;
        RECT 513.890 47.360 1008.250 47.500 ;
        RECT 513.890 47.300 514.210 47.360 ;
        RECT 1007.930 47.300 1008.250 47.360 ;
      LAYER via ;
        RECT 1007.960 1196.500 1008.220 1196.760 ;
        RECT 1012.100 1196.500 1012.360 1196.760 ;
        RECT 513.920 47.300 514.180 47.560 ;
        RECT 1007.960 47.300 1008.220 47.560 ;
      LAYER met2 ;
        RECT 1013.950 1220.330 1014.510 1228.680 ;
        RECT 1012.160 1220.190 1014.510 1220.330 ;
        RECT 1012.160 1196.790 1012.300 1220.190 ;
        RECT 1013.950 1219.680 1014.510 1220.190 ;
        RECT 1007.960 1196.470 1008.220 1196.790 ;
        RECT 1012.100 1196.470 1012.360 1196.790 ;
        RECT 1008.020 47.590 1008.160 1196.470 ;
        RECT 513.920 47.270 514.180 47.590 ;
        RECT 1007.960 47.270 1008.220 47.590 ;
        RECT 513.980 2.400 514.120 47.270 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.830 47.840 532.150 47.900 ;
        RECT 1021.730 47.840 1022.050 47.900 ;
        RECT 531.830 47.700 1022.050 47.840 ;
        RECT 531.830 47.640 532.150 47.700 ;
        RECT 1021.730 47.640 1022.050 47.700 ;
      LAYER via ;
        RECT 531.860 47.640 532.120 47.900 ;
        RECT 1021.760 47.640 1022.020 47.900 ;
      LAYER met2 ;
        RECT 1023.150 1220.330 1023.710 1228.680 ;
        RECT 1021.820 1220.190 1023.710 1220.330 ;
        RECT 1021.820 47.930 1021.960 1220.190 ;
        RECT 1023.150 1219.680 1023.710 1220.190 ;
        RECT 531.860 47.610 532.120 47.930 ;
        RECT 1021.760 47.610 1022.020 47.930 ;
        RECT 531.920 2.400 532.060 47.610 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1030.085 786.505 1030.255 814.215 ;
        RECT 1030.085 469.285 1030.255 517.395 ;
        RECT 1030.085 427.805 1030.255 435.115 ;
      LAYER mcon ;
        RECT 1030.085 814.045 1030.255 814.215 ;
        RECT 1030.085 517.225 1030.255 517.395 ;
        RECT 1030.085 434.945 1030.255 435.115 ;
      LAYER met1 ;
        RECT 1029.090 1111.020 1029.410 1111.080 ;
        RECT 1029.550 1111.020 1029.870 1111.080 ;
        RECT 1029.090 1110.880 1029.870 1111.020 ;
        RECT 1029.090 1110.820 1029.410 1110.880 ;
        RECT 1029.550 1110.820 1029.870 1110.880 ;
        RECT 1029.550 1031.460 1029.870 1031.520 ;
        RECT 1030.470 1031.460 1030.790 1031.520 ;
        RECT 1029.550 1031.320 1030.790 1031.460 ;
        RECT 1029.550 1031.260 1029.870 1031.320 ;
        RECT 1030.470 1031.260 1030.790 1031.320 ;
        RECT 1029.550 1007.120 1029.870 1007.380 ;
        RECT 1029.640 1006.980 1029.780 1007.120 ;
        RECT 1030.010 1006.980 1030.330 1007.040 ;
        RECT 1029.640 1006.840 1030.330 1006.980 ;
        RECT 1030.010 1006.780 1030.330 1006.840 ;
        RECT 1029.550 869.620 1029.870 869.680 ;
        RECT 1030.470 869.620 1030.790 869.680 ;
        RECT 1029.550 869.480 1030.790 869.620 ;
        RECT 1029.550 869.420 1029.870 869.480 ;
        RECT 1030.470 869.420 1030.790 869.480 ;
        RECT 1030.010 814.200 1030.330 814.260 ;
        RECT 1029.815 814.060 1030.330 814.200 ;
        RECT 1030.010 814.000 1030.330 814.060 ;
        RECT 1030.010 786.660 1030.330 786.720 ;
        RECT 1029.815 786.520 1030.330 786.660 ;
        RECT 1030.010 786.460 1030.330 786.520 ;
        RECT 1029.550 724.440 1029.870 724.500 ;
        RECT 1030.010 724.440 1030.330 724.500 ;
        RECT 1029.550 724.300 1030.330 724.440 ;
        RECT 1029.550 724.240 1029.870 724.300 ;
        RECT 1030.010 724.240 1030.330 724.300 ;
        RECT 1029.550 717.640 1029.870 717.700 ;
        RECT 1030.470 717.640 1030.790 717.700 ;
        RECT 1029.550 717.500 1030.790 717.640 ;
        RECT 1029.550 717.440 1029.870 717.500 ;
        RECT 1030.470 717.440 1030.790 717.500 ;
        RECT 1029.090 627.880 1029.410 627.940 ;
        RECT 1030.010 627.880 1030.330 627.940 ;
        RECT 1029.090 627.740 1030.330 627.880 ;
        RECT 1029.090 627.680 1029.410 627.740 ;
        RECT 1030.010 627.680 1030.330 627.740 ;
        RECT 1029.090 524.520 1029.410 524.580 ;
        RECT 1030.010 524.520 1030.330 524.580 ;
        RECT 1029.090 524.380 1030.330 524.520 ;
        RECT 1029.090 524.320 1029.410 524.380 ;
        RECT 1030.010 524.320 1030.330 524.380 ;
        RECT 1030.010 517.380 1030.330 517.440 ;
        RECT 1029.815 517.240 1030.330 517.380 ;
        RECT 1030.010 517.180 1030.330 517.240 ;
        RECT 1030.010 469.440 1030.330 469.500 ;
        RECT 1029.815 469.300 1030.330 469.440 ;
        RECT 1030.010 469.240 1030.330 469.300 ;
        RECT 1030.010 435.100 1030.330 435.160 ;
        RECT 1029.815 434.960 1030.330 435.100 ;
        RECT 1030.010 434.900 1030.330 434.960 ;
        RECT 1030.010 427.960 1030.330 428.020 ;
        RECT 1029.815 427.820 1030.330 427.960 ;
        RECT 1030.010 427.760 1030.330 427.820 ;
        RECT 1028.630 145.080 1028.950 145.140 ;
        RECT 1029.090 145.080 1029.410 145.140 ;
        RECT 1028.630 144.940 1029.410 145.080 ;
        RECT 1028.630 144.880 1028.950 144.940 ;
        RECT 1029.090 144.880 1029.410 144.940 ;
        RECT 1029.090 137.940 1029.410 138.000 ;
        RECT 1029.550 137.940 1029.870 138.000 ;
        RECT 1029.090 137.800 1029.870 137.940 ;
        RECT 1029.090 137.740 1029.410 137.800 ;
        RECT 1029.550 137.740 1029.870 137.800 ;
        RECT 549.770 48.180 550.090 48.240 ;
        RECT 1029.090 48.180 1029.410 48.240 ;
        RECT 549.770 48.040 1029.410 48.180 ;
        RECT 549.770 47.980 550.090 48.040 ;
        RECT 1029.090 47.980 1029.410 48.040 ;
      LAYER via ;
        RECT 1029.120 1110.820 1029.380 1111.080 ;
        RECT 1029.580 1110.820 1029.840 1111.080 ;
        RECT 1029.580 1031.260 1029.840 1031.520 ;
        RECT 1030.500 1031.260 1030.760 1031.520 ;
        RECT 1029.580 1007.120 1029.840 1007.380 ;
        RECT 1030.040 1006.780 1030.300 1007.040 ;
        RECT 1029.580 869.420 1029.840 869.680 ;
        RECT 1030.500 869.420 1030.760 869.680 ;
        RECT 1030.040 814.000 1030.300 814.260 ;
        RECT 1030.040 786.460 1030.300 786.720 ;
        RECT 1029.580 724.240 1029.840 724.500 ;
        RECT 1030.040 724.240 1030.300 724.500 ;
        RECT 1029.580 717.440 1029.840 717.700 ;
        RECT 1030.500 717.440 1030.760 717.700 ;
        RECT 1029.120 627.680 1029.380 627.940 ;
        RECT 1030.040 627.680 1030.300 627.940 ;
        RECT 1029.120 524.320 1029.380 524.580 ;
        RECT 1030.040 524.320 1030.300 524.580 ;
        RECT 1030.040 517.180 1030.300 517.440 ;
        RECT 1030.040 469.240 1030.300 469.500 ;
        RECT 1030.040 434.900 1030.300 435.160 ;
        RECT 1030.040 427.760 1030.300 428.020 ;
        RECT 1028.660 144.880 1028.920 145.140 ;
        RECT 1029.120 144.880 1029.380 145.140 ;
        RECT 1029.120 137.740 1029.380 138.000 ;
        RECT 1029.580 137.740 1029.840 138.000 ;
        RECT 549.800 47.980 550.060 48.240 ;
        RECT 1029.120 47.980 1029.380 48.240 ;
      LAYER met2 ;
        RECT 1032.350 1221.010 1032.910 1228.680 ;
        RECT 1030.100 1220.870 1032.910 1221.010 ;
        RECT 1030.100 1196.530 1030.240 1220.870 ;
        RECT 1032.350 1219.680 1032.910 1220.870 ;
        RECT 1029.640 1196.390 1030.240 1196.530 ;
        RECT 1029.640 1111.110 1029.780 1196.390 ;
        RECT 1029.120 1110.790 1029.380 1111.110 ;
        RECT 1029.580 1110.790 1029.840 1111.110 ;
        RECT 1029.180 1097.250 1029.320 1110.790 ;
        RECT 1029.180 1097.110 1029.780 1097.250 ;
        RECT 1029.640 1031.550 1029.780 1097.110 ;
        RECT 1029.580 1031.230 1029.840 1031.550 ;
        RECT 1030.500 1031.230 1030.760 1031.550 ;
        RECT 1030.560 1007.605 1030.700 1031.230 ;
        RECT 1029.570 1007.235 1029.850 1007.605 ;
        RECT 1030.490 1007.235 1030.770 1007.605 ;
        RECT 1029.580 1007.090 1029.840 1007.235 ;
        RECT 1030.040 1006.750 1030.300 1007.070 ;
        RECT 1030.100 893.930 1030.240 1006.750 ;
        RECT 1030.100 893.790 1030.700 893.930 ;
        RECT 1030.560 869.710 1030.700 893.790 ;
        RECT 1029.580 869.390 1029.840 869.710 ;
        RECT 1030.500 869.390 1030.760 869.710 ;
        RECT 1029.640 847.010 1029.780 869.390 ;
        RECT 1029.640 846.870 1030.240 847.010 ;
        RECT 1030.100 814.290 1030.240 846.870 ;
        RECT 1030.040 813.970 1030.300 814.290 ;
        RECT 1030.040 786.430 1030.300 786.750 ;
        RECT 1030.100 724.530 1030.240 786.430 ;
        RECT 1029.580 724.210 1029.840 724.530 ;
        RECT 1030.040 724.210 1030.300 724.530 ;
        RECT 1029.640 717.730 1029.780 724.210 ;
        RECT 1029.580 717.410 1029.840 717.730 ;
        RECT 1030.500 717.410 1030.760 717.730 ;
        RECT 1030.560 641.650 1030.700 717.410 ;
        RECT 1030.100 641.510 1030.700 641.650 ;
        RECT 1030.100 627.970 1030.240 641.510 ;
        RECT 1029.120 627.650 1029.380 627.970 ;
        RECT 1030.040 627.650 1030.300 627.970 ;
        RECT 1029.180 593.370 1029.320 627.650 ;
        RECT 1029.180 593.230 1029.780 593.370 ;
        RECT 1029.640 548.490 1029.780 593.230 ;
        RECT 1029.180 548.350 1029.780 548.490 ;
        RECT 1029.180 524.610 1029.320 548.350 ;
        RECT 1029.120 524.290 1029.380 524.610 ;
        RECT 1030.040 524.290 1030.300 524.610 ;
        RECT 1030.100 517.470 1030.240 524.290 ;
        RECT 1030.040 517.150 1030.300 517.470 ;
        RECT 1030.040 469.210 1030.300 469.530 ;
        RECT 1030.100 435.190 1030.240 469.210 ;
        RECT 1030.040 434.870 1030.300 435.190 ;
        RECT 1030.040 427.730 1030.300 428.050 ;
        RECT 1030.100 410.450 1030.240 427.730 ;
        RECT 1029.640 410.310 1030.240 410.450 ;
        RECT 1029.640 255.410 1029.780 410.310 ;
        RECT 1029.180 255.270 1029.780 255.410 ;
        RECT 1029.180 207.130 1029.320 255.270 ;
        RECT 1028.720 206.990 1029.320 207.130 ;
        RECT 1028.720 145.170 1028.860 206.990 ;
        RECT 1028.660 144.850 1028.920 145.170 ;
        RECT 1029.120 144.850 1029.380 145.170 ;
        RECT 1029.180 138.030 1029.320 144.850 ;
        RECT 1029.120 137.710 1029.380 138.030 ;
        RECT 1029.580 137.710 1029.840 138.030 ;
        RECT 1029.640 61.610 1029.780 137.710 ;
        RECT 1029.180 61.470 1029.780 61.610 ;
        RECT 1029.180 48.270 1029.320 61.470 ;
        RECT 549.800 47.950 550.060 48.270 ;
        RECT 1029.120 47.950 1029.380 48.270 ;
        RECT 549.860 2.400 550.000 47.950 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 1029.570 1007.280 1029.850 1007.560 ;
        RECT 1030.490 1007.280 1030.770 1007.560 ;
      LAYER met3 ;
        RECT 1029.545 1007.570 1029.875 1007.585 ;
        RECT 1030.465 1007.570 1030.795 1007.585 ;
        RECT 1029.545 1007.270 1030.795 1007.570 ;
        RECT 1029.545 1007.255 1029.875 1007.270 ;
        RECT 1030.465 1007.255 1030.795 1007.270 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 804.150 1207.580 804.470 1207.640 ;
        RECT 1041.050 1207.580 1041.370 1207.640 ;
        RECT 804.150 1207.440 1041.370 1207.580 ;
        RECT 804.150 1207.380 804.470 1207.440 ;
        RECT 1041.050 1207.380 1041.370 1207.440 ;
        RECT 567.710 27.780 568.030 27.840 ;
        RECT 803.690 27.780 804.010 27.840 ;
        RECT 567.710 27.640 804.010 27.780 ;
        RECT 567.710 27.580 568.030 27.640 ;
        RECT 803.690 27.580 804.010 27.640 ;
      LAYER via ;
        RECT 804.180 1207.380 804.440 1207.640 ;
        RECT 1041.080 1207.380 1041.340 1207.640 ;
        RECT 567.740 27.580 568.000 27.840 ;
        RECT 803.720 27.580 803.980 27.840 ;
      LAYER met2 ;
        RECT 1041.090 1219.680 1041.650 1228.680 ;
        RECT 1041.140 1207.670 1041.280 1219.680 ;
        RECT 804.180 1207.350 804.440 1207.670 ;
        RECT 1041.080 1207.350 1041.340 1207.670 ;
        RECT 804.240 1182.930 804.380 1207.350 ;
        RECT 803.780 1182.790 804.380 1182.930 ;
        RECT 803.780 27.870 803.920 1182.790 ;
        RECT 567.740 27.550 568.000 27.870 ;
        RECT 803.720 27.550 803.980 27.870 ;
        RECT 567.800 2.400 567.940 27.550 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 44.440 585.970 44.500 ;
        RECT 1049.330 44.440 1049.650 44.500 ;
        RECT 585.650 44.300 1049.650 44.440 ;
        RECT 585.650 44.240 585.970 44.300 ;
        RECT 1049.330 44.240 1049.650 44.300 ;
      LAYER via ;
        RECT 585.680 44.240 585.940 44.500 ;
        RECT 1049.360 44.240 1049.620 44.500 ;
      LAYER met2 ;
        RECT 1050.290 1220.330 1050.850 1228.680 ;
        RECT 1049.420 1220.190 1050.850 1220.330 ;
        RECT 1049.420 44.530 1049.560 1220.190 ;
        RECT 1050.290 1219.680 1050.850 1220.190 ;
        RECT 585.680 44.210 585.940 44.530 ;
        RECT 1049.360 44.210 1049.620 44.530 ;
        RECT 585.740 2.400 585.880 44.210 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 31.860 91.930 31.920 ;
        RECT 794.490 31.860 794.810 31.920 ;
        RECT 91.610 31.720 794.810 31.860 ;
        RECT 91.610 31.660 91.930 31.720 ;
        RECT 794.490 31.660 794.810 31.720 ;
      LAYER via ;
        RECT 91.640 31.660 91.900 31.920 ;
        RECT 794.520 31.660 794.780 31.920 ;
      LAYER met2 ;
        RECT 796.830 1220.330 797.390 1228.680 ;
        RECT 794.580 1220.190 797.390 1220.330 ;
        RECT 794.580 31.950 794.720 1220.190 ;
        RECT 796.830 1219.680 797.390 1220.190 ;
        RECT 91.640 31.630 91.900 31.950 ;
        RECT 794.520 31.630 794.780 31.950 ;
        RECT 91.700 2.400 91.840 31.630 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1056.765 427.805 1056.935 475.915 ;
        RECT 1056.305 324.785 1056.475 372.555 ;
        RECT 1056.765 276.165 1056.935 324.275 ;
        RECT 1056.305 227.885 1056.475 236.555 ;
        RECT 1056.765 96.645 1056.935 137.955 ;
      LAYER mcon ;
        RECT 1056.765 475.745 1056.935 475.915 ;
        RECT 1056.305 372.385 1056.475 372.555 ;
        RECT 1056.765 324.105 1056.935 324.275 ;
        RECT 1056.305 236.385 1056.475 236.555 ;
        RECT 1056.765 137.785 1056.935 137.955 ;
      LAYER met1 ;
        RECT 1056.230 1159.300 1056.550 1159.360 ;
        RECT 1057.610 1159.300 1057.930 1159.360 ;
        RECT 1056.230 1159.160 1057.930 1159.300 ;
        RECT 1056.230 1159.100 1056.550 1159.160 ;
        RECT 1057.610 1159.100 1057.930 1159.160 ;
        RECT 1056.230 1014.460 1056.550 1014.520 ;
        RECT 1056.690 1014.460 1057.010 1014.520 ;
        RECT 1056.230 1014.320 1057.010 1014.460 ;
        RECT 1056.230 1014.260 1056.550 1014.320 ;
        RECT 1056.690 1014.260 1057.010 1014.320 ;
        RECT 1056.230 869.620 1056.550 869.680 ;
        RECT 1056.690 869.620 1057.010 869.680 ;
        RECT 1056.230 869.480 1057.010 869.620 ;
        RECT 1056.230 869.420 1056.550 869.480 ;
        RECT 1056.690 869.420 1057.010 869.480 ;
        RECT 1056.230 786.800 1056.550 787.060 ;
        RECT 1056.320 786.380 1056.460 786.800 ;
        RECT 1056.230 786.120 1056.550 786.380 ;
        RECT 1056.230 724.440 1056.550 724.500 ;
        RECT 1057.150 724.440 1057.470 724.500 ;
        RECT 1056.230 724.300 1057.470 724.440 ;
        RECT 1056.230 724.240 1056.550 724.300 ;
        RECT 1057.150 724.240 1057.470 724.300 ;
        RECT 1056.230 627.680 1056.550 627.940 ;
        RECT 1056.320 627.540 1056.460 627.680 ;
        RECT 1056.690 627.540 1057.010 627.600 ;
        RECT 1056.320 627.400 1057.010 627.540 ;
        RECT 1056.690 627.340 1057.010 627.400 ;
        RECT 1056.690 531.460 1057.010 531.720 ;
        RECT 1056.780 530.700 1056.920 531.460 ;
        RECT 1056.690 530.440 1057.010 530.700 ;
        RECT 1056.690 475.900 1057.010 475.960 ;
        RECT 1056.495 475.760 1057.010 475.900 ;
        RECT 1056.690 475.700 1057.010 475.760 ;
        RECT 1056.690 427.960 1057.010 428.020 ;
        RECT 1056.495 427.820 1057.010 427.960 ;
        RECT 1056.690 427.760 1057.010 427.820 ;
        RECT 1056.230 372.540 1056.550 372.600 ;
        RECT 1056.035 372.400 1056.550 372.540 ;
        RECT 1056.230 372.340 1056.550 372.400 ;
        RECT 1056.245 324.940 1056.535 324.985 ;
        RECT 1056.690 324.940 1057.010 325.000 ;
        RECT 1056.245 324.800 1057.010 324.940 ;
        RECT 1056.245 324.755 1056.535 324.800 ;
        RECT 1056.690 324.740 1057.010 324.800 ;
        RECT 1056.690 324.260 1057.010 324.320 ;
        RECT 1056.495 324.120 1057.010 324.260 ;
        RECT 1056.690 324.060 1057.010 324.120 ;
        RECT 1056.705 276.320 1056.995 276.365 ;
        RECT 1057.610 276.320 1057.930 276.380 ;
        RECT 1056.705 276.180 1057.930 276.320 ;
        RECT 1056.705 276.135 1056.995 276.180 ;
        RECT 1057.610 276.120 1057.930 276.180 ;
        RECT 1056.245 236.540 1056.535 236.585 ;
        RECT 1057.610 236.540 1057.930 236.600 ;
        RECT 1056.245 236.400 1057.930 236.540 ;
        RECT 1056.245 236.355 1056.535 236.400 ;
        RECT 1057.610 236.340 1057.930 236.400 ;
        RECT 1056.230 228.040 1056.550 228.100 ;
        RECT 1056.035 227.900 1056.550 228.040 ;
        RECT 1056.230 227.840 1056.550 227.900 ;
        RECT 1056.230 137.940 1056.550 138.000 ;
        RECT 1056.705 137.940 1056.995 137.985 ;
        RECT 1056.230 137.800 1056.995 137.940 ;
        RECT 1056.230 137.740 1056.550 137.800 ;
        RECT 1056.705 137.755 1056.995 137.800 ;
        RECT 1056.690 96.800 1057.010 96.860 ;
        RECT 1056.495 96.660 1057.010 96.800 ;
        RECT 1056.690 96.600 1057.010 96.660 ;
        RECT 603.130 44.100 603.450 44.160 ;
        RECT 1056.690 44.100 1057.010 44.160 ;
        RECT 603.130 43.960 1057.010 44.100 ;
        RECT 603.130 43.900 603.450 43.960 ;
        RECT 1056.690 43.900 1057.010 43.960 ;
      LAYER via ;
        RECT 1056.260 1159.100 1056.520 1159.360 ;
        RECT 1057.640 1159.100 1057.900 1159.360 ;
        RECT 1056.260 1014.260 1056.520 1014.520 ;
        RECT 1056.720 1014.260 1056.980 1014.520 ;
        RECT 1056.260 869.420 1056.520 869.680 ;
        RECT 1056.720 869.420 1056.980 869.680 ;
        RECT 1056.260 786.800 1056.520 787.060 ;
        RECT 1056.260 786.120 1056.520 786.380 ;
        RECT 1056.260 724.240 1056.520 724.500 ;
        RECT 1057.180 724.240 1057.440 724.500 ;
        RECT 1056.260 627.680 1056.520 627.940 ;
        RECT 1056.720 627.340 1056.980 627.600 ;
        RECT 1056.720 531.460 1056.980 531.720 ;
        RECT 1056.720 530.440 1056.980 530.700 ;
        RECT 1056.720 475.700 1056.980 475.960 ;
        RECT 1056.720 427.760 1056.980 428.020 ;
        RECT 1056.260 372.340 1056.520 372.600 ;
        RECT 1056.720 324.740 1056.980 325.000 ;
        RECT 1056.720 324.060 1056.980 324.320 ;
        RECT 1057.640 276.120 1057.900 276.380 ;
        RECT 1057.640 236.340 1057.900 236.600 ;
        RECT 1056.260 227.840 1056.520 228.100 ;
        RECT 1056.260 137.740 1056.520 138.000 ;
        RECT 1056.720 96.600 1056.980 96.860 ;
        RECT 603.160 43.900 603.420 44.160 ;
        RECT 1056.720 43.900 1056.980 44.160 ;
      LAYER met2 ;
        RECT 1059.490 1221.010 1060.050 1228.680 ;
        RECT 1057.700 1220.870 1060.050 1221.010 ;
        RECT 1057.700 1159.390 1057.840 1220.870 ;
        RECT 1059.490 1219.680 1060.050 1220.870 ;
        RECT 1056.260 1159.070 1056.520 1159.390 ;
        RECT 1057.640 1159.070 1057.900 1159.390 ;
        RECT 1056.320 1014.550 1056.460 1159.070 ;
        RECT 1056.260 1014.230 1056.520 1014.550 ;
        RECT 1056.720 1014.230 1056.980 1014.550 ;
        RECT 1056.780 942.210 1056.920 1014.230 ;
        RECT 1056.320 942.070 1056.920 942.210 ;
        RECT 1056.320 869.710 1056.460 942.070 ;
        RECT 1056.260 869.390 1056.520 869.710 ;
        RECT 1056.720 869.390 1056.980 869.710 ;
        RECT 1056.780 814.370 1056.920 869.390 ;
        RECT 1056.320 814.230 1056.920 814.370 ;
        RECT 1056.320 787.090 1056.460 814.230 ;
        RECT 1056.260 786.770 1056.520 787.090 ;
        RECT 1056.260 786.090 1056.520 786.410 ;
        RECT 1056.320 724.530 1056.460 786.090 ;
        RECT 1056.260 724.210 1056.520 724.530 ;
        RECT 1057.180 724.210 1057.440 724.530 ;
        RECT 1057.240 688.570 1057.380 724.210 ;
        RECT 1056.780 688.430 1057.380 688.570 ;
        RECT 1056.780 651.850 1056.920 688.430 ;
        RECT 1056.320 651.710 1056.920 651.850 ;
        RECT 1056.320 627.970 1056.460 651.710 ;
        RECT 1056.260 627.650 1056.520 627.970 ;
        RECT 1056.720 627.310 1056.980 627.630 ;
        RECT 1056.780 531.750 1056.920 627.310 ;
        RECT 1056.720 531.430 1056.980 531.750 ;
        RECT 1056.720 530.410 1056.980 530.730 ;
        RECT 1056.780 475.990 1056.920 530.410 ;
        RECT 1056.720 475.670 1056.980 475.990 ;
        RECT 1056.720 427.730 1056.980 428.050 ;
        RECT 1056.780 373.050 1056.920 427.730 ;
        RECT 1056.320 372.910 1056.920 373.050 ;
        RECT 1056.320 372.630 1056.460 372.910 ;
        RECT 1056.260 372.310 1056.520 372.630 ;
        RECT 1056.720 324.710 1056.980 325.030 ;
        RECT 1056.780 324.350 1056.920 324.710 ;
        RECT 1056.720 324.030 1056.980 324.350 ;
        RECT 1057.640 276.090 1057.900 276.410 ;
        RECT 1057.700 236.630 1057.840 276.090 ;
        RECT 1057.640 236.310 1057.900 236.630 ;
        RECT 1056.260 227.810 1056.520 228.130 ;
        RECT 1056.320 138.030 1056.460 227.810 ;
        RECT 1056.260 137.710 1056.520 138.030 ;
        RECT 1056.720 96.570 1056.980 96.890 ;
        RECT 1056.780 44.190 1056.920 96.570 ;
        RECT 603.160 43.870 603.420 44.190 ;
        RECT 1056.720 43.870 1056.980 44.190 ;
        RECT 603.220 2.400 603.360 43.870 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1063.130 1196.700 1063.450 1196.760 ;
        RECT 1067.270 1196.700 1067.590 1196.760 ;
        RECT 1063.130 1196.560 1067.590 1196.700 ;
        RECT 1063.130 1196.500 1063.450 1196.560 ;
        RECT 1067.270 1196.500 1067.590 1196.560 ;
        RECT 621.070 43.760 621.390 43.820 ;
        RECT 1063.130 43.760 1063.450 43.820 ;
        RECT 621.070 43.620 1063.450 43.760 ;
        RECT 621.070 43.560 621.390 43.620 ;
        RECT 1063.130 43.560 1063.450 43.620 ;
      LAYER via ;
        RECT 1063.160 1196.500 1063.420 1196.760 ;
        RECT 1067.300 1196.500 1067.560 1196.760 ;
        RECT 621.100 43.560 621.360 43.820 ;
        RECT 1063.160 43.560 1063.420 43.820 ;
      LAYER met2 ;
        RECT 1068.690 1220.330 1069.250 1228.680 ;
        RECT 1067.360 1220.190 1069.250 1220.330 ;
        RECT 1067.360 1196.790 1067.500 1220.190 ;
        RECT 1068.690 1219.680 1069.250 1220.190 ;
        RECT 1063.160 1196.470 1063.420 1196.790 ;
        RECT 1067.300 1196.470 1067.560 1196.790 ;
        RECT 1063.220 43.850 1063.360 1196.470 ;
        RECT 621.100 43.530 621.360 43.850 ;
        RECT 1063.160 43.530 1063.420 43.850 ;
        RECT 621.160 2.400 621.300 43.530 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 115.530 37.980 115.850 38.040 ;
        RECT 807.830 37.980 808.150 38.040 ;
        RECT 115.530 37.840 808.150 37.980 ;
        RECT 115.530 37.780 115.850 37.840 ;
        RECT 807.830 37.780 808.150 37.840 ;
      LAYER via ;
        RECT 115.560 37.780 115.820 38.040 ;
        RECT 807.860 37.780 808.120 38.040 ;
      LAYER met2 ;
        RECT 809.250 1220.330 809.810 1228.680 ;
        RECT 807.920 1220.190 809.810 1220.330 ;
        RECT 807.920 38.070 808.060 1220.190 ;
        RECT 809.250 1219.680 809.810 1220.190 ;
        RECT 115.560 37.750 115.820 38.070 ;
        RECT 807.860 37.750 808.120 38.070 ;
        RECT 115.620 2.400 115.760 37.750 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 821.210 1220.330 821.770 1228.680 ;
        RECT 821.210 1220.190 822.320 1220.330 ;
        RECT 821.210 1219.680 821.770 1220.190 ;
        RECT 822.180 44.725 822.320 1220.190 ;
        RECT 139.470 44.355 139.750 44.725 ;
        RECT 822.110 44.355 822.390 44.725 ;
        RECT 139.540 2.400 139.680 44.355 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 139.470 44.400 139.750 44.680 ;
        RECT 822.110 44.400 822.390 44.680 ;
      LAYER met3 ;
        RECT 139.445 44.690 139.775 44.705 ;
        RECT 822.085 44.690 822.415 44.705 ;
        RECT 139.445 44.390 822.415 44.690 ;
        RECT 139.445 44.375 139.775 44.390 ;
        RECT 822.085 44.375 822.415 44.390 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 157.390 44.780 157.710 44.840 ;
        RECT 828.530 44.780 828.850 44.840 ;
        RECT 157.390 44.640 828.850 44.780 ;
        RECT 157.390 44.580 157.710 44.640 ;
        RECT 828.530 44.580 828.850 44.640 ;
      LAYER via ;
        RECT 157.420 44.580 157.680 44.840 ;
        RECT 828.560 44.580 828.820 44.840 ;
      LAYER met2 ;
        RECT 830.410 1220.330 830.970 1228.680 ;
        RECT 828.620 1220.190 830.970 1220.330 ;
        RECT 828.620 44.870 828.760 1220.190 ;
        RECT 830.410 1219.680 830.970 1220.190 ;
        RECT 157.420 44.550 157.680 44.870 ;
        RECT 828.560 44.550 828.820 44.870 ;
        RECT 157.480 2.400 157.620 44.550 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.970 1196.700 835.290 1196.760 ;
        RECT 838.190 1196.700 838.510 1196.760 ;
        RECT 834.970 1196.560 838.510 1196.700 ;
        RECT 834.970 1196.500 835.290 1196.560 ;
        RECT 838.190 1196.500 838.510 1196.560 ;
        RECT 174.870 18.940 175.190 19.000 ;
        RECT 834.970 18.940 835.290 19.000 ;
        RECT 174.870 18.800 835.290 18.940 ;
        RECT 174.870 18.740 175.190 18.800 ;
        RECT 834.970 18.740 835.290 18.800 ;
      LAYER via ;
        RECT 835.000 1196.500 835.260 1196.760 ;
        RECT 838.220 1196.500 838.480 1196.760 ;
        RECT 174.900 18.740 175.160 19.000 ;
        RECT 835.000 18.740 835.260 19.000 ;
      LAYER met2 ;
        RECT 839.610 1220.330 840.170 1228.680 ;
        RECT 838.280 1220.190 840.170 1220.330 ;
        RECT 838.280 1196.790 838.420 1220.190 ;
        RECT 839.610 1219.680 840.170 1220.190 ;
        RECT 835.000 1196.470 835.260 1196.790 ;
        RECT 838.220 1196.470 838.480 1196.790 ;
        RECT 835.060 19.030 835.200 1196.470 ;
        RECT 174.900 18.710 175.160 19.030 ;
        RECT 835.000 18.710 835.260 19.030 ;
        RECT 174.960 2.400 175.100 18.710 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 355.190 1214.380 355.510 1214.440 ;
        RECT 848.770 1214.380 849.090 1214.440 ;
        RECT 355.190 1214.240 849.090 1214.380 ;
        RECT 355.190 1214.180 355.510 1214.240 ;
        RECT 848.770 1214.180 849.090 1214.240 ;
        RECT 192.810 16.560 193.130 16.620 ;
        RECT 355.190 16.560 355.510 16.620 ;
        RECT 192.810 16.420 355.510 16.560 ;
        RECT 192.810 16.360 193.130 16.420 ;
        RECT 355.190 16.360 355.510 16.420 ;
      LAYER via ;
        RECT 355.220 1214.180 355.480 1214.440 ;
        RECT 848.800 1214.180 849.060 1214.440 ;
        RECT 192.840 16.360 193.100 16.620 ;
        RECT 355.220 16.360 355.480 16.620 ;
      LAYER met2 ;
        RECT 848.810 1219.680 849.370 1228.680 ;
        RECT 848.860 1214.470 849.000 1219.680 ;
        RECT 355.220 1214.150 355.480 1214.470 ;
        RECT 848.800 1214.150 849.060 1214.470 ;
        RECT 355.280 16.650 355.420 1214.150 ;
        RECT 192.840 16.330 193.100 16.650 ;
        RECT 355.220 16.330 355.480 16.650 ;
        RECT 192.900 2.400 193.040 16.330 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.750 19.620 211.070 19.680 ;
        RECT 856.130 19.620 856.450 19.680 ;
        RECT 210.750 19.480 856.450 19.620 ;
        RECT 210.750 19.420 211.070 19.480 ;
        RECT 856.130 19.420 856.450 19.480 ;
      LAYER via ;
        RECT 210.780 19.420 211.040 19.680 ;
        RECT 856.160 19.420 856.420 19.680 ;
      LAYER met2 ;
        RECT 858.010 1220.330 858.570 1228.680 ;
        RECT 856.220 1220.190 858.570 1220.330 ;
        RECT 856.220 19.710 856.360 1220.190 ;
        RECT 858.010 1219.680 858.570 1220.190 ;
        RECT 210.780 19.390 211.040 19.710 ;
        RECT 856.160 19.390 856.420 19.710 ;
        RECT 210.840 2.400 210.980 19.390 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 375.890 1209.960 376.210 1210.020 ;
        RECT 867.170 1209.960 867.490 1210.020 ;
        RECT 375.890 1209.820 867.490 1209.960 ;
        RECT 375.890 1209.760 376.210 1209.820 ;
        RECT 867.170 1209.760 867.490 1209.820 ;
        RECT 228.690 16.220 229.010 16.280 ;
        RECT 375.890 16.220 376.210 16.280 ;
        RECT 228.690 16.080 376.210 16.220 ;
        RECT 228.690 16.020 229.010 16.080 ;
        RECT 375.890 16.020 376.210 16.080 ;
      LAYER via ;
        RECT 375.920 1209.760 376.180 1210.020 ;
        RECT 867.200 1209.760 867.460 1210.020 ;
        RECT 228.720 16.020 228.980 16.280 ;
        RECT 375.920 16.020 376.180 16.280 ;
      LAYER met2 ;
        RECT 867.210 1219.680 867.770 1228.680 ;
        RECT 867.260 1210.050 867.400 1219.680 ;
        RECT 375.920 1209.730 376.180 1210.050 ;
        RECT 867.200 1209.730 867.460 1210.050 ;
        RECT 375.980 16.310 376.120 1209.730 ;
        RECT 228.720 15.990 228.980 16.310 ;
        RECT 375.920 15.990 376.180 16.310 ;
        RECT 228.780 2.400 228.920 15.990 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 17.240 50.530 17.300 ;
        RECT 773.330 17.240 773.650 17.300 ;
        RECT 50.210 17.100 773.650 17.240 ;
        RECT 50.210 17.040 50.530 17.100 ;
        RECT 773.330 17.040 773.650 17.100 ;
      LAYER via ;
        RECT 50.240 17.040 50.500 17.300 ;
        RECT 773.360 17.040 773.620 17.300 ;
      LAYER met2 ;
        RECT 775.670 1220.330 776.230 1228.680 ;
        RECT 773.420 1220.190 776.230 1220.330 ;
        RECT 773.420 17.330 773.560 1220.190 ;
        RECT 775.670 1219.680 776.230 1220.190 ;
        RECT 50.240 17.010 50.500 17.330 ;
        RECT 773.360 17.010 773.620 17.330 ;
        RECT 50.300 2.400 50.440 17.010 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 389.690 1210.300 390.010 1210.360 ;
        RECT 879.130 1210.300 879.450 1210.360 ;
        RECT 389.690 1210.160 879.450 1210.300 ;
        RECT 389.690 1210.100 390.010 1210.160 ;
        RECT 879.130 1210.100 879.450 1210.160 ;
        RECT 252.610 15.880 252.930 15.940 ;
        RECT 389.690 15.880 390.010 15.940 ;
        RECT 252.610 15.740 390.010 15.880 ;
        RECT 252.610 15.680 252.930 15.740 ;
        RECT 389.690 15.680 390.010 15.740 ;
      LAYER via ;
        RECT 389.720 1210.100 389.980 1210.360 ;
        RECT 879.160 1210.100 879.420 1210.360 ;
        RECT 252.640 15.680 252.900 15.940 ;
        RECT 389.720 15.680 389.980 15.940 ;
      LAYER met2 ;
        RECT 879.170 1219.680 879.730 1228.680 ;
        RECT 879.220 1210.390 879.360 1219.680 ;
        RECT 389.720 1210.070 389.980 1210.390 ;
        RECT 879.160 1210.070 879.420 1210.390 ;
        RECT 389.780 15.970 389.920 1210.070 ;
        RECT 252.640 15.650 252.900 15.970 ;
        RECT 389.720 15.650 389.980 15.970 ;
        RECT 252.700 2.400 252.840 15.650 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 872.690 1208.260 873.010 1208.320 ;
        RECT 888.330 1208.260 888.650 1208.320 ;
        RECT 872.690 1208.120 888.650 1208.260 ;
        RECT 872.690 1208.060 873.010 1208.120 ;
        RECT 888.330 1208.060 888.650 1208.120 ;
        RECT 270.090 20.300 270.410 20.360 ;
        RECT 872.690 20.300 873.010 20.360 ;
        RECT 270.090 20.160 873.010 20.300 ;
        RECT 270.090 20.100 270.410 20.160 ;
        RECT 872.690 20.100 873.010 20.160 ;
      LAYER via ;
        RECT 872.720 1208.060 872.980 1208.320 ;
        RECT 888.360 1208.060 888.620 1208.320 ;
        RECT 270.120 20.100 270.380 20.360 ;
        RECT 872.720 20.100 872.980 20.360 ;
      LAYER met2 ;
        RECT 888.370 1219.680 888.930 1228.680 ;
        RECT 888.420 1208.350 888.560 1219.680 ;
        RECT 872.720 1208.030 872.980 1208.350 ;
        RECT 888.360 1208.030 888.620 1208.350 ;
        RECT 872.780 20.390 872.920 1208.030 ;
        RECT 270.120 20.070 270.380 20.390 ;
        RECT 872.720 20.070 872.980 20.390 ;
        RECT 270.180 2.400 270.320 20.070 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 424.190 1209.280 424.510 1209.340 ;
        RECT 897.530 1209.280 897.850 1209.340 ;
        RECT 424.190 1209.140 897.850 1209.280 ;
        RECT 424.190 1209.080 424.510 1209.140 ;
        RECT 897.530 1209.080 897.850 1209.140 ;
        RECT 288.030 15.540 288.350 15.600 ;
        RECT 424.190 15.540 424.510 15.600 ;
        RECT 288.030 15.400 424.510 15.540 ;
        RECT 288.030 15.340 288.350 15.400 ;
        RECT 424.190 15.340 424.510 15.400 ;
      LAYER via ;
        RECT 424.220 1209.080 424.480 1209.340 ;
        RECT 897.560 1209.080 897.820 1209.340 ;
        RECT 288.060 15.340 288.320 15.600 ;
        RECT 424.220 15.340 424.480 15.600 ;
      LAYER met2 ;
        RECT 897.570 1219.680 898.130 1228.680 ;
        RECT 897.620 1209.370 897.760 1219.680 ;
        RECT 424.220 1209.050 424.480 1209.370 ;
        RECT 897.560 1209.050 897.820 1209.370 ;
        RECT 424.280 15.630 424.420 1209.050 ;
        RECT 288.060 15.310 288.320 15.630 ;
        RECT 424.220 15.310 424.480 15.630 ;
        RECT 288.120 2.400 288.260 15.310 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 880.510 1212.340 880.830 1212.400 ;
        RECT 906.730 1212.340 907.050 1212.400 ;
        RECT 880.510 1212.200 907.050 1212.340 ;
        RECT 880.510 1212.140 880.830 1212.200 ;
        RECT 906.730 1212.140 907.050 1212.200 ;
        RECT 305.970 20.640 306.290 20.700 ;
        RECT 879.590 20.640 879.910 20.700 ;
        RECT 305.970 20.500 879.910 20.640 ;
        RECT 305.970 20.440 306.290 20.500 ;
        RECT 879.590 20.440 879.910 20.500 ;
      LAYER via ;
        RECT 880.540 1212.140 880.800 1212.400 ;
        RECT 906.760 1212.140 907.020 1212.400 ;
        RECT 306.000 20.440 306.260 20.700 ;
        RECT 879.620 20.440 879.880 20.700 ;
      LAYER met2 ;
        RECT 906.770 1219.680 907.330 1228.680 ;
        RECT 906.820 1212.430 906.960 1219.680 ;
        RECT 880.540 1212.110 880.800 1212.430 ;
        RECT 906.760 1212.110 907.020 1212.430 ;
        RECT 880.600 1192.450 880.740 1212.110 ;
        RECT 879.680 1192.310 880.740 1192.450 ;
        RECT 879.680 20.730 879.820 1192.310 ;
        RECT 306.000 20.410 306.260 20.730 ;
        RECT 879.620 20.410 879.880 20.730 ;
        RECT 306.060 2.400 306.200 20.410 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 534.590 1207.920 534.910 1207.980 ;
        RECT 915.930 1207.920 916.250 1207.980 ;
        RECT 534.590 1207.780 916.250 1207.920 ;
        RECT 534.590 1207.720 534.910 1207.780 ;
        RECT 915.930 1207.720 916.250 1207.780 ;
        RECT 323.910 14.520 324.230 14.580 ;
        RECT 534.590 14.520 534.910 14.580 ;
        RECT 323.910 14.380 534.910 14.520 ;
        RECT 323.910 14.320 324.230 14.380 ;
        RECT 534.590 14.320 534.910 14.380 ;
      LAYER via ;
        RECT 534.620 1207.720 534.880 1207.980 ;
        RECT 915.960 1207.720 916.220 1207.980 ;
        RECT 323.940 14.320 324.200 14.580 ;
        RECT 534.620 14.320 534.880 14.580 ;
      LAYER met2 ;
        RECT 915.970 1219.680 916.530 1228.680 ;
        RECT 916.020 1208.010 916.160 1219.680 ;
        RECT 534.620 1207.690 534.880 1208.010 ;
        RECT 915.960 1207.690 916.220 1208.010 ;
        RECT 534.680 14.610 534.820 1207.690 ;
        RECT 323.940 14.290 324.200 14.610 ;
        RECT 534.620 14.290 534.880 14.610 ;
        RECT 324.000 2.400 324.140 14.290 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 886.490 1209.960 886.810 1210.020 ;
        RECT 925.130 1209.960 925.450 1210.020 ;
        RECT 886.490 1209.820 925.450 1209.960 ;
        RECT 886.490 1209.760 886.810 1209.820 ;
        RECT 925.130 1209.760 925.450 1209.820 ;
        RECT 341.390 16.900 341.710 16.960 ;
        RECT 886.490 16.900 886.810 16.960 ;
        RECT 341.390 16.760 886.810 16.900 ;
        RECT 341.390 16.700 341.710 16.760 ;
        RECT 886.490 16.700 886.810 16.760 ;
      LAYER via ;
        RECT 886.520 1209.760 886.780 1210.020 ;
        RECT 925.160 1209.760 925.420 1210.020 ;
        RECT 341.420 16.700 341.680 16.960 ;
        RECT 886.520 16.700 886.780 16.960 ;
      LAYER met2 ;
        RECT 925.170 1219.680 925.730 1228.680 ;
        RECT 925.220 1210.050 925.360 1219.680 ;
        RECT 886.520 1209.730 886.780 1210.050 ;
        RECT 925.160 1209.730 925.420 1210.050 ;
        RECT 886.580 16.990 886.720 1209.730 ;
        RECT 341.420 16.670 341.680 16.990 ;
        RECT 886.520 16.670 886.780 16.990 ;
        RECT 341.480 2.400 341.620 16.670 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 916.465 1214.225 917.555 1214.395 ;
        RECT 916.465 1213.545 916.635 1214.225 ;
        RECT 917.385 1213.885 917.555 1214.225 ;
        RECT 921.065 1213.545 921.235 1215.075 ;
      LAYER mcon ;
        RECT 921.065 1214.905 921.235 1215.075 ;
      LAYER met1 ;
        RECT 921.005 1215.060 921.295 1215.105 ;
        RECT 934.330 1215.060 934.650 1215.120 ;
        RECT 921.005 1214.920 934.650 1215.060 ;
        RECT 921.005 1214.875 921.295 1214.920 ;
        RECT 934.330 1214.860 934.650 1214.920 ;
        RECT 917.325 1213.855 917.615 1214.085 ;
        RECT 431.090 1213.700 431.410 1213.760 ;
        RECT 916.405 1213.700 916.695 1213.745 ;
        RECT 431.090 1213.560 916.695 1213.700 ;
        RECT 917.400 1213.700 917.540 1213.855 ;
        RECT 921.005 1213.700 921.295 1213.745 ;
        RECT 917.400 1213.560 921.295 1213.700 ;
        RECT 431.090 1213.500 431.410 1213.560 ;
        RECT 916.405 1213.515 916.695 1213.560 ;
        RECT 921.005 1213.515 921.295 1213.560 ;
        RECT 359.330 14.860 359.650 14.920 ;
        RECT 431.090 14.860 431.410 14.920 ;
        RECT 359.330 14.720 431.410 14.860 ;
        RECT 359.330 14.660 359.650 14.720 ;
        RECT 431.090 14.660 431.410 14.720 ;
      LAYER via ;
        RECT 934.360 1214.860 934.620 1215.120 ;
        RECT 431.120 1213.500 431.380 1213.760 ;
        RECT 359.360 14.660 359.620 14.920 ;
        RECT 431.120 14.660 431.380 14.920 ;
      LAYER met2 ;
        RECT 934.370 1219.680 934.930 1228.680 ;
        RECT 934.420 1215.150 934.560 1219.680 ;
        RECT 934.360 1214.830 934.620 1215.150 ;
        RECT 431.120 1213.470 431.380 1213.790 ;
        RECT 431.180 14.950 431.320 1213.470 ;
        RECT 359.360 14.630 359.620 14.950 ;
        RECT 431.120 14.630 431.380 14.950 ;
        RECT 359.420 2.400 359.560 14.630 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 900.290 1212.680 900.610 1212.740 ;
        RECT 943.530 1212.680 943.850 1212.740 ;
        RECT 900.290 1212.540 943.850 1212.680 ;
        RECT 900.290 1212.480 900.610 1212.540 ;
        RECT 943.530 1212.480 943.850 1212.540 ;
        RECT 377.270 16.560 377.590 16.620 ;
        RECT 900.290 16.560 900.610 16.620 ;
        RECT 377.270 16.420 900.610 16.560 ;
        RECT 377.270 16.360 377.590 16.420 ;
        RECT 900.290 16.360 900.610 16.420 ;
      LAYER via ;
        RECT 900.320 1212.480 900.580 1212.740 ;
        RECT 943.560 1212.480 943.820 1212.740 ;
        RECT 377.300 16.360 377.560 16.620 ;
        RECT 900.320 16.360 900.580 16.620 ;
      LAYER met2 ;
        RECT 943.570 1219.680 944.130 1228.680 ;
        RECT 943.620 1212.770 943.760 1219.680 ;
        RECT 900.320 1212.450 900.580 1212.770 ;
        RECT 943.560 1212.450 943.820 1212.770 ;
        RECT 900.380 16.650 900.520 1212.450 ;
        RECT 377.300 16.330 377.560 16.650 ;
        RECT 900.320 16.330 900.580 16.650 ;
        RECT 377.360 2.400 377.500 16.330 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 893.925 1213.205 894.095 1214.395 ;
      LAYER mcon ;
        RECT 893.925 1214.225 894.095 1214.395 ;
      LAYER met1 ;
        RECT 893.865 1214.380 894.155 1214.425 ;
        RECT 952.730 1214.380 953.050 1214.440 ;
        RECT 893.865 1214.240 953.050 1214.380 ;
        RECT 893.865 1214.195 894.155 1214.240 ;
        RECT 952.730 1214.180 953.050 1214.240 ;
        RECT 444.890 1213.360 445.210 1213.420 ;
        RECT 893.865 1213.360 894.155 1213.405 ;
        RECT 444.890 1213.220 894.155 1213.360 ;
        RECT 444.890 1213.160 445.210 1213.220 ;
        RECT 893.865 1213.175 894.155 1213.220 ;
        RECT 395.210 14.180 395.530 14.240 ;
        RECT 444.890 14.180 445.210 14.240 ;
        RECT 395.210 14.040 445.210 14.180 ;
        RECT 395.210 13.980 395.530 14.040 ;
        RECT 444.890 13.980 445.210 14.040 ;
      LAYER via ;
        RECT 952.760 1214.180 953.020 1214.440 ;
        RECT 444.920 1213.160 445.180 1213.420 ;
        RECT 395.240 13.980 395.500 14.240 ;
        RECT 444.920 13.980 445.180 14.240 ;
      LAYER met2 ;
        RECT 952.770 1219.680 953.330 1228.680 ;
        RECT 952.820 1214.470 952.960 1219.680 ;
        RECT 952.760 1214.150 953.020 1214.470 ;
        RECT 444.920 1213.130 445.180 1213.450 ;
        RECT 444.980 14.270 445.120 1213.130 ;
        RECT 395.240 13.950 395.500 14.270 ;
        RECT 444.920 13.950 445.180 14.270 ;
        RECT 395.300 2.400 395.440 13.950 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 908.110 1210.980 908.430 1211.040 ;
        RECT 961.930 1210.980 962.250 1211.040 ;
        RECT 908.110 1210.840 962.250 1210.980 ;
        RECT 908.110 1210.780 908.430 1210.840 ;
        RECT 961.930 1210.780 962.250 1210.840 ;
        RECT 413.150 16.220 413.470 16.280 ;
        RECT 907.190 16.220 907.510 16.280 ;
        RECT 413.150 16.080 907.510 16.220 ;
        RECT 413.150 16.020 413.470 16.080 ;
        RECT 907.190 16.020 907.510 16.080 ;
      LAYER via ;
        RECT 908.140 1210.780 908.400 1211.040 ;
        RECT 961.960 1210.780 962.220 1211.040 ;
        RECT 413.180 16.020 413.440 16.280 ;
        RECT 907.220 16.020 907.480 16.280 ;
      LAYER met2 ;
        RECT 961.970 1219.680 962.530 1228.680 ;
        RECT 962.020 1211.070 962.160 1219.680 ;
        RECT 908.140 1210.750 908.400 1211.070 ;
        RECT 961.960 1210.750 962.220 1211.070 ;
        RECT 908.200 1191.770 908.340 1210.750 ;
        RECT 907.280 1191.630 908.340 1191.770 ;
        RECT 907.280 16.310 907.420 1191.630 ;
        RECT 413.180 15.990 413.440 16.310 ;
        RECT 907.220 15.990 907.480 16.310 ;
        RECT 413.240 2.400 413.380 15.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 86.090 1210.980 86.410 1211.040 ;
        RECT 787.590 1210.980 787.910 1211.040 ;
        RECT 86.090 1210.840 787.910 1210.980 ;
        RECT 86.090 1210.780 86.410 1210.840 ;
        RECT 787.590 1210.780 787.910 1210.840 ;
        RECT 74.130 19.960 74.450 20.020 ;
        RECT 86.090 19.960 86.410 20.020 ;
        RECT 74.130 19.820 86.410 19.960 ;
        RECT 74.130 19.760 74.450 19.820 ;
        RECT 86.090 19.760 86.410 19.820 ;
      LAYER via ;
        RECT 86.120 1210.780 86.380 1211.040 ;
        RECT 787.620 1210.780 787.880 1211.040 ;
        RECT 74.160 19.760 74.420 20.020 ;
        RECT 86.120 19.760 86.380 20.020 ;
      LAYER met2 ;
        RECT 787.630 1219.680 788.190 1228.680 ;
        RECT 787.680 1211.070 787.820 1219.680 ;
        RECT 86.120 1210.750 86.380 1211.070 ;
        RECT 787.620 1210.750 787.880 1211.070 ;
        RECT 86.180 20.050 86.320 1210.750 ;
        RECT 74.160 19.730 74.420 20.050 ;
        RECT 86.120 19.730 86.380 20.050 ;
        RECT 74.220 2.400 74.360 19.730 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 920.990 1212.340 921.310 1212.400 ;
        RECT 971.130 1212.340 971.450 1212.400 ;
        RECT 920.990 1212.200 971.450 1212.340 ;
        RECT 920.990 1212.140 921.310 1212.200 ;
        RECT 971.130 1212.140 971.450 1212.200 ;
        RECT 920.990 15.880 921.310 15.940 ;
        RECT 466.140 15.740 921.310 15.880 ;
        RECT 430.630 15.540 430.950 15.600 ;
        RECT 466.140 15.540 466.280 15.740 ;
        RECT 920.990 15.680 921.310 15.740 ;
        RECT 430.630 15.400 466.280 15.540 ;
        RECT 430.630 15.340 430.950 15.400 ;
      LAYER via ;
        RECT 921.020 1212.140 921.280 1212.400 ;
        RECT 971.160 1212.140 971.420 1212.400 ;
        RECT 430.660 15.340 430.920 15.600 ;
        RECT 921.020 15.680 921.280 15.940 ;
      LAYER met2 ;
        RECT 971.170 1219.680 971.730 1228.680 ;
        RECT 971.220 1212.430 971.360 1219.680 ;
        RECT 921.020 1212.110 921.280 1212.430 ;
        RECT 971.160 1212.110 971.420 1212.430 ;
        RECT 921.080 15.970 921.220 1212.110 ;
        RECT 921.020 15.650 921.280 15.970 ;
        RECT 430.660 15.310 430.920 15.630 ;
        RECT 430.720 2.400 430.860 15.310 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 465.590 1213.020 465.910 1213.080 ;
        RECT 980.330 1213.020 980.650 1213.080 ;
        RECT 465.590 1212.880 980.650 1213.020 ;
        RECT 465.590 1212.820 465.910 1212.880 ;
        RECT 980.330 1212.820 980.650 1212.880 ;
        RECT 448.570 15.880 448.890 15.940 ;
        RECT 465.590 15.880 465.910 15.940 ;
        RECT 448.570 15.740 465.910 15.880 ;
        RECT 448.570 15.680 448.890 15.740 ;
        RECT 465.590 15.680 465.910 15.740 ;
      LAYER via ;
        RECT 465.620 1212.820 465.880 1213.080 ;
        RECT 980.360 1212.820 980.620 1213.080 ;
        RECT 448.600 15.680 448.860 15.940 ;
        RECT 465.620 15.680 465.880 15.940 ;
      LAYER met2 ;
        RECT 980.370 1219.680 980.930 1228.680 ;
        RECT 980.420 1213.110 980.560 1219.680 ;
        RECT 465.620 1212.790 465.880 1213.110 ;
        RECT 980.360 1212.790 980.620 1213.110 ;
        RECT 465.680 15.970 465.820 1212.790 ;
        RECT 448.600 15.650 448.860 15.970 ;
        RECT 465.620 15.650 465.880 15.970 ;
        RECT 448.660 2.400 448.800 15.650 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 927.890 1211.660 928.210 1211.720 ;
        RECT 989.530 1211.660 989.850 1211.720 ;
        RECT 927.890 1211.520 989.850 1211.660 ;
        RECT 927.890 1211.460 928.210 1211.520 ;
        RECT 989.530 1211.460 989.850 1211.520 ;
        RECT 466.510 15.540 466.830 15.600 ;
        RECT 927.890 15.540 928.210 15.600 ;
        RECT 466.510 15.400 928.210 15.540 ;
        RECT 466.510 15.340 466.830 15.400 ;
        RECT 927.890 15.340 928.210 15.400 ;
      LAYER via ;
        RECT 927.920 1211.460 928.180 1211.720 ;
        RECT 989.560 1211.460 989.820 1211.720 ;
        RECT 466.540 15.340 466.800 15.600 ;
        RECT 927.920 15.340 928.180 15.600 ;
      LAYER met2 ;
        RECT 989.570 1219.680 990.130 1228.680 ;
        RECT 989.620 1211.750 989.760 1219.680 ;
        RECT 927.920 1211.430 928.180 1211.750 ;
        RECT 989.560 1211.430 989.820 1211.750 ;
        RECT 927.980 15.630 928.120 1211.430 ;
        RECT 466.540 15.310 466.800 15.630 ;
        RECT 927.920 15.310 928.180 15.630 ;
        RECT 466.600 2.400 466.740 15.310 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 565.945 1208.445 566.115 1214.055 ;
        RECT 613.785 1208.615 613.955 1214.055 ;
        RECT 662.545 1213.885 662.715 1214.735 ;
        RECT 711.305 1212.525 711.475 1214.735 ;
        RECT 762.365 1212.525 762.535 1214.055 ;
        RECT 810.665 1211.505 810.835 1214.055 ;
        RECT 858.965 1211.505 859.135 1214.395 ;
        RECT 917.845 1213.205 918.015 1215.415 ;
        RECT 953.265 1214.225 953.435 1215.415 ;
        RECT 613.325 1208.445 613.955 1208.615 ;
      LAYER mcon ;
        RECT 917.845 1215.245 918.015 1215.415 ;
        RECT 662.545 1214.565 662.715 1214.735 ;
        RECT 565.945 1213.885 566.115 1214.055 ;
        RECT 613.785 1213.885 613.955 1214.055 ;
        RECT 711.305 1214.565 711.475 1214.735 ;
        RECT 858.965 1214.225 859.135 1214.395 ;
        RECT 762.365 1213.885 762.535 1214.055 ;
        RECT 810.665 1213.885 810.835 1214.055 ;
        RECT 953.265 1215.245 953.435 1215.415 ;
      LAYER met1 ;
        RECT 917.785 1215.400 918.075 1215.445 ;
        RECT 953.205 1215.400 953.495 1215.445 ;
        RECT 917.785 1215.260 953.495 1215.400 ;
        RECT 917.785 1215.215 918.075 1215.260 ;
        RECT 953.205 1215.215 953.495 1215.260 ;
        RECT 662.485 1214.720 662.775 1214.765 ;
        RECT 711.245 1214.720 711.535 1214.765 ;
        RECT 662.485 1214.580 711.535 1214.720 ;
        RECT 662.485 1214.535 662.775 1214.580 ;
        RECT 711.245 1214.535 711.535 1214.580 ;
        RECT 858.905 1214.380 859.195 1214.425 ;
        RECT 953.205 1214.380 953.495 1214.425 ;
        RECT 998.270 1214.380 998.590 1214.440 ;
        RECT 858.905 1214.240 893.620 1214.380 ;
        RECT 858.905 1214.195 859.195 1214.240 ;
        RECT 517.110 1214.040 517.430 1214.100 ;
        RECT 565.885 1214.040 566.175 1214.085 ;
        RECT 517.110 1213.900 566.175 1214.040 ;
        RECT 517.110 1213.840 517.430 1213.900 ;
        RECT 565.885 1213.855 566.175 1213.900 ;
        RECT 613.725 1214.040 614.015 1214.085 ;
        RECT 662.485 1214.040 662.775 1214.085 ;
        RECT 613.725 1213.900 662.775 1214.040 ;
        RECT 613.725 1213.855 614.015 1213.900 ;
        RECT 662.485 1213.855 662.775 1213.900 ;
        RECT 762.305 1214.040 762.595 1214.085 ;
        RECT 810.605 1214.040 810.895 1214.085 ;
        RECT 762.305 1213.900 810.895 1214.040 ;
        RECT 893.480 1214.040 893.620 1214.240 ;
        RECT 953.205 1214.240 998.590 1214.380 ;
        RECT 953.205 1214.195 953.495 1214.240 ;
        RECT 998.270 1214.180 998.590 1214.240 ;
        RECT 916.850 1214.040 917.170 1214.100 ;
        RECT 893.480 1213.900 917.170 1214.040 ;
        RECT 762.305 1213.855 762.595 1213.900 ;
        RECT 810.605 1213.855 810.895 1213.900 ;
        RECT 916.850 1213.840 917.170 1213.900 ;
        RECT 917.310 1213.360 917.630 1213.420 ;
        RECT 917.785 1213.360 918.075 1213.405 ;
        RECT 917.310 1213.220 918.075 1213.360 ;
        RECT 917.310 1213.160 917.630 1213.220 ;
        RECT 917.785 1213.175 918.075 1213.220 ;
        RECT 711.245 1212.680 711.535 1212.725 ;
        RECT 762.305 1212.680 762.595 1212.725 ;
        RECT 711.245 1212.540 762.595 1212.680 ;
        RECT 711.245 1212.495 711.535 1212.540 ;
        RECT 762.305 1212.495 762.595 1212.540 ;
        RECT 810.605 1211.660 810.895 1211.705 ;
        RECT 858.905 1211.660 859.195 1211.705 ;
        RECT 810.605 1211.520 859.195 1211.660 ;
        RECT 810.605 1211.475 810.895 1211.520 ;
        RECT 858.905 1211.475 859.195 1211.520 ;
        RECT 493.190 1210.640 493.510 1210.700 ;
        RECT 517.110 1210.640 517.430 1210.700 ;
        RECT 493.190 1210.500 517.430 1210.640 ;
        RECT 493.190 1210.440 493.510 1210.500 ;
        RECT 517.110 1210.440 517.430 1210.500 ;
        RECT 565.885 1208.600 566.175 1208.645 ;
        RECT 613.265 1208.600 613.555 1208.645 ;
        RECT 565.885 1208.460 613.555 1208.600 ;
        RECT 565.885 1208.415 566.175 1208.460 ;
        RECT 613.265 1208.415 613.555 1208.460 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 493.190 15.200 493.510 15.260 ;
        RECT 484.450 15.060 493.510 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
        RECT 493.190 15.000 493.510 15.060 ;
      LAYER via ;
        RECT 517.140 1213.840 517.400 1214.100 ;
        RECT 998.300 1214.180 998.560 1214.440 ;
        RECT 916.880 1213.840 917.140 1214.100 ;
        RECT 917.340 1213.160 917.600 1213.420 ;
        RECT 493.220 1210.440 493.480 1210.700 ;
        RECT 517.140 1210.440 517.400 1210.700 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 493.220 15.000 493.480 15.260 ;
      LAYER met2 ;
        RECT 998.310 1219.680 998.870 1228.680 ;
        RECT 998.360 1214.470 998.500 1219.680 ;
        RECT 998.300 1214.150 998.560 1214.470 ;
        RECT 517.140 1213.810 517.400 1214.130 ;
        RECT 916.880 1213.810 917.140 1214.130 ;
        RECT 517.200 1210.730 517.340 1213.810 ;
        RECT 916.940 1213.530 917.080 1213.810 ;
        RECT 916.940 1213.450 917.540 1213.530 ;
        RECT 916.940 1213.390 917.600 1213.450 ;
        RECT 917.340 1213.130 917.600 1213.390 ;
        RECT 493.220 1210.410 493.480 1210.730 ;
        RECT 517.140 1210.410 517.400 1210.730 ;
        RECT 493.280 15.290 493.420 1210.410 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 493.220 14.970 493.480 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 935.710 1212.000 936.030 1212.060 ;
        RECT 1007.470 1212.000 1007.790 1212.060 ;
        RECT 935.710 1211.860 1007.790 1212.000 ;
        RECT 935.710 1211.800 936.030 1211.860 ;
        RECT 1007.470 1211.800 1007.790 1211.860 ;
        RECT 934.790 15.200 935.110 15.260 ;
        RECT 559.060 15.060 935.110 15.200 ;
        RECT 502.390 14.860 502.710 14.920 ;
        RECT 559.060 14.860 559.200 15.060 ;
        RECT 934.790 15.000 935.110 15.060 ;
        RECT 502.390 14.720 559.200 14.860 ;
        RECT 502.390 14.660 502.710 14.720 ;
      LAYER via ;
        RECT 935.740 1211.800 936.000 1212.060 ;
        RECT 1007.500 1211.800 1007.760 1212.060 ;
        RECT 502.420 14.660 502.680 14.920 ;
        RECT 934.820 15.000 935.080 15.260 ;
      LAYER met2 ;
        RECT 1007.510 1219.680 1008.070 1228.680 ;
        RECT 1007.560 1212.090 1007.700 1219.680 ;
        RECT 935.740 1211.770 936.000 1212.090 ;
        RECT 1007.500 1211.770 1007.760 1212.090 ;
        RECT 935.800 1192.450 935.940 1211.770 ;
        RECT 934.880 1192.310 935.940 1192.450 ;
        RECT 934.880 15.290 935.020 1192.310 ;
        RECT 934.820 14.970 935.080 15.290 ;
        RECT 502.420 14.630 502.680 14.950 ;
        RECT 502.480 2.400 502.620 14.630 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 1210.640 524.330 1210.700 ;
        RECT 1016.670 1210.640 1016.990 1210.700 ;
        RECT 524.010 1210.500 1016.990 1210.640 ;
        RECT 524.010 1210.440 524.330 1210.500 ;
        RECT 1016.670 1210.440 1016.990 1210.500 ;
        RECT 519.870 15.200 520.190 15.260 ;
        RECT 524.010 15.200 524.330 15.260 ;
        RECT 519.870 15.060 524.330 15.200 ;
        RECT 519.870 15.000 520.190 15.060 ;
        RECT 524.010 15.000 524.330 15.060 ;
      LAYER via ;
        RECT 524.040 1210.440 524.300 1210.700 ;
        RECT 1016.700 1210.440 1016.960 1210.700 ;
        RECT 519.900 15.000 520.160 15.260 ;
        RECT 524.040 15.000 524.300 15.260 ;
      LAYER met2 ;
        RECT 1016.710 1219.680 1017.270 1228.680 ;
        RECT 1016.760 1210.730 1016.900 1219.680 ;
        RECT 524.040 1210.410 524.300 1210.730 ;
        RECT 1016.700 1210.410 1016.960 1210.730 ;
        RECT 524.100 15.290 524.240 1210.410 ;
        RECT 519.900 14.970 520.160 15.290 ;
        RECT 524.040 14.970 524.300 15.290 ;
        RECT 519.960 2.400 520.100 14.970 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 1209.280 942.470 1209.340 ;
        RECT 1024.030 1209.280 1024.350 1209.340 ;
        RECT 942.150 1209.140 1024.350 1209.280 ;
        RECT 942.150 1209.080 942.470 1209.140 ;
        RECT 1024.030 1209.080 1024.350 1209.140 ;
        RECT 943.070 14.860 943.390 14.920 ;
        RECT 559.520 14.720 943.390 14.860 ;
        RECT 537.810 14.180 538.130 14.240 ;
        RECT 559.520 14.180 559.660 14.720 ;
        RECT 943.070 14.660 943.390 14.720 ;
        RECT 537.810 14.040 559.660 14.180 ;
        RECT 537.810 13.980 538.130 14.040 ;
      LAYER via ;
        RECT 942.180 1209.080 942.440 1209.340 ;
        RECT 1024.060 1209.080 1024.320 1209.340 ;
        RECT 537.840 13.980 538.100 14.240 ;
        RECT 943.100 14.660 943.360 14.920 ;
      LAYER met2 ;
        RECT 1025.910 1220.330 1026.470 1228.680 ;
        RECT 1024.120 1220.190 1026.470 1220.330 ;
        RECT 1024.120 1209.370 1024.260 1220.190 ;
        RECT 1025.910 1219.680 1026.470 1220.190 ;
        RECT 942.180 1209.050 942.440 1209.370 ;
        RECT 1024.060 1209.050 1024.320 1209.370 ;
        RECT 942.240 24.210 942.380 1209.050 ;
        RECT 942.240 24.070 943.300 24.210 ;
        RECT 943.160 14.950 943.300 24.070 ;
        RECT 943.100 14.630 943.360 14.950 ;
        RECT 537.840 13.950 538.100 14.270 ;
        RECT 537.900 2.400 538.040 13.950 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 1209.620 558.830 1209.680 ;
        RECT 1035.070 1209.620 1035.390 1209.680 ;
        RECT 558.510 1209.480 1035.390 1209.620 ;
        RECT 558.510 1209.420 558.830 1209.480 ;
        RECT 1035.070 1209.420 1035.390 1209.480 ;
        RECT 555.750 15.200 556.070 15.260 ;
        RECT 558.510 15.200 558.830 15.260 ;
        RECT 555.750 15.060 558.830 15.200 ;
        RECT 555.750 15.000 556.070 15.060 ;
        RECT 558.510 15.000 558.830 15.060 ;
      LAYER via ;
        RECT 558.540 1209.420 558.800 1209.680 ;
        RECT 1035.100 1209.420 1035.360 1209.680 ;
        RECT 555.780 15.000 556.040 15.260 ;
        RECT 558.540 15.000 558.800 15.260 ;
      LAYER met2 ;
        RECT 1035.110 1219.680 1035.670 1228.680 ;
        RECT 1035.160 1209.710 1035.300 1219.680 ;
        RECT 558.540 1209.390 558.800 1209.710 ;
        RECT 1035.100 1209.390 1035.360 1209.710 ;
        RECT 558.600 15.290 558.740 1209.390 ;
        RECT 555.780 14.970 556.040 15.290 ;
        RECT 558.540 14.970 558.800 15.290 ;
        RECT 555.840 2.400 555.980 14.970 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 1208.940 579.530 1209.000 ;
        RECT 1044.270 1208.940 1044.590 1209.000 ;
        RECT 579.210 1208.800 1044.590 1208.940 ;
        RECT 579.210 1208.740 579.530 1208.800 ;
        RECT 1044.270 1208.740 1044.590 1208.800 ;
        RECT 573.690 14.520 574.010 14.580 ;
        RECT 579.210 14.520 579.530 14.580 ;
        RECT 573.690 14.380 579.530 14.520 ;
        RECT 573.690 14.320 574.010 14.380 ;
        RECT 579.210 14.320 579.530 14.380 ;
      LAYER via ;
        RECT 579.240 1208.740 579.500 1209.000 ;
        RECT 1044.300 1208.740 1044.560 1209.000 ;
        RECT 573.720 14.320 573.980 14.580 ;
        RECT 579.240 14.320 579.500 14.580 ;
      LAYER met2 ;
        RECT 1044.310 1219.680 1044.870 1228.680 ;
        RECT 1044.360 1209.030 1044.500 1219.680 ;
        RECT 579.240 1208.710 579.500 1209.030 ;
        RECT 1044.300 1208.710 1044.560 1209.030 ;
        RECT 579.300 14.610 579.440 1208.710 ;
        RECT 573.720 14.290 573.980 14.610 ;
        RECT 579.240 14.290 579.500 14.610 ;
        RECT 573.780 2.400 573.920 14.290 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1003.865 1213.205 1004.035 1214.395 ;
        RECT 637.245 14.365 638.335 14.535 ;
        RECT 637.245 14.025 637.415 14.365 ;
      LAYER mcon ;
        RECT 1003.865 1214.225 1004.035 1214.395 ;
        RECT 638.165 14.365 638.335 14.535 ;
      LAYER met1 ;
        RECT 1003.805 1214.380 1004.095 1214.425 ;
        RECT 1053.470 1214.380 1053.790 1214.440 ;
        RECT 1003.805 1214.240 1053.790 1214.380 ;
        RECT 1003.805 1214.195 1004.095 1214.240 ;
        RECT 1053.470 1214.180 1053.790 1214.240 ;
        RECT 941.690 1213.360 942.010 1213.420 ;
        RECT 1003.805 1213.360 1004.095 1213.405 ;
        RECT 941.690 1213.220 1004.095 1213.360 ;
        RECT 941.690 1213.160 942.010 1213.220 ;
        RECT 1003.805 1213.175 1004.095 1213.220 ;
        RECT 638.105 14.520 638.395 14.565 ;
        RECT 941.690 14.520 942.010 14.580 ;
        RECT 638.105 14.380 942.010 14.520 ;
        RECT 638.105 14.335 638.395 14.380 ;
        RECT 941.690 14.320 942.010 14.380 ;
        RECT 591.170 14.180 591.490 14.240 ;
        RECT 637.185 14.180 637.475 14.225 ;
        RECT 591.170 14.040 637.475 14.180 ;
        RECT 591.170 13.980 591.490 14.040 ;
        RECT 637.185 13.995 637.475 14.040 ;
      LAYER via ;
        RECT 1053.500 1214.180 1053.760 1214.440 ;
        RECT 941.720 1213.160 941.980 1213.420 ;
        RECT 941.720 14.320 941.980 14.580 ;
        RECT 591.200 13.980 591.460 14.240 ;
      LAYER met2 ;
        RECT 1053.510 1219.680 1054.070 1228.680 ;
        RECT 1053.560 1214.470 1053.700 1219.680 ;
        RECT 1053.500 1214.150 1053.760 1214.470 ;
        RECT 941.720 1213.130 941.980 1213.450 ;
        RECT 941.780 14.610 941.920 1213.130 ;
        RECT 941.720 14.290 941.980 14.610 ;
        RECT 591.200 13.950 591.460 14.270 ;
        RECT 591.260 2.400 591.400 13.950 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 793.570 1196.700 793.890 1196.760 ;
        RECT 798.630 1196.700 798.950 1196.760 ;
        RECT 793.570 1196.560 798.950 1196.700 ;
        RECT 793.570 1196.500 793.890 1196.560 ;
        RECT 798.630 1196.500 798.950 1196.560 ;
        RECT 97.590 17.920 97.910 17.980 ;
        RECT 793.570 17.920 793.890 17.980 ;
        RECT 97.590 17.780 793.890 17.920 ;
        RECT 97.590 17.720 97.910 17.780 ;
        RECT 793.570 17.720 793.890 17.780 ;
      LAYER via ;
        RECT 793.600 1196.500 793.860 1196.760 ;
        RECT 798.660 1196.500 798.920 1196.760 ;
        RECT 97.620 17.720 97.880 17.980 ;
        RECT 793.600 17.720 793.860 17.980 ;
      LAYER met2 ;
        RECT 800.050 1220.330 800.610 1228.680 ;
        RECT 798.720 1220.190 800.610 1220.330 ;
        RECT 798.720 1196.790 798.860 1220.190 ;
        RECT 800.050 1219.680 800.610 1220.190 ;
        RECT 793.600 1196.470 793.860 1196.790 ;
        RECT 798.660 1196.470 798.920 1196.790 ;
        RECT 793.660 18.010 793.800 1196.470 ;
        RECT 97.620 17.690 97.880 18.010 ;
        RECT 793.600 17.690 793.860 18.010 ;
        RECT 97.680 2.400 97.820 17.690 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 1208.600 614.030 1208.660 ;
        RECT 1062.670 1208.600 1062.990 1208.660 ;
        RECT 613.710 1208.460 1062.990 1208.600 ;
        RECT 613.710 1208.400 614.030 1208.460 ;
        RECT 1062.670 1208.400 1062.990 1208.460 ;
        RECT 609.110 14.520 609.430 14.580 ;
        RECT 613.710 14.520 614.030 14.580 ;
        RECT 609.110 14.380 614.030 14.520 ;
        RECT 609.110 14.320 609.430 14.380 ;
        RECT 613.710 14.320 614.030 14.380 ;
      LAYER via ;
        RECT 613.740 1208.400 614.000 1208.660 ;
        RECT 1062.700 1208.400 1062.960 1208.660 ;
        RECT 609.140 14.320 609.400 14.580 ;
        RECT 613.740 14.320 614.000 14.580 ;
      LAYER met2 ;
        RECT 1062.710 1219.680 1063.270 1228.680 ;
        RECT 1062.760 1208.690 1062.900 1219.680 ;
        RECT 613.740 1208.370 614.000 1208.690 ;
        RECT 1062.700 1208.370 1062.960 1208.690 ;
        RECT 613.800 14.610 613.940 1208.370 ;
        RECT 609.140 14.290 609.400 14.610 ;
        RECT 613.740 14.290 614.000 14.610 ;
        RECT 609.200 2.400 609.340 14.290 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 955.490 1208.260 955.810 1208.320 ;
        RECT 1071.870 1208.260 1072.190 1208.320 ;
        RECT 955.490 1208.120 1072.190 1208.260 ;
        RECT 955.490 1208.060 955.810 1208.120 ;
        RECT 1071.870 1208.060 1072.190 1208.120 ;
        RECT 627.050 14.520 627.370 14.580 ;
        RECT 627.050 14.380 637.860 14.520 ;
        RECT 627.050 14.320 627.370 14.380 ;
        RECT 637.720 13.840 637.860 14.380 ;
        RECT 955.490 14.180 955.810 14.240 ;
        RECT 638.640 14.040 955.810 14.180 ;
        RECT 638.640 13.840 638.780 14.040 ;
        RECT 955.490 13.980 955.810 14.040 ;
        RECT 637.720 13.700 638.780 13.840 ;
      LAYER via ;
        RECT 955.520 1208.060 955.780 1208.320 ;
        RECT 1071.900 1208.060 1072.160 1208.320 ;
        RECT 627.080 14.320 627.340 14.580 ;
        RECT 955.520 13.980 955.780 14.240 ;
      LAYER met2 ;
        RECT 1071.910 1219.680 1072.470 1228.680 ;
        RECT 1071.960 1208.350 1072.100 1219.680 ;
        RECT 955.520 1208.030 955.780 1208.350 ;
        RECT 1071.900 1208.030 1072.160 1208.350 ;
        RECT 627.080 14.290 627.340 14.610 ;
        RECT 627.140 2.400 627.280 14.290 ;
        RECT 955.580 14.270 955.720 1208.030 ;
        RECT 955.520 13.950 955.780 14.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 141.290 1211.320 141.610 1211.380 ;
        RECT 811.970 1211.320 812.290 1211.380 ;
        RECT 141.290 1211.180 812.290 1211.320 ;
        RECT 141.290 1211.120 141.610 1211.180 ;
        RECT 811.970 1211.120 812.290 1211.180 ;
        RECT 121.510 19.620 121.830 19.680 ;
        RECT 141.290 19.620 141.610 19.680 ;
        RECT 121.510 19.480 141.610 19.620 ;
        RECT 121.510 19.420 121.830 19.480 ;
        RECT 141.290 19.420 141.610 19.480 ;
      LAYER via ;
        RECT 141.320 1211.120 141.580 1211.380 ;
        RECT 812.000 1211.120 812.260 1211.380 ;
        RECT 121.540 19.420 121.800 19.680 ;
        RECT 141.320 19.420 141.580 19.680 ;
      LAYER met2 ;
        RECT 812.010 1219.680 812.570 1228.680 ;
        RECT 812.060 1211.410 812.200 1219.680 ;
        RECT 141.320 1211.090 141.580 1211.410 ;
        RECT 812.000 1211.090 812.260 1211.410 ;
        RECT 141.380 19.710 141.520 1211.090 ;
        RECT 121.540 19.390 121.800 19.710 ;
        RECT 141.320 19.390 141.580 19.710 ;
        RECT 121.600 2.400 121.740 19.390 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 821.170 1173.920 821.490 1173.980 ;
        RECT 822.550 1173.920 822.870 1173.980 ;
        RECT 821.170 1173.780 822.870 1173.920 ;
        RECT 821.170 1173.720 821.490 1173.780 ;
        RECT 822.550 1173.720 822.870 1173.780 ;
        RECT 145.430 18.600 145.750 18.660 ;
        RECT 821.170 18.600 821.490 18.660 ;
        RECT 145.430 18.460 821.490 18.600 ;
        RECT 145.430 18.400 145.750 18.460 ;
        RECT 821.170 18.400 821.490 18.460 ;
      LAYER via ;
        RECT 821.200 1173.720 821.460 1173.980 ;
        RECT 822.580 1173.720 822.840 1173.980 ;
        RECT 145.460 18.400 145.720 18.660 ;
        RECT 821.200 18.400 821.460 18.660 ;
      LAYER met2 ;
        RECT 824.430 1220.330 824.990 1228.680 ;
        RECT 822.640 1220.190 824.990 1220.330 ;
        RECT 822.640 1174.010 822.780 1220.190 ;
        RECT 824.430 1219.680 824.990 1220.190 ;
        RECT 821.200 1173.690 821.460 1174.010 ;
        RECT 822.580 1173.690 822.840 1174.010 ;
        RECT 821.260 18.690 821.400 1173.690 ;
        RECT 145.460 18.370 145.720 18.690 ;
        RECT 821.200 18.370 821.460 18.690 ;
        RECT 145.520 2.400 145.660 18.370 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 1212.340 176.110 1212.400 ;
        RECT 833.590 1212.340 833.910 1212.400 ;
        RECT 175.790 1212.200 833.910 1212.340 ;
        RECT 175.790 1212.140 176.110 1212.200 ;
        RECT 833.590 1212.140 833.910 1212.200 ;
        RECT 163.370 16.900 163.690 16.960 ;
        RECT 175.790 16.900 176.110 16.960 ;
        RECT 163.370 16.760 176.110 16.900 ;
        RECT 163.370 16.700 163.690 16.760 ;
        RECT 175.790 16.700 176.110 16.760 ;
      LAYER via ;
        RECT 175.820 1212.140 176.080 1212.400 ;
        RECT 833.620 1212.140 833.880 1212.400 ;
        RECT 163.400 16.700 163.660 16.960 ;
        RECT 175.820 16.700 176.080 16.960 ;
      LAYER met2 ;
        RECT 833.630 1219.680 834.190 1228.680 ;
        RECT 833.680 1212.430 833.820 1219.680 ;
        RECT 175.820 1212.110 176.080 1212.430 ;
        RECT 833.620 1212.110 833.880 1212.430 ;
        RECT 175.880 16.990 176.020 1212.110 ;
        RECT 163.400 16.670 163.660 16.990 ;
        RECT 175.820 16.670 176.080 16.990 ;
        RECT 163.460 2.400 163.600 16.670 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 19.280 181.170 19.340 ;
        RECT 841.870 19.280 842.190 19.340 ;
        RECT 180.850 19.140 842.190 19.280 ;
        RECT 180.850 19.080 181.170 19.140 ;
        RECT 841.870 19.080 842.190 19.140 ;
      LAYER via ;
        RECT 180.880 19.080 181.140 19.340 ;
        RECT 841.900 19.080 842.160 19.340 ;
      LAYER met2 ;
        RECT 842.830 1220.330 843.390 1228.680 ;
        RECT 841.960 1220.190 843.390 1220.330 ;
        RECT 841.960 19.370 842.100 1220.190 ;
        RECT 842.830 1219.680 843.390 1220.190 ;
        RECT 180.880 19.050 181.140 19.370 ;
        RECT 841.900 19.050 842.160 19.370 ;
        RECT 180.940 2.400 181.080 19.050 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 241.645 1213.885 241.815 1214.735 ;
        RECT 289.485 1213.545 289.655 1214.735 ;
        RECT 338.245 1213.885 338.415 1214.735 ;
        RECT 303.285 1213.545 303.915 1213.715 ;
        RECT 386.085 1213.545 386.255 1214.735 ;
        RECT 410.465 1213.545 410.635 1214.735 ;
        RECT 434.385 1212.525 434.555 1214.735 ;
        RECT 448.185 1212.525 448.355 1214.055 ;
        RECT 472.565 1212.525 472.735 1214.055 ;
        RECT 517.645 1208.785 517.815 1212.695 ;
        RECT 565.485 1208.785 565.655 1212.695 ;
        RECT 710.845 1207.425 711.015 1212.695 ;
        RECT 762.825 1207.425 762.995 1212.695 ;
      LAYER mcon ;
        RECT 241.645 1214.565 241.815 1214.735 ;
        RECT 289.485 1214.565 289.655 1214.735 ;
        RECT 338.245 1214.565 338.415 1214.735 ;
        RECT 386.085 1214.565 386.255 1214.735 ;
        RECT 303.745 1213.545 303.915 1213.715 ;
        RECT 410.465 1214.565 410.635 1214.735 ;
        RECT 434.385 1214.565 434.555 1214.735 ;
        RECT 448.185 1213.885 448.355 1214.055 ;
        RECT 472.565 1213.885 472.735 1214.055 ;
        RECT 517.645 1212.525 517.815 1212.695 ;
        RECT 565.485 1212.525 565.655 1212.695 ;
        RECT 710.845 1212.525 711.015 1212.695 ;
        RECT 762.825 1212.525 762.995 1212.695 ;
      LAYER met1 ;
        RECT 241.585 1214.720 241.875 1214.765 ;
        RECT 289.425 1214.720 289.715 1214.765 ;
        RECT 241.585 1214.580 289.715 1214.720 ;
        RECT 241.585 1214.535 241.875 1214.580 ;
        RECT 289.425 1214.535 289.715 1214.580 ;
        RECT 338.185 1214.720 338.475 1214.765 ;
        RECT 386.025 1214.720 386.315 1214.765 ;
        RECT 338.185 1214.580 386.315 1214.720 ;
        RECT 338.185 1214.535 338.475 1214.580 ;
        RECT 386.025 1214.535 386.315 1214.580 ;
        RECT 410.405 1214.720 410.695 1214.765 ;
        RECT 434.325 1214.720 434.615 1214.765 ;
        RECT 410.405 1214.580 434.615 1214.720 ;
        RECT 410.405 1214.535 410.695 1214.580 ;
        RECT 434.325 1214.535 434.615 1214.580 ;
        RECT 210.290 1214.040 210.610 1214.100 ;
        RECT 241.585 1214.040 241.875 1214.085 ;
        RECT 338.185 1214.040 338.475 1214.085 ;
        RECT 210.290 1213.900 241.875 1214.040 ;
        RECT 210.290 1213.840 210.610 1213.900 ;
        RECT 241.585 1213.855 241.875 1213.900 ;
        RECT 309.740 1213.900 338.475 1214.040 ;
        RECT 289.425 1213.700 289.715 1213.745 ;
        RECT 303.225 1213.700 303.515 1213.745 ;
        RECT 289.425 1213.560 303.515 1213.700 ;
        RECT 289.425 1213.515 289.715 1213.560 ;
        RECT 303.225 1213.515 303.515 1213.560 ;
        RECT 303.685 1213.700 303.975 1213.745 ;
        RECT 309.740 1213.700 309.880 1213.900 ;
        RECT 338.185 1213.855 338.475 1213.900 ;
        RECT 448.125 1214.040 448.415 1214.085 ;
        RECT 472.505 1214.040 472.795 1214.085 ;
        RECT 448.125 1213.900 472.795 1214.040 ;
        RECT 448.125 1213.855 448.415 1213.900 ;
        RECT 472.505 1213.855 472.795 1213.900 ;
        RECT 303.685 1213.560 309.880 1213.700 ;
        RECT 386.025 1213.700 386.315 1213.745 ;
        RECT 410.405 1213.700 410.695 1213.745 ;
        RECT 386.025 1213.560 410.695 1213.700 ;
        RECT 303.685 1213.515 303.975 1213.560 ;
        RECT 386.025 1213.515 386.315 1213.560 ;
        RECT 410.405 1213.515 410.695 1213.560 ;
        RECT 434.325 1212.680 434.615 1212.725 ;
        RECT 448.125 1212.680 448.415 1212.725 ;
        RECT 434.325 1212.540 448.415 1212.680 ;
        RECT 434.325 1212.495 434.615 1212.540 ;
        RECT 448.125 1212.495 448.415 1212.540 ;
        RECT 472.505 1212.680 472.795 1212.725 ;
        RECT 517.585 1212.680 517.875 1212.725 ;
        RECT 472.505 1212.540 517.875 1212.680 ;
        RECT 472.505 1212.495 472.795 1212.540 ;
        RECT 517.585 1212.495 517.875 1212.540 ;
        RECT 565.425 1212.680 565.715 1212.725 ;
        RECT 565.870 1212.680 566.190 1212.740 ;
        RECT 565.425 1212.540 566.190 1212.680 ;
        RECT 565.425 1212.495 565.715 1212.540 ;
        RECT 565.870 1212.480 566.190 1212.540 ;
        RECT 613.710 1212.680 614.030 1212.740 ;
        RECT 710.785 1212.680 711.075 1212.725 ;
        RECT 613.710 1212.540 711.075 1212.680 ;
        RECT 613.710 1212.480 614.030 1212.540 ;
        RECT 710.785 1212.495 711.075 1212.540 ;
        RECT 762.765 1212.680 763.055 1212.725 ;
        RECT 851.990 1212.680 852.310 1212.740 ;
        RECT 762.765 1212.540 852.310 1212.680 ;
        RECT 762.765 1212.495 763.055 1212.540 ;
        RECT 851.990 1212.480 852.310 1212.540 ;
        RECT 517.585 1208.940 517.875 1208.985 ;
        RECT 565.425 1208.940 565.715 1208.985 ;
        RECT 517.585 1208.800 565.715 1208.940 ;
        RECT 517.585 1208.755 517.875 1208.800 ;
        RECT 565.425 1208.755 565.715 1208.800 ;
        RECT 565.870 1207.580 566.190 1207.640 ;
        RECT 613.250 1207.580 613.570 1207.640 ;
        RECT 565.870 1207.440 613.570 1207.580 ;
        RECT 565.870 1207.380 566.190 1207.440 ;
        RECT 613.250 1207.380 613.570 1207.440 ;
        RECT 710.785 1207.580 711.075 1207.625 ;
        RECT 762.765 1207.580 763.055 1207.625 ;
        RECT 710.785 1207.440 763.055 1207.580 ;
        RECT 710.785 1207.395 711.075 1207.440 ;
        RECT 762.765 1207.395 763.055 1207.440 ;
        RECT 198.790 20.640 199.110 20.700 ;
        RECT 210.290 20.640 210.610 20.700 ;
        RECT 198.790 20.500 210.610 20.640 ;
        RECT 198.790 20.440 199.110 20.500 ;
        RECT 210.290 20.440 210.610 20.500 ;
      LAYER via ;
        RECT 210.320 1213.840 210.580 1214.100 ;
        RECT 565.900 1212.480 566.160 1212.740 ;
        RECT 613.740 1212.480 614.000 1212.740 ;
        RECT 852.020 1212.480 852.280 1212.740 ;
        RECT 565.900 1207.380 566.160 1207.640 ;
        RECT 613.280 1207.380 613.540 1207.640 ;
        RECT 198.820 20.440 199.080 20.700 ;
        RECT 210.320 20.440 210.580 20.700 ;
      LAYER met2 ;
        RECT 852.030 1219.680 852.590 1228.680 ;
        RECT 210.320 1213.810 210.580 1214.130 ;
        RECT 210.380 20.730 210.520 1213.810 ;
        RECT 852.080 1212.770 852.220 1219.680 ;
        RECT 565.900 1212.450 566.160 1212.770 ;
        RECT 613.740 1212.450 614.000 1212.770 ;
        RECT 852.020 1212.450 852.280 1212.770 ;
        RECT 565.960 1207.670 566.100 1212.450 ;
        RECT 613.800 1209.450 613.940 1212.450 ;
        RECT 613.340 1209.310 613.940 1209.450 ;
        RECT 613.340 1207.670 613.480 1209.310 ;
        RECT 565.900 1207.350 566.160 1207.670 ;
        RECT 613.280 1207.350 613.540 1207.670 ;
        RECT 198.820 20.410 199.080 20.730 ;
        RECT 210.320 20.410 210.580 20.730 ;
        RECT 198.880 2.400 199.020 20.410 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.670 1196.700 855.990 1196.760 ;
        RECT 859.350 1196.700 859.670 1196.760 ;
        RECT 855.670 1196.560 859.670 1196.700 ;
        RECT 855.670 1196.500 855.990 1196.560 ;
        RECT 859.350 1196.500 859.670 1196.560 ;
        RECT 216.730 19.960 217.050 20.020 ;
        RECT 855.670 19.960 855.990 20.020 ;
        RECT 216.730 19.820 855.990 19.960 ;
        RECT 216.730 19.760 217.050 19.820 ;
        RECT 855.670 19.760 855.990 19.820 ;
      LAYER via ;
        RECT 855.700 1196.500 855.960 1196.760 ;
        RECT 859.380 1196.500 859.640 1196.760 ;
        RECT 216.760 19.760 217.020 20.020 ;
        RECT 855.700 19.760 855.960 20.020 ;
      LAYER met2 ;
        RECT 861.230 1220.330 861.790 1228.680 ;
        RECT 859.440 1220.190 861.790 1220.330 ;
        RECT 859.440 1196.790 859.580 1220.190 ;
        RECT 861.230 1219.680 861.790 1220.190 ;
        RECT 855.700 1196.470 855.960 1196.790 ;
        RECT 859.380 1196.470 859.640 1196.790 ;
        RECT 855.760 20.050 855.900 1196.470 ;
        RECT 216.760 19.730 217.020 20.050 ;
        RECT 855.700 19.730 855.960 20.050 ;
        RECT 216.820 2.400 216.960 19.730 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 479.390 1208.260 479.710 1208.320 ;
        RECT 870.390 1208.260 870.710 1208.320 ;
        RECT 479.390 1208.120 870.710 1208.260 ;
        RECT 479.390 1208.060 479.710 1208.120 ;
        RECT 870.390 1208.060 870.710 1208.120 ;
        RECT 234.670 15.200 234.990 15.260 ;
        RECT 479.390 15.200 479.710 15.260 ;
        RECT 234.670 15.060 479.710 15.200 ;
        RECT 234.670 15.000 234.990 15.060 ;
        RECT 479.390 15.000 479.710 15.060 ;
      LAYER via ;
        RECT 479.420 1208.060 479.680 1208.320 ;
        RECT 870.420 1208.060 870.680 1208.320 ;
        RECT 234.700 15.000 234.960 15.260 ;
        RECT 479.420 15.000 479.680 15.260 ;
      LAYER met2 ;
        RECT 870.430 1219.680 870.990 1228.680 ;
        RECT 870.480 1208.350 870.620 1219.680 ;
        RECT 479.420 1208.030 479.680 1208.350 ;
        RECT 870.420 1208.030 870.680 1208.350 ;
        RECT 479.480 15.290 479.620 1208.030 ;
        RECT 234.700 14.970 234.960 15.290 ;
        RECT 479.420 14.970 479.680 15.290 ;
        RECT 234.760 2.400 234.900 14.970 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 774.325 1110.865 774.495 1124.975 ;
        RECT 773.865 483.565 774.035 530.995 ;
        RECT 773.865 338.045 774.035 386.155 ;
        RECT 773.865 241.825 774.035 289.595 ;
        RECT 773.865 218.365 774.035 241.315 ;
        RECT 774.325 61.965 774.495 89.675 ;
      LAYER mcon ;
        RECT 774.325 1124.805 774.495 1124.975 ;
        RECT 773.865 530.825 774.035 530.995 ;
        RECT 773.865 385.985 774.035 386.155 ;
        RECT 773.865 289.425 774.035 289.595 ;
        RECT 773.865 241.145 774.035 241.315 ;
        RECT 774.325 89.505 774.495 89.675 ;
      LAYER met1 ;
        RECT 774.250 1124.960 774.570 1125.020 ;
        RECT 774.055 1124.820 774.570 1124.960 ;
        RECT 774.250 1124.760 774.570 1124.820 ;
        RECT 774.250 1111.020 774.570 1111.080 ;
        RECT 774.055 1110.880 774.570 1111.020 ;
        RECT 774.250 1110.820 774.570 1110.880 ;
        RECT 773.790 1062.740 774.110 1062.800 ;
        RECT 774.250 1062.740 774.570 1062.800 ;
        RECT 773.790 1062.600 774.570 1062.740 ;
        RECT 773.790 1062.540 774.110 1062.600 ;
        RECT 774.250 1062.540 774.570 1062.600 ;
        RECT 774.250 869.960 774.570 870.020 ;
        RECT 774.710 869.960 775.030 870.020 ;
        RECT 774.250 869.820 775.030 869.960 ;
        RECT 774.250 869.760 774.570 869.820 ;
        RECT 774.710 869.760 775.030 869.820 ;
        RECT 773.790 530.980 774.110 531.040 ;
        RECT 773.595 530.840 774.110 530.980 ;
        RECT 773.790 530.780 774.110 530.840 ;
        RECT 773.790 483.720 774.110 483.780 ;
        RECT 773.595 483.580 774.110 483.720 ;
        RECT 773.790 483.520 774.110 483.580 ;
        RECT 773.790 483.040 774.110 483.100 ;
        RECT 774.710 483.040 775.030 483.100 ;
        RECT 773.790 482.900 775.030 483.040 ;
        RECT 773.790 482.840 774.110 482.900 ;
        RECT 774.710 482.840 775.030 482.900 ;
        RECT 773.790 386.140 774.110 386.200 ;
        RECT 773.595 386.000 774.110 386.140 ;
        RECT 773.790 385.940 774.110 386.000 ;
        RECT 773.790 338.200 774.110 338.260 ;
        RECT 773.595 338.060 774.110 338.200 ;
        RECT 773.790 338.000 774.110 338.060 ;
        RECT 773.790 289.580 774.110 289.640 ;
        RECT 773.595 289.440 774.110 289.580 ;
        RECT 773.790 289.380 774.110 289.440 ;
        RECT 773.790 241.980 774.110 242.040 ;
        RECT 773.595 241.840 774.110 241.980 ;
        RECT 773.790 241.780 774.110 241.840 ;
        RECT 773.790 241.300 774.110 241.360 ;
        RECT 773.595 241.160 774.110 241.300 ;
        RECT 773.790 241.100 774.110 241.160 ;
        RECT 773.805 218.520 774.095 218.565 ;
        RECT 775.170 218.520 775.490 218.580 ;
        RECT 773.805 218.380 775.490 218.520 ;
        RECT 773.805 218.335 774.095 218.380 ;
        RECT 775.170 218.320 775.490 218.380 ;
        RECT 774.250 89.660 774.570 89.720 ;
        RECT 774.055 89.520 774.570 89.660 ;
        RECT 774.250 89.460 774.570 89.520 ;
        RECT 774.250 62.120 774.570 62.180 ;
        RECT 774.055 61.980 774.570 62.120 ;
        RECT 774.250 61.920 774.570 61.980 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 774.250 17.580 774.570 17.640 ;
        RECT 56.190 17.440 774.570 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 774.250 17.380 774.570 17.440 ;
      LAYER via ;
        RECT 774.280 1124.760 774.540 1125.020 ;
        RECT 774.280 1110.820 774.540 1111.080 ;
        RECT 773.820 1062.540 774.080 1062.800 ;
        RECT 774.280 1062.540 774.540 1062.800 ;
        RECT 774.280 869.760 774.540 870.020 ;
        RECT 774.740 869.760 775.000 870.020 ;
        RECT 773.820 530.780 774.080 531.040 ;
        RECT 773.820 483.520 774.080 483.780 ;
        RECT 773.820 482.840 774.080 483.100 ;
        RECT 774.740 482.840 775.000 483.100 ;
        RECT 773.820 385.940 774.080 386.200 ;
        RECT 773.820 338.000 774.080 338.260 ;
        RECT 773.820 289.380 774.080 289.640 ;
        RECT 773.820 241.780 774.080 242.040 ;
        RECT 773.820 241.100 774.080 241.360 ;
        RECT 775.200 218.320 775.460 218.580 ;
        RECT 774.280 89.460 774.540 89.720 ;
        RECT 774.280 61.920 774.540 62.180 ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 774.280 17.380 774.540 17.640 ;
      LAYER met2 ;
        RECT 778.430 1220.330 778.990 1228.680 ;
        RECT 776.640 1220.190 778.990 1220.330 ;
        RECT 776.640 1196.530 776.780 1220.190 ;
        RECT 778.430 1219.680 778.990 1220.190 ;
        RECT 774.340 1196.390 776.780 1196.530 ;
        RECT 774.340 1125.050 774.480 1196.390 ;
        RECT 774.280 1124.730 774.540 1125.050 ;
        RECT 774.340 1111.110 774.480 1111.265 ;
        RECT 774.280 1110.850 774.540 1111.110 ;
        RECT 773.880 1110.790 774.540 1110.850 ;
        RECT 773.880 1110.710 774.480 1110.790 ;
        RECT 773.880 1062.830 774.020 1110.710 ;
        RECT 773.820 1062.510 774.080 1062.830 ;
        RECT 774.280 1062.510 774.540 1062.830 ;
        RECT 774.340 980.290 774.480 1062.510 ;
        RECT 773.880 980.150 774.480 980.290 ;
        RECT 773.880 917.845 774.020 980.150 ;
        RECT 773.810 917.475 774.090 917.845 ;
        RECT 774.730 917.475 775.010 917.845 ;
        RECT 774.800 870.050 774.940 917.475 ;
        RECT 774.280 869.730 774.540 870.050 ;
        RECT 774.740 869.730 775.000 870.050 ;
        RECT 774.340 869.565 774.480 869.730 ;
        RECT 774.270 869.195 774.550 869.565 ;
        RECT 775.190 869.195 775.470 869.565 ;
        RECT 775.260 821.285 775.400 869.195 ;
        RECT 774.270 820.915 774.550 821.285 ;
        RECT 775.190 820.915 775.470 821.285 ;
        RECT 774.340 772.890 774.480 820.915 ;
        RECT 773.880 772.750 774.480 772.890 ;
        RECT 773.880 531.070 774.020 772.750 ;
        RECT 773.820 530.750 774.080 531.070 ;
        RECT 773.820 483.490 774.080 483.810 ;
        RECT 773.880 483.130 774.020 483.490 ;
        RECT 773.820 482.810 774.080 483.130 ;
        RECT 774.740 482.810 775.000 483.130 ;
        RECT 774.800 435.045 774.940 482.810 ;
        RECT 773.810 434.675 774.090 435.045 ;
        RECT 774.730 434.675 775.010 435.045 ;
        RECT 773.880 386.230 774.020 434.675 ;
        RECT 773.820 385.910 774.080 386.230 ;
        RECT 773.820 337.970 774.080 338.290 ;
        RECT 773.880 289.670 774.020 337.970 ;
        RECT 773.820 289.350 774.080 289.670 ;
        RECT 773.820 241.750 774.080 242.070 ;
        RECT 773.880 241.390 774.020 241.750 ;
        RECT 773.820 241.070 774.080 241.390 ;
        RECT 775.200 218.290 775.460 218.610 ;
        RECT 775.260 145.250 775.400 218.290 ;
        RECT 774.340 145.110 775.400 145.250 ;
        RECT 774.340 89.750 774.480 145.110 ;
        RECT 774.280 89.430 774.540 89.750 ;
        RECT 774.280 61.890 774.540 62.210 ;
        RECT 774.340 17.670 774.480 61.890 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 774.280 17.350 774.540 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 773.810 917.520 774.090 917.800 ;
        RECT 774.730 917.520 775.010 917.800 ;
        RECT 774.270 869.240 774.550 869.520 ;
        RECT 775.190 869.240 775.470 869.520 ;
        RECT 774.270 820.960 774.550 821.240 ;
        RECT 775.190 820.960 775.470 821.240 ;
        RECT 773.810 434.720 774.090 435.000 ;
        RECT 774.730 434.720 775.010 435.000 ;
      LAYER met3 ;
        RECT 773.785 917.810 774.115 917.825 ;
        RECT 774.705 917.810 775.035 917.825 ;
        RECT 773.785 917.510 775.035 917.810 ;
        RECT 773.785 917.495 774.115 917.510 ;
        RECT 774.705 917.495 775.035 917.510 ;
        RECT 774.245 869.530 774.575 869.545 ;
        RECT 775.165 869.530 775.495 869.545 ;
        RECT 774.245 869.230 775.495 869.530 ;
        RECT 774.245 869.215 774.575 869.230 ;
        RECT 775.165 869.215 775.495 869.230 ;
        RECT 774.245 821.250 774.575 821.265 ;
        RECT 775.165 821.250 775.495 821.265 ;
        RECT 774.245 820.950 775.495 821.250 ;
        RECT 774.245 820.935 774.575 820.950 ;
        RECT 775.165 820.935 775.495 820.950 ;
        RECT 773.785 435.010 774.115 435.025 ;
        RECT 774.705 435.010 775.035 435.025 ;
        RECT 773.785 434.710 775.035 435.010 ;
        RECT 773.785 434.695 774.115 434.710 ;
        RECT 774.705 434.695 775.035 434.710 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 120.590 1211.660 120.910 1211.720 ;
        RECT 790.810 1211.660 791.130 1211.720 ;
        RECT 120.590 1211.520 791.130 1211.660 ;
        RECT 120.590 1211.460 120.910 1211.520 ;
        RECT 790.810 1211.460 791.130 1211.520 ;
        RECT 80.110 18.600 80.430 18.660 ;
        RECT 120.590 18.600 120.910 18.660 ;
        RECT 80.110 18.460 120.910 18.600 ;
        RECT 80.110 18.400 80.430 18.460 ;
        RECT 120.590 18.400 120.910 18.460 ;
      LAYER via ;
        RECT 120.620 1211.460 120.880 1211.720 ;
        RECT 790.840 1211.460 791.100 1211.720 ;
        RECT 80.140 18.400 80.400 18.660 ;
        RECT 120.620 18.400 120.880 18.660 ;
      LAYER met2 ;
        RECT 790.850 1219.680 791.410 1228.680 ;
        RECT 790.900 1211.750 791.040 1219.680 ;
        RECT 120.620 1211.430 120.880 1211.750 ;
        RECT 790.840 1211.430 791.100 1211.750 ;
        RECT 120.680 18.690 120.820 1211.430 ;
        RECT 80.140 18.370 80.400 18.690 ;
        RECT 120.620 18.370 120.880 18.690 ;
        RECT 80.200 2.400 80.340 18.370 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 103.570 18.260 103.890 18.320 ;
        RECT 800.470 18.260 800.790 18.320 ;
        RECT 103.570 18.120 800.790 18.260 ;
        RECT 103.570 18.060 103.890 18.120 ;
        RECT 800.470 18.060 800.790 18.120 ;
      LAYER via ;
        RECT 103.600 18.060 103.860 18.320 ;
        RECT 800.500 18.060 800.760 18.320 ;
      LAYER met2 ;
        RECT 802.810 1220.330 803.370 1228.680 ;
        RECT 801.020 1220.190 803.370 1220.330 ;
        RECT 801.020 1196.700 801.160 1220.190 ;
        RECT 802.810 1219.680 803.370 1220.190 ;
        RECT 800.560 1196.560 801.160 1196.700 ;
        RECT 800.560 18.350 800.700 1196.560 ;
        RECT 103.600 18.030 103.860 18.350 ;
        RECT 800.500 18.030 800.760 18.350 ;
        RECT 103.660 2.400 103.800 18.030 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 155.090 1212.000 155.410 1212.060 ;
        RECT 815.190 1212.000 815.510 1212.060 ;
        RECT 155.090 1211.860 815.510 1212.000 ;
        RECT 155.090 1211.800 155.410 1211.860 ;
        RECT 815.190 1211.800 815.510 1211.860 ;
        RECT 127.490 18.940 127.810 19.000 ;
        RECT 155.090 18.940 155.410 19.000 ;
        RECT 127.490 18.800 155.410 18.940 ;
        RECT 127.490 18.740 127.810 18.800 ;
        RECT 155.090 18.740 155.410 18.800 ;
      LAYER via ;
        RECT 155.120 1211.800 155.380 1212.060 ;
        RECT 815.220 1211.800 815.480 1212.060 ;
        RECT 127.520 18.740 127.780 19.000 ;
        RECT 155.120 18.740 155.380 19.000 ;
      LAYER met2 ;
        RECT 815.230 1219.680 815.790 1228.680 ;
        RECT 815.280 1212.090 815.420 1219.680 ;
        RECT 155.120 1211.770 155.380 1212.090 ;
        RECT 815.220 1211.770 815.480 1212.090 ;
        RECT 155.180 19.030 155.320 1211.770 ;
        RECT 127.520 18.710 127.780 19.030 ;
        RECT 155.120 18.710 155.380 19.030 ;
        RECT 127.580 2.400 127.720 18.710 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 760.985 655.605 761.155 703.715 ;
        RECT 760.065 559.045 760.235 607.155 ;
        RECT 760.065 462.485 760.235 510.595 ;
        RECT 760.065 365.925 760.235 414.035 ;
      LAYER mcon ;
        RECT 760.985 703.545 761.155 703.715 ;
        RECT 760.065 606.985 760.235 607.155 ;
        RECT 760.065 510.425 760.235 510.595 ;
        RECT 760.065 413.865 760.235 414.035 ;
      LAYER met1 ;
        RECT 759.070 917.900 759.390 917.960 ;
        RECT 759.990 917.900 760.310 917.960 ;
        RECT 759.070 917.760 760.310 917.900 ;
        RECT 759.070 917.700 759.390 917.760 ;
        RECT 759.990 917.700 760.310 917.760 ;
        RECT 759.990 910.760 760.310 910.820 ;
        RECT 760.910 910.760 761.230 910.820 ;
        RECT 759.990 910.620 761.230 910.760 ;
        RECT 759.990 910.560 760.310 910.620 ;
        RECT 760.910 910.560 761.230 910.620 ;
        RECT 759.990 821.340 760.310 821.400 ;
        RECT 760.910 821.340 761.230 821.400 ;
        RECT 759.990 821.200 761.230 821.340 ;
        RECT 759.990 821.140 760.310 821.200 ;
        RECT 760.910 821.140 761.230 821.200 ;
        RECT 759.990 710.500 760.310 710.560 ;
        RECT 760.910 710.500 761.230 710.560 ;
        RECT 759.990 710.360 761.230 710.500 ;
        RECT 759.990 710.300 760.310 710.360 ;
        RECT 760.910 710.300 761.230 710.360 ;
        RECT 760.910 703.700 761.230 703.760 ;
        RECT 760.715 703.560 761.230 703.700 ;
        RECT 760.910 703.500 761.230 703.560 ;
        RECT 760.910 655.760 761.230 655.820 ;
        RECT 760.715 655.620 761.230 655.760 ;
        RECT 760.910 655.560 761.230 655.620 ;
        RECT 759.990 614.280 760.310 614.340 ;
        RECT 760.450 614.280 760.770 614.340 ;
        RECT 759.990 614.140 760.770 614.280 ;
        RECT 759.990 614.080 760.310 614.140 ;
        RECT 760.450 614.080 760.770 614.140 ;
        RECT 759.990 607.140 760.310 607.200 ;
        RECT 759.795 607.000 760.310 607.140 ;
        RECT 759.990 606.940 760.310 607.000 ;
        RECT 759.990 559.200 760.310 559.260 ;
        RECT 759.795 559.060 760.310 559.200 ;
        RECT 759.990 559.000 760.310 559.060 ;
        RECT 759.990 510.580 760.310 510.640 ;
        RECT 759.795 510.440 760.310 510.580 ;
        RECT 759.990 510.380 760.310 510.440 ;
        RECT 759.990 462.640 760.310 462.700 ;
        RECT 759.795 462.500 760.310 462.640 ;
        RECT 759.990 462.440 760.310 462.500 ;
        RECT 759.990 414.020 760.310 414.080 ;
        RECT 759.795 413.880 760.310 414.020 ;
        RECT 759.990 413.820 760.310 413.880 ;
        RECT 759.990 366.080 760.310 366.140 ;
        RECT 759.795 365.940 760.310 366.080 ;
        RECT 759.990 365.880 760.310 365.940 ;
        RECT 759.990 131.480 760.310 131.540 ;
        RECT 760.450 131.480 760.770 131.540 ;
        RECT 759.990 131.340 760.770 131.480 ;
        RECT 759.990 131.280 760.310 131.340 ;
        RECT 760.450 131.280 760.770 131.340 ;
      LAYER via ;
        RECT 759.100 917.700 759.360 917.960 ;
        RECT 760.020 917.700 760.280 917.960 ;
        RECT 760.020 910.560 760.280 910.820 ;
        RECT 760.940 910.560 761.200 910.820 ;
        RECT 760.020 821.140 760.280 821.400 ;
        RECT 760.940 821.140 761.200 821.400 ;
        RECT 760.020 710.300 760.280 710.560 ;
        RECT 760.940 710.300 761.200 710.560 ;
        RECT 760.940 703.500 761.200 703.760 ;
        RECT 760.940 655.560 761.200 655.820 ;
        RECT 760.020 614.080 760.280 614.340 ;
        RECT 760.480 614.080 760.740 614.340 ;
        RECT 760.020 606.940 760.280 607.200 ;
        RECT 760.020 559.000 760.280 559.260 ;
        RECT 760.020 510.380 760.280 510.640 ;
        RECT 760.020 462.440 760.280 462.700 ;
        RECT 760.020 413.820 760.280 414.080 ;
        RECT 760.020 365.880 760.280 366.140 ;
        RECT 760.020 131.280 760.280 131.540 ;
        RECT 760.480 131.280 760.740 131.540 ;
      LAYER met2 ;
        RECT 763.250 1220.330 763.810 1228.680 ;
        RECT 761.000 1220.190 763.810 1220.330 ;
        RECT 761.000 1196.530 761.140 1220.190 ;
        RECT 763.250 1219.680 763.810 1220.190 ;
        RECT 760.080 1196.390 761.140 1196.530 ;
        RECT 760.080 1172.730 760.220 1196.390 ;
        RECT 760.080 1172.590 760.680 1172.730 ;
        RECT 760.540 980.290 760.680 1172.590 ;
        RECT 760.080 980.150 760.680 980.290 ;
        RECT 760.080 966.125 760.220 980.150 ;
        RECT 759.090 965.755 759.370 966.125 ;
        RECT 760.010 965.755 760.290 966.125 ;
        RECT 759.160 917.990 759.300 965.755 ;
        RECT 759.100 917.670 759.360 917.990 ;
        RECT 760.020 917.670 760.280 917.990 ;
        RECT 760.080 910.850 760.220 917.670 ;
        RECT 760.020 910.530 760.280 910.850 ;
        RECT 760.940 910.530 761.200 910.850 ;
        RECT 761.000 821.430 761.140 910.530 ;
        RECT 760.020 821.110 760.280 821.430 ;
        RECT 760.940 821.110 761.200 821.430 ;
        RECT 760.080 710.590 760.220 821.110 ;
        RECT 760.020 710.270 760.280 710.590 ;
        RECT 760.940 710.270 761.200 710.590 ;
        RECT 761.000 703.790 761.140 710.270 ;
        RECT 760.940 703.470 761.200 703.790 ;
        RECT 760.940 655.530 761.200 655.850 ;
        RECT 761.000 621.930 761.140 655.530 ;
        RECT 760.540 621.790 761.140 621.930 ;
        RECT 760.540 614.370 760.680 621.790 ;
        RECT 760.020 614.050 760.280 614.370 ;
        RECT 760.480 614.050 760.740 614.370 ;
        RECT 760.080 607.230 760.220 614.050 ;
        RECT 760.020 606.910 760.280 607.230 ;
        RECT 760.020 558.970 760.280 559.290 ;
        RECT 760.080 510.670 760.220 558.970 ;
        RECT 760.020 510.350 760.280 510.670 ;
        RECT 760.020 462.410 760.280 462.730 ;
        RECT 760.080 414.110 760.220 462.410 ;
        RECT 760.020 413.790 760.280 414.110 ;
        RECT 760.020 365.850 760.280 366.170 ;
        RECT 760.080 131.570 760.220 365.850 ;
        RECT 760.020 131.250 760.280 131.570 ;
        RECT 760.480 131.250 760.740 131.570 ;
        RECT 760.540 76.005 760.680 131.250 ;
        RECT 760.470 75.635 760.750 76.005 ;
        RECT 761.390 75.635 761.670 76.005 ;
        RECT 761.460 28.405 761.600 75.635 ;
        RECT 760.010 28.035 760.290 28.405 ;
        RECT 761.390 28.035 761.670 28.405 ;
        RECT 760.080 16.845 760.220 28.035 ;
        RECT 26.310 16.475 26.590 16.845 ;
        RECT 760.010 16.475 760.290 16.845 ;
        RECT 26.380 2.400 26.520 16.475 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 759.090 965.800 759.370 966.080 ;
        RECT 760.010 965.800 760.290 966.080 ;
        RECT 760.470 75.680 760.750 75.960 ;
        RECT 761.390 75.680 761.670 75.960 ;
        RECT 760.010 28.080 760.290 28.360 ;
        RECT 761.390 28.080 761.670 28.360 ;
        RECT 26.310 16.520 26.590 16.800 ;
        RECT 760.010 16.520 760.290 16.800 ;
      LAYER met3 ;
        RECT 759.065 966.090 759.395 966.105 ;
        RECT 759.985 966.090 760.315 966.105 ;
        RECT 759.065 965.790 760.315 966.090 ;
        RECT 759.065 965.775 759.395 965.790 ;
        RECT 759.985 965.775 760.315 965.790 ;
        RECT 760.445 75.970 760.775 75.985 ;
        RECT 761.365 75.970 761.695 75.985 ;
        RECT 760.445 75.670 761.695 75.970 ;
        RECT 760.445 75.655 760.775 75.670 ;
        RECT 761.365 75.655 761.695 75.670 ;
        RECT 759.985 28.370 760.315 28.385 ;
        RECT 761.365 28.370 761.695 28.385 ;
        RECT 759.985 28.070 761.695 28.370 ;
        RECT 759.985 28.055 760.315 28.070 ;
        RECT 761.365 28.055 761.695 28.070 ;
        RECT 26.285 16.810 26.615 16.825 ;
        RECT 759.985 16.810 760.315 16.825 ;
        RECT 26.285 16.510 760.315 16.810 ;
        RECT 26.285 16.495 26.615 16.510 ;
        RECT 759.985 16.495 760.315 16.510 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.920 32.590 17.980 ;
        RECT 65.390 17.920 65.710 17.980 ;
        RECT 32.270 17.780 65.710 17.920 ;
        RECT 32.270 17.720 32.590 17.780 ;
        RECT 65.390 17.720 65.710 17.780 ;
      LAYER via ;
        RECT 32.300 17.720 32.560 17.980 ;
        RECT 65.420 17.720 65.680 17.980 ;
      LAYER met2 ;
        RECT 766.470 1219.680 767.030 1228.680 ;
        RECT 766.520 1210.925 766.660 1219.680 ;
        RECT 65.410 1210.555 65.690 1210.925 ;
        RECT 766.450 1210.555 766.730 1210.925 ;
        RECT 65.480 18.010 65.620 1210.555 ;
        RECT 32.300 17.690 32.560 18.010 ;
        RECT 65.420 17.690 65.680 18.010 ;
        RECT 32.360 2.400 32.500 17.690 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 65.410 1210.600 65.690 1210.880 ;
        RECT 766.450 1210.600 766.730 1210.880 ;
      LAYER met3 ;
        RECT 65.385 1210.890 65.715 1210.905 ;
        RECT 766.425 1210.890 766.755 1210.905 ;
        RECT 65.385 1210.590 766.755 1210.890 ;
        RECT 65.385 1210.575 65.715 1210.590 ;
        RECT 766.425 1210.575 766.755 1210.590 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 2735.680 907.020 3528.900 ;
        RECT 1084.020 2735.680 1087.020 3528.900 ;
        RECT 1264.020 2735.680 1267.020 3528.900 ;
        RECT 1444.020 2735.680 1447.020 3528.900 ;
        RECT 1624.020 2735.680 1627.020 3528.900 ;
        RECT 1804.020 2735.680 1807.020 3528.900 ;
        RECT 1984.020 2735.680 1987.020 3528.900 ;
        RECT 2164.020 2735.680 2167.020 3528.900 ;
        RECT 904.020 -9.220 907.020 1215.680 ;
        RECT 1084.020 -9.220 1087.020 1215.680 ;
        RECT 1264.020 -9.220 1267.020 1215.680 ;
        RECT 1444.020 -9.220 1447.020 1215.680 ;
        RECT 1624.020 -9.220 1627.020 1215.680 ;
        RECT 1804.020 -9.220 1807.020 1215.680 ;
        RECT 1984.020 -9.220 1987.020 1215.680 ;
        RECT 2164.020 -9.220 2167.020 1215.680 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 739.960 2712.380 ;
        RECT 2259.960 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 739.960 2532.380 ;
        RECT 2259.960 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 739.960 2352.380 ;
        RECT 2259.960 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 739.960 2172.380 ;
        RECT 2259.960 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 739.960 1992.380 ;
        RECT 2259.960 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 739.960 1812.380 ;
        RECT 2259.960 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 739.960 1632.380 ;
        RECT 2259.960 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 739.960 1452.380 ;
        RECT 2259.960 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 739.960 1272.380 ;
        RECT 2259.960 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 2735.680 817.020 3528.900 ;
        RECT 994.020 2735.680 997.020 3528.900 ;
        RECT 1174.020 2735.680 1177.020 3528.900 ;
        RECT 1354.020 2735.680 1357.020 3528.900 ;
        RECT 1534.020 2735.680 1537.020 3528.900 ;
        RECT 1714.020 2735.680 1717.020 3528.900 ;
        RECT 1894.020 2735.680 1897.020 3528.900 ;
        RECT 2074.020 2735.680 2077.020 3528.900 ;
        RECT 2254.020 2735.680 2257.020 3528.900 ;
        RECT 814.020 -9.220 817.020 1215.680 ;
        RECT 994.020 -9.220 997.020 1215.680 ;
        RECT 1174.020 -9.220 1177.020 1215.680 ;
        RECT 1354.020 -9.220 1357.020 1215.680 ;
        RECT 1534.020 -9.220 1537.020 1215.680 ;
        RECT 1714.020 -9.220 1717.020 1215.680 ;
        RECT 1894.020 -9.220 1897.020 1215.680 ;
        RECT 2074.020 -9.220 2077.020 1215.680 ;
        RECT 2254.020 -9.220 2257.020 1215.680 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 739.960 2622.380 ;
        RECT 2259.960 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 739.960 2442.380 ;
        RECT 2259.960 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 739.960 2262.380 ;
        RECT 2259.960 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 739.960 2082.380 ;
        RECT 2259.960 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 739.960 1902.380 ;
        RECT 2259.960 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 739.960 1722.380 ;
        RECT 2259.960 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 739.960 1542.380 ;
        RECT 2259.960 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 739.960 1362.380 ;
        RECT 2259.960 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 2735.680 745.020 3538.100 ;
        RECT 922.020 2735.680 925.020 3538.100 ;
        RECT 1102.020 2735.680 1105.020 3538.100 ;
        RECT 1282.020 2735.680 1285.020 3538.100 ;
        RECT 1462.020 2735.680 1465.020 3538.100 ;
        RECT 1642.020 2735.680 1645.020 3538.100 ;
        RECT 1822.020 2735.680 1825.020 3538.100 ;
        RECT 2002.020 2735.680 2005.020 3538.100 ;
        RECT 2182.020 2735.680 2185.020 3538.100 ;
        RECT 742.020 -18.420 745.020 1215.680 ;
        RECT 922.020 -18.420 925.020 1215.680 ;
        RECT 1102.020 -18.420 1105.020 1215.680 ;
        RECT 1282.020 -18.420 1285.020 1215.680 ;
        RECT 1462.020 -18.420 1465.020 1215.680 ;
        RECT 1642.020 -18.420 1645.020 1215.680 ;
        RECT 1822.020 -18.420 1825.020 1215.680 ;
        RECT 2002.020 -18.420 2005.020 1215.680 ;
        RECT 2182.020 -18.420 2185.020 1215.680 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 739.960 2730.380 ;
        RECT 2259.960 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 739.960 2550.380 ;
        RECT 2259.960 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 739.960 2370.380 ;
        RECT 2259.960 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 739.960 2190.380 ;
        RECT 2259.960 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 739.960 2010.380 ;
        RECT 2259.960 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 739.960 1830.380 ;
        RECT 2259.960 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 739.960 1650.380 ;
        RECT 2259.960 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 739.960 1470.380 ;
        RECT 2259.960 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 739.960 1290.380 ;
        RECT 2259.960 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 2735.680 835.020 3538.100 ;
        RECT 1012.020 2735.680 1015.020 3538.100 ;
        RECT 1192.020 2735.680 1195.020 3538.100 ;
        RECT 1372.020 2735.680 1375.020 3538.100 ;
        RECT 1552.020 2735.680 1555.020 3538.100 ;
        RECT 1732.020 2735.680 1735.020 3538.100 ;
        RECT 1912.020 2735.680 1915.020 3538.100 ;
        RECT 2092.020 2735.680 2095.020 3538.100 ;
        RECT 832.020 -18.420 835.020 1215.680 ;
        RECT 1012.020 -18.420 1015.020 1215.680 ;
        RECT 1192.020 -18.420 1195.020 1215.680 ;
        RECT 1372.020 -18.420 1375.020 1215.680 ;
        RECT 1552.020 -18.420 1555.020 1215.680 ;
        RECT 1732.020 -18.420 1735.020 1215.680 ;
        RECT 1912.020 -18.420 1915.020 1215.680 ;
        RECT 2092.020 -18.420 2095.020 1215.680 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 739.960 2640.380 ;
        RECT 2259.960 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 739.960 2460.380 ;
        RECT 2259.960 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 739.960 2280.380 ;
        RECT 2259.960 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 739.960 2100.380 ;
        RECT 2259.960 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 739.960 1920.380 ;
        RECT 2259.960 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 739.960 1740.380 ;
        RECT 2259.960 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 739.960 1560.380 ;
        RECT 2259.960 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 739.960 1380.380 ;
        RECT 2259.960 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 2735.680 763.020 3547.300 ;
        RECT 940.020 2735.680 943.020 3547.300 ;
        RECT 1120.020 2735.680 1123.020 3547.300 ;
        RECT 1300.020 2735.680 1303.020 3547.300 ;
        RECT 1480.020 2735.680 1483.020 3547.300 ;
        RECT 1660.020 2735.680 1663.020 3547.300 ;
        RECT 1840.020 2735.680 1843.020 3547.300 ;
        RECT 2020.020 2735.680 2023.020 3547.300 ;
        RECT 2200.020 2735.680 2203.020 3547.300 ;
        RECT 760.020 -27.620 763.020 1215.680 ;
        RECT 940.020 -27.620 943.020 1215.680 ;
        RECT 1120.020 -27.620 1123.020 1215.680 ;
        RECT 1300.020 -27.620 1303.020 1215.680 ;
        RECT 1480.020 -27.620 1483.020 1215.680 ;
        RECT 1660.020 -27.620 1663.020 1215.680 ;
        RECT 1840.020 -27.620 1843.020 1215.680 ;
        RECT 2020.020 -27.620 2023.020 1215.680 ;
        RECT 2200.020 -27.620 2203.020 1215.680 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 739.960 2568.380 ;
        RECT 2259.960 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 739.960 2388.380 ;
        RECT 2259.960 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 739.960 2208.380 ;
        RECT 2259.960 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 739.960 2028.380 ;
        RECT 2259.960 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 739.960 1848.380 ;
        RECT 2259.960 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 739.960 1668.380 ;
        RECT 2259.960 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 739.960 1488.380 ;
        RECT 2259.960 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 739.960 1308.380 ;
        RECT 2259.960 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 2735.680 853.020 3547.300 ;
        RECT 1030.020 2735.680 1033.020 3547.300 ;
        RECT 1210.020 2735.680 1213.020 3547.300 ;
        RECT 1390.020 2735.680 1393.020 3547.300 ;
        RECT 1570.020 2735.680 1573.020 3547.300 ;
        RECT 1750.020 2735.680 1753.020 3547.300 ;
        RECT 1930.020 2735.680 1933.020 3547.300 ;
        RECT 2110.020 2735.680 2113.020 3547.300 ;
        RECT 850.020 -27.620 853.020 1215.680 ;
        RECT 1030.020 -27.620 1033.020 1215.680 ;
        RECT 1210.020 -27.620 1213.020 1215.680 ;
        RECT 1390.020 -27.620 1393.020 1215.680 ;
        RECT 1570.020 -27.620 1573.020 1215.680 ;
        RECT 1750.020 -27.620 1753.020 1215.680 ;
        RECT 1930.020 -27.620 1933.020 1215.680 ;
        RECT 2110.020 -27.620 2113.020 1215.680 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 739.960 2658.380 ;
        RECT 2259.960 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 739.960 2478.380 ;
        RECT 2259.960 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 739.960 2298.380 ;
        RECT 2259.960 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 739.960 2118.380 ;
        RECT 2259.960 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 739.960 1938.380 ;
        RECT 2259.960 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 739.960 1758.380 ;
        RECT 2259.960 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 739.960 1578.380 ;
        RECT 2259.960 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 739.960 1398.380 ;
        RECT 2259.960 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 739.960 1218.380 ;
        RECT 2259.960 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 2735.680 781.020 3556.500 ;
        RECT 958.020 2735.680 961.020 3556.500 ;
        RECT 1138.020 2735.680 1141.020 3556.500 ;
        RECT 1318.020 2735.680 1321.020 3556.500 ;
        RECT 1498.020 2735.680 1501.020 3556.500 ;
        RECT 1678.020 2735.680 1681.020 3556.500 ;
        RECT 1858.020 2735.680 1861.020 3556.500 ;
        RECT 2038.020 2735.680 2041.020 3556.500 ;
        RECT 2218.020 2735.680 2221.020 3556.500 ;
        RECT 778.020 -36.820 781.020 1215.680 ;
        RECT 958.020 -36.820 961.020 1215.680 ;
        RECT 1138.020 -36.820 1141.020 1215.680 ;
        RECT 1318.020 -36.820 1321.020 1215.680 ;
        RECT 1498.020 -36.820 1501.020 1215.680 ;
        RECT 1678.020 -36.820 1681.020 1215.680 ;
        RECT 1858.020 -36.820 1861.020 1215.680 ;
        RECT 2038.020 -36.820 2041.020 1215.680 ;
        RECT 2218.020 -36.820 2221.020 1215.680 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 739.960 2586.380 ;
        RECT 2259.960 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 739.960 2406.380 ;
        RECT 2259.960 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 739.960 2226.380 ;
        RECT 2259.960 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 739.960 2046.380 ;
        RECT 2259.960 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 739.960 1866.380 ;
        RECT 2259.960 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 739.960 1686.380 ;
        RECT 2259.960 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 739.960 1506.380 ;
        RECT 2259.960 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 739.960 1326.380 ;
        RECT 2259.960 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 2735.680 871.020 3556.500 ;
        RECT 1048.020 2735.680 1051.020 3556.500 ;
        RECT 1228.020 2735.680 1231.020 3556.500 ;
        RECT 1408.020 2735.680 1411.020 3556.500 ;
        RECT 1588.020 2735.680 1591.020 3556.500 ;
        RECT 1768.020 2735.680 1771.020 3556.500 ;
        RECT 1948.020 2735.680 1951.020 3556.500 ;
        RECT 2128.020 2735.680 2131.020 3556.500 ;
        RECT 868.020 -36.820 871.020 1215.680 ;
        RECT 1048.020 -36.820 1051.020 1215.680 ;
        RECT 1228.020 -36.820 1231.020 1215.680 ;
        RECT 1408.020 -36.820 1411.020 1215.680 ;
        RECT 1588.020 -36.820 1591.020 1215.680 ;
        RECT 1768.020 -36.820 1771.020 1215.680 ;
        RECT 1948.020 -36.820 1951.020 1215.680 ;
        RECT 2128.020 -36.820 2131.020 1215.680 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 739.960 2676.380 ;
        RECT 2259.960 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 739.960 2496.380 ;
        RECT 2259.960 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 739.960 2316.380 ;
        RECT 2259.960 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 739.960 2136.380 ;
        RECT 2259.960 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 739.960 1956.380 ;
        RECT 2259.960 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 739.960 1776.380 ;
        RECT 2259.960 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 739.960 1596.380 ;
        RECT 2259.960 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 739.960 1416.380 ;
        RECT 2259.960 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 739.960 1236.380 ;
        RECT 2259.960 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 755.480 1236.475 2244.040 2713.605 ;
      LAYER met1 ;
        RECT 751.410 1236.320 2244.040 2713.760 ;
      LAYER met2 ;
        RECT 2230.190 2722.680 2230.750 2731.680 ;
        RECT 2243.070 2722.680 2243.630 2731.680 ;
      LAYER met2 ;
        RECT 751.440 2722.400 756.070 2722.680 ;
        RECT 757.190 2722.400 768.950 2722.680 ;
        RECT 770.070 2722.400 781.830 2722.680 ;
        RECT 782.950 2722.400 794.710 2722.680 ;
        RECT 795.830 2722.400 807.590 2722.680 ;
        RECT 808.710 2722.400 820.470 2722.680 ;
        RECT 821.590 2722.400 833.350 2722.680 ;
        RECT 834.470 2722.400 846.230 2722.680 ;
        RECT 847.350 2722.400 859.110 2722.680 ;
        RECT 860.230 2722.400 872.450 2722.680 ;
        RECT 873.570 2722.400 885.330 2722.680 ;
        RECT 886.450 2722.400 898.210 2722.680 ;
        RECT 899.330 2722.400 911.090 2722.680 ;
        RECT 912.210 2722.400 923.970 2722.680 ;
        RECT 925.090 2722.400 936.850 2722.680 ;
        RECT 937.970 2722.400 949.730 2722.680 ;
        RECT 950.850 2722.400 962.610 2722.680 ;
        RECT 963.730 2722.400 975.490 2722.680 ;
        RECT 976.610 2722.400 988.830 2722.680 ;
        RECT 989.950 2722.400 1001.710 2722.680 ;
        RECT 1002.830 2722.400 1014.590 2722.680 ;
        RECT 1015.710 2722.400 1027.470 2722.680 ;
        RECT 1028.590 2722.400 1040.350 2722.680 ;
        RECT 1041.470 2722.400 1053.230 2722.680 ;
        RECT 1054.350 2722.400 1066.110 2722.680 ;
        RECT 1067.230 2722.400 1078.990 2722.680 ;
        RECT 1080.110 2722.400 1091.870 2722.680 ;
        RECT 1092.990 2722.400 1105.210 2722.680 ;
        RECT 1106.330 2722.400 1118.090 2722.680 ;
        RECT 1119.210 2722.400 1130.970 2722.680 ;
        RECT 1132.090 2722.400 1143.850 2722.680 ;
        RECT 1144.970 2722.400 1156.730 2722.680 ;
        RECT 1157.850 2722.400 1169.610 2722.680 ;
        RECT 1170.730 2722.400 1182.490 2722.680 ;
        RECT 1183.610 2722.400 1195.370 2722.680 ;
        RECT 1196.490 2722.400 1208.250 2722.680 ;
        RECT 1209.370 2722.400 1221.590 2722.680 ;
        RECT 1222.710 2722.400 1234.470 2722.680 ;
        RECT 1235.590 2722.400 1247.350 2722.680 ;
        RECT 1248.470 2722.400 1260.230 2722.680 ;
        RECT 1261.350 2722.400 1273.110 2722.680 ;
        RECT 1274.230 2722.400 1285.990 2722.680 ;
        RECT 1287.110 2722.400 1298.870 2722.680 ;
        RECT 1299.990 2722.400 1311.750 2722.680 ;
        RECT 1312.870 2722.400 1324.630 2722.680 ;
        RECT 1325.750 2722.400 1337.970 2722.680 ;
        RECT 1339.090 2722.400 1350.850 2722.680 ;
        RECT 1351.970 2722.400 1363.730 2722.680 ;
        RECT 1364.850 2722.400 1376.610 2722.680 ;
        RECT 1377.730 2722.400 1389.490 2722.680 ;
        RECT 1390.610 2722.400 1402.370 2722.680 ;
        RECT 1403.490 2722.400 1415.250 2722.680 ;
        RECT 1416.370 2722.400 1428.130 2722.680 ;
        RECT 1429.250 2722.400 1441.010 2722.680 ;
        RECT 1442.130 2722.400 1454.350 2722.680 ;
        RECT 1455.470 2722.400 1467.230 2722.680 ;
        RECT 1468.350 2722.400 1480.110 2722.680 ;
        RECT 1481.230 2722.400 1492.990 2722.680 ;
        RECT 1494.110 2722.400 1505.870 2722.680 ;
        RECT 1506.990 2722.400 1518.750 2722.680 ;
        RECT 1519.870 2722.400 1531.630 2722.680 ;
        RECT 1532.750 2722.400 1544.510 2722.680 ;
        RECT 1545.630 2722.400 1557.390 2722.680 ;
        RECT 1558.510 2722.400 1570.730 2722.680 ;
        RECT 1571.850 2722.400 1583.610 2722.680 ;
        RECT 1584.730 2722.400 1596.490 2722.680 ;
        RECT 1597.610 2722.400 1609.370 2722.680 ;
        RECT 1610.490 2722.400 1622.250 2722.680 ;
        RECT 1623.370 2722.400 1635.130 2722.680 ;
        RECT 1636.250 2722.400 1648.010 2722.680 ;
        RECT 1649.130 2722.400 1660.890 2722.680 ;
        RECT 1662.010 2722.400 1673.770 2722.680 ;
        RECT 1674.890 2722.400 1687.110 2722.680 ;
        RECT 1688.230 2722.400 1699.990 2722.680 ;
        RECT 1701.110 2722.400 1712.870 2722.680 ;
        RECT 1713.990 2722.400 1725.750 2722.680 ;
        RECT 1726.870 2722.400 1738.630 2722.680 ;
        RECT 1739.750 2722.400 1751.510 2722.680 ;
        RECT 1752.630 2722.400 1764.390 2722.680 ;
        RECT 1765.510 2722.400 1777.270 2722.680 ;
        RECT 1778.390 2722.400 1790.150 2722.680 ;
        RECT 1791.270 2722.400 1803.490 2722.680 ;
        RECT 1804.610 2722.400 1816.370 2722.680 ;
        RECT 1817.490 2722.400 1829.250 2722.680 ;
        RECT 1830.370 2722.400 1842.130 2722.680 ;
        RECT 1843.250 2722.400 1855.010 2722.680 ;
        RECT 1856.130 2722.400 1867.890 2722.680 ;
        RECT 1869.010 2722.400 1880.770 2722.680 ;
        RECT 1881.890 2722.400 1893.650 2722.680 ;
        RECT 1894.770 2722.400 1906.530 2722.680 ;
        RECT 1907.650 2722.400 1919.870 2722.680 ;
        RECT 1920.990 2722.400 1932.750 2722.680 ;
        RECT 1933.870 2722.400 1945.630 2722.680 ;
        RECT 1946.750 2722.400 1958.510 2722.680 ;
        RECT 1959.630 2722.400 1971.390 2722.680 ;
        RECT 1972.510 2722.400 1984.270 2722.680 ;
        RECT 1985.390 2722.400 1997.150 2722.680 ;
        RECT 1998.270 2722.400 2010.030 2722.680 ;
        RECT 2011.150 2722.400 2022.910 2722.680 ;
        RECT 2024.030 2722.400 2036.250 2722.680 ;
        RECT 2037.370 2722.400 2049.130 2722.680 ;
        RECT 2050.250 2722.400 2062.010 2722.680 ;
        RECT 2063.130 2722.400 2074.890 2722.680 ;
        RECT 2076.010 2722.400 2087.770 2722.680 ;
        RECT 2088.890 2722.400 2100.650 2722.680 ;
        RECT 2101.770 2722.400 2113.530 2722.680 ;
        RECT 2114.650 2722.400 2126.410 2722.680 ;
        RECT 2127.530 2722.400 2139.290 2722.680 ;
        RECT 2140.410 2722.400 2152.630 2722.680 ;
        RECT 2153.750 2722.400 2165.510 2722.680 ;
        RECT 2166.630 2722.400 2178.390 2722.680 ;
        RECT 2179.510 2722.400 2191.270 2722.680 ;
        RECT 2192.390 2722.400 2204.150 2722.680 ;
        RECT 2205.270 2722.400 2217.030 2722.680 ;
        RECT 2218.150 2722.400 2229.910 2722.680 ;
        RECT 2231.030 2722.400 2242.560 2722.680 ;
        RECT 751.440 1228.960 2242.560 2722.400 ;
        RECT 752.130 1228.670 753.770 1228.960 ;
        RECT 754.890 1228.670 756.990 1228.960 ;
        RECT 758.110 1228.670 759.750 1228.960 ;
        RECT 760.870 1228.670 762.970 1228.960 ;
        RECT 764.090 1228.670 766.190 1228.960 ;
        RECT 767.310 1228.670 768.950 1228.960 ;
        RECT 770.070 1228.670 772.170 1228.960 ;
        RECT 773.290 1228.670 775.390 1228.960 ;
        RECT 776.510 1228.670 778.150 1228.960 ;
        RECT 779.270 1228.670 781.370 1228.960 ;
        RECT 782.490 1228.670 784.590 1228.960 ;
        RECT 785.710 1228.670 787.350 1228.960 ;
        RECT 788.470 1228.670 790.570 1228.960 ;
        RECT 791.690 1228.670 793.330 1228.960 ;
        RECT 794.450 1228.670 796.550 1228.960 ;
        RECT 797.670 1228.670 799.770 1228.960 ;
        RECT 800.890 1228.670 802.530 1228.960 ;
        RECT 803.650 1228.670 805.750 1228.960 ;
        RECT 806.870 1228.670 808.970 1228.960 ;
        RECT 810.090 1228.670 811.730 1228.960 ;
        RECT 812.850 1228.670 814.950 1228.960 ;
        RECT 816.070 1228.670 818.170 1228.960 ;
        RECT 819.290 1228.670 820.930 1228.960 ;
        RECT 822.050 1228.670 824.150 1228.960 ;
        RECT 825.270 1228.670 827.370 1228.960 ;
        RECT 828.490 1228.670 830.130 1228.960 ;
        RECT 831.250 1228.670 833.350 1228.960 ;
        RECT 834.470 1228.670 836.110 1228.960 ;
        RECT 837.230 1228.670 839.330 1228.960 ;
        RECT 840.450 1228.670 842.550 1228.960 ;
        RECT 843.670 1228.670 845.310 1228.960 ;
        RECT 846.430 1228.670 848.530 1228.960 ;
        RECT 849.650 1228.670 851.750 1228.960 ;
        RECT 852.870 1228.670 854.510 1228.960 ;
        RECT 855.630 1228.670 857.730 1228.960 ;
        RECT 858.850 1228.670 860.950 1228.960 ;
        RECT 862.070 1228.670 863.710 1228.960 ;
        RECT 864.830 1228.670 866.930 1228.960 ;
        RECT 868.050 1228.670 870.150 1228.960 ;
        RECT 871.270 1228.670 872.910 1228.960 ;
        RECT 874.030 1228.670 876.130 1228.960 ;
        RECT 877.250 1228.670 878.890 1228.960 ;
        RECT 880.010 1228.670 882.110 1228.960 ;
        RECT 883.230 1228.670 885.330 1228.960 ;
        RECT 886.450 1228.670 888.090 1228.960 ;
        RECT 889.210 1228.670 891.310 1228.960 ;
        RECT 892.430 1228.670 894.530 1228.960 ;
        RECT 895.650 1228.670 897.290 1228.960 ;
        RECT 898.410 1228.670 900.510 1228.960 ;
        RECT 901.630 1228.670 903.730 1228.960 ;
        RECT 904.850 1228.670 906.490 1228.960 ;
        RECT 907.610 1228.670 909.710 1228.960 ;
        RECT 910.830 1228.670 912.930 1228.960 ;
        RECT 914.050 1228.670 915.690 1228.960 ;
        RECT 916.810 1228.670 918.910 1228.960 ;
        RECT 920.030 1228.670 921.670 1228.960 ;
        RECT 922.790 1228.670 924.890 1228.960 ;
        RECT 926.010 1228.670 928.110 1228.960 ;
        RECT 929.230 1228.670 930.870 1228.960 ;
        RECT 931.990 1228.670 934.090 1228.960 ;
        RECT 935.210 1228.670 937.310 1228.960 ;
        RECT 938.430 1228.670 940.070 1228.960 ;
        RECT 941.190 1228.670 943.290 1228.960 ;
        RECT 944.410 1228.670 946.510 1228.960 ;
        RECT 947.630 1228.670 949.270 1228.960 ;
        RECT 950.390 1228.670 952.490 1228.960 ;
        RECT 953.610 1228.670 955.250 1228.960 ;
        RECT 956.370 1228.670 958.470 1228.960 ;
        RECT 959.590 1228.670 961.690 1228.960 ;
        RECT 962.810 1228.670 964.450 1228.960 ;
        RECT 965.570 1228.670 967.670 1228.960 ;
        RECT 968.790 1228.670 970.890 1228.960 ;
        RECT 972.010 1228.670 973.650 1228.960 ;
        RECT 974.770 1228.670 976.870 1228.960 ;
        RECT 977.990 1228.670 980.090 1228.960 ;
        RECT 981.210 1228.670 982.850 1228.960 ;
        RECT 983.970 1228.670 986.070 1228.960 ;
        RECT 987.190 1228.670 989.290 1228.960 ;
        RECT 990.410 1228.670 992.050 1228.960 ;
        RECT 993.170 1228.670 995.270 1228.960 ;
        RECT 996.390 1228.670 998.030 1228.960 ;
        RECT 999.150 1228.670 1001.250 1228.960 ;
        RECT 1002.370 1228.670 1004.470 1228.960 ;
        RECT 1005.590 1228.670 1007.230 1228.960 ;
        RECT 1008.350 1228.670 1010.450 1228.960 ;
        RECT 1011.570 1228.670 1013.670 1228.960 ;
        RECT 1014.790 1228.670 1016.430 1228.960 ;
        RECT 1017.550 1228.670 1019.650 1228.960 ;
        RECT 1020.770 1228.670 1022.870 1228.960 ;
        RECT 1023.990 1228.670 1025.630 1228.960 ;
        RECT 1026.750 1228.670 1028.850 1228.960 ;
        RECT 1029.970 1228.670 1032.070 1228.960 ;
        RECT 1033.190 1228.670 1034.830 1228.960 ;
        RECT 1035.950 1228.670 1038.050 1228.960 ;
        RECT 1039.170 1228.670 1040.810 1228.960 ;
        RECT 1041.930 1228.670 1044.030 1228.960 ;
        RECT 1045.150 1228.670 1047.250 1228.960 ;
        RECT 1048.370 1228.670 1050.010 1228.960 ;
        RECT 1051.130 1228.670 1053.230 1228.960 ;
        RECT 1054.350 1228.670 1056.450 1228.960 ;
        RECT 1057.570 1228.670 1059.210 1228.960 ;
        RECT 1060.330 1228.670 1062.430 1228.960 ;
        RECT 1063.550 1228.670 1065.650 1228.960 ;
        RECT 1066.770 1228.670 1068.410 1228.960 ;
        RECT 1069.530 1228.670 1071.630 1228.960 ;
        RECT 1072.750 1228.670 1074.850 1228.960 ;
        RECT 1075.970 1228.670 1077.610 1228.960 ;
        RECT 1078.730 1228.670 1080.830 1228.960 ;
        RECT 1081.950 1228.670 1083.590 1228.960 ;
        RECT 1084.710 1228.670 1086.810 1228.960 ;
        RECT 1087.930 1228.670 1090.030 1228.960 ;
        RECT 1091.150 1228.670 1092.790 1228.960 ;
        RECT 1093.910 1228.670 1096.010 1228.960 ;
        RECT 1097.130 1228.670 1099.230 1228.960 ;
        RECT 1100.350 1228.670 1101.990 1228.960 ;
        RECT 1103.110 1228.670 1105.210 1228.960 ;
        RECT 1106.330 1228.670 1108.430 1228.960 ;
        RECT 1109.550 1228.670 1111.190 1228.960 ;
        RECT 1112.310 1228.670 1114.410 1228.960 ;
        RECT 1115.530 1228.670 1117.170 1228.960 ;
        RECT 1118.290 1228.670 1120.390 1228.960 ;
        RECT 1121.510 1228.670 1123.610 1228.960 ;
        RECT 1124.730 1228.670 1126.370 1228.960 ;
        RECT 1127.490 1228.670 1129.590 1228.960 ;
        RECT 1130.710 1228.670 1132.810 1228.960 ;
        RECT 1133.930 1228.670 1135.570 1228.960 ;
        RECT 1136.690 1228.670 1138.790 1228.960 ;
        RECT 1139.910 1228.670 1142.010 1228.960 ;
        RECT 1143.130 1228.670 1144.770 1228.960 ;
        RECT 1145.890 1228.670 1147.990 1228.960 ;
        RECT 1149.110 1228.670 1151.210 1228.960 ;
        RECT 1152.330 1228.670 1153.970 1228.960 ;
        RECT 1155.090 1228.670 1157.190 1228.960 ;
        RECT 1158.310 1228.670 1159.950 1228.960 ;
        RECT 1161.070 1228.670 1163.170 1228.960 ;
        RECT 1164.290 1228.670 1166.390 1228.960 ;
        RECT 1167.510 1228.670 1169.150 1228.960 ;
        RECT 1170.270 1228.670 1172.370 1228.960 ;
        RECT 1173.490 1228.670 1175.590 1228.960 ;
        RECT 1176.710 1228.670 1178.350 1228.960 ;
        RECT 1179.470 1228.670 1181.570 1228.960 ;
        RECT 1182.690 1228.670 1184.790 1228.960 ;
        RECT 1185.910 1228.670 1187.550 1228.960 ;
        RECT 1188.670 1228.670 1190.770 1228.960 ;
        RECT 1191.890 1228.670 1193.990 1228.960 ;
        RECT 1195.110 1228.670 1196.750 1228.960 ;
        RECT 1197.870 1228.670 1199.970 1228.960 ;
        RECT 1201.090 1228.670 1202.730 1228.960 ;
        RECT 1203.850 1228.670 1205.950 1228.960 ;
        RECT 1207.070 1228.670 1209.170 1228.960 ;
        RECT 1210.290 1228.670 1211.930 1228.960 ;
        RECT 1213.050 1228.670 1215.150 1228.960 ;
        RECT 1216.270 1228.670 1218.370 1228.960 ;
        RECT 1219.490 1228.670 1221.130 1228.960 ;
        RECT 1222.250 1228.670 1224.350 1228.960 ;
        RECT 1225.470 1228.670 1227.570 1228.960 ;
        RECT 1228.690 1228.670 1230.330 1228.960 ;
        RECT 1231.450 1228.670 1233.550 1228.960 ;
        RECT 1234.670 1228.670 1236.770 1228.960 ;
        RECT 1237.890 1228.670 1239.530 1228.960 ;
        RECT 1240.650 1228.670 1242.750 1228.960 ;
        RECT 1243.870 1228.670 1245.510 1228.960 ;
        RECT 1246.630 1228.670 1248.730 1228.960 ;
        RECT 1249.850 1228.670 1251.950 1228.960 ;
        RECT 1253.070 1228.670 1254.710 1228.960 ;
        RECT 1255.830 1228.670 1257.930 1228.960 ;
        RECT 1259.050 1228.670 1261.150 1228.960 ;
        RECT 1262.270 1228.670 1263.910 1228.960 ;
        RECT 1265.030 1228.670 1267.130 1228.960 ;
        RECT 1268.250 1228.670 1270.350 1228.960 ;
        RECT 1271.470 1228.670 1273.110 1228.960 ;
        RECT 1274.230 1228.670 1276.330 1228.960 ;
        RECT 1277.450 1228.670 1279.090 1228.960 ;
        RECT 1280.210 1228.670 1282.310 1228.960 ;
        RECT 1283.430 1228.670 1285.530 1228.960 ;
        RECT 1286.650 1228.670 1288.290 1228.960 ;
        RECT 1289.410 1228.670 1291.510 1228.960 ;
        RECT 1292.630 1228.670 1294.730 1228.960 ;
        RECT 1295.850 1228.670 1297.490 1228.960 ;
        RECT 1298.610 1228.670 1300.710 1228.960 ;
        RECT 1301.830 1228.670 1303.930 1228.960 ;
        RECT 1305.050 1228.670 1306.690 1228.960 ;
        RECT 1307.810 1228.670 1309.910 1228.960 ;
        RECT 1311.030 1228.670 1313.130 1228.960 ;
        RECT 1314.250 1228.670 1315.890 1228.960 ;
        RECT 1317.010 1228.670 1319.110 1228.960 ;
        RECT 1320.230 1228.670 1321.870 1228.960 ;
        RECT 1322.990 1228.670 1325.090 1228.960 ;
        RECT 1326.210 1228.670 1328.310 1228.960 ;
        RECT 1329.430 1228.670 1331.070 1228.960 ;
        RECT 1332.190 1228.670 1334.290 1228.960 ;
        RECT 1335.410 1228.670 1337.510 1228.960 ;
        RECT 1338.630 1228.670 1340.270 1228.960 ;
        RECT 1341.390 1228.670 1343.490 1228.960 ;
        RECT 1344.610 1228.670 1346.710 1228.960 ;
        RECT 1347.830 1228.670 1349.470 1228.960 ;
        RECT 1350.590 1228.670 1352.690 1228.960 ;
        RECT 1353.810 1228.670 1355.910 1228.960 ;
        RECT 1357.030 1228.670 1358.670 1228.960 ;
        RECT 1359.790 1228.670 1361.890 1228.960 ;
        RECT 1363.010 1228.670 1364.650 1228.960 ;
        RECT 1365.770 1228.670 1367.870 1228.960 ;
        RECT 1368.990 1228.670 1371.090 1228.960 ;
        RECT 1372.210 1228.670 1373.850 1228.960 ;
        RECT 1374.970 1228.670 1377.070 1228.960 ;
        RECT 1378.190 1228.670 1380.290 1228.960 ;
        RECT 1381.410 1228.670 1383.050 1228.960 ;
        RECT 1384.170 1228.670 1386.270 1228.960 ;
        RECT 1387.390 1228.670 1389.490 1228.960 ;
        RECT 1390.610 1228.670 1392.250 1228.960 ;
        RECT 1393.370 1228.670 1395.470 1228.960 ;
        RECT 1396.590 1228.670 1398.690 1228.960 ;
        RECT 1399.810 1228.670 1401.450 1228.960 ;
        RECT 1402.570 1228.670 1404.670 1228.960 ;
        RECT 1405.790 1228.670 1407.430 1228.960 ;
        RECT 1408.550 1228.670 1410.650 1228.960 ;
        RECT 1411.770 1228.670 1413.870 1228.960 ;
        RECT 1414.990 1228.670 1416.630 1228.960 ;
        RECT 1417.750 1228.670 1419.850 1228.960 ;
        RECT 1420.970 1228.670 1423.070 1228.960 ;
        RECT 1424.190 1228.670 1425.830 1228.960 ;
        RECT 1426.950 1228.670 1429.050 1228.960 ;
        RECT 1430.170 1228.670 1432.270 1228.960 ;
        RECT 1433.390 1228.670 1435.030 1228.960 ;
        RECT 1436.150 1228.670 1438.250 1228.960 ;
        RECT 1439.370 1228.670 1441.010 1228.960 ;
        RECT 1442.130 1228.670 1444.230 1228.960 ;
        RECT 1445.350 1228.670 1447.450 1228.960 ;
        RECT 1448.570 1228.670 1450.210 1228.960 ;
        RECT 1451.330 1228.670 1453.430 1228.960 ;
        RECT 1454.550 1228.670 1456.650 1228.960 ;
        RECT 1457.770 1228.670 1459.410 1228.960 ;
        RECT 1460.530 1228.670 1462.630 1228.960 ;
        RECT 1463.750 1228.670 1465.850 1228.960 ;
        RECT 1466.970 1228.670 1468.610 1228.960 ;
        RECT 1469.730 1228.670 1471.830 1228.960 ;
        RECT 1472.950 1228.670 1475.050 1228.960 ;
        RECT 1476.170 1228.670 1477.810 1228.960 ;
        RECT 1478.930 1228.670 1481.030 1228.960 ;
        RECT 1482.150 1228.670 1483.790 1228.960 ;
        RECT 1484.910 1228.670 1487.010 1228.960 ;
        RECT 1488.130 1228.670 1490.230 1228.960 ;
        RECT 1491.350 1228.670 1492.990 1228.960 ;
        RECT 1494.110 1228.670 1496.210 1228.960 ;
        RECT 1497.330 1228.670 1499.430 1228.960 ;
        RECT 1500.550 1228.670 1502.190 1228.960 ;
        RECT 1503.310 1228.670 1505.410 1228.960 ;
        RECT 1506.530 1228.670 1508.630 1228.960 ;
        RECT 1509.750 1228.670 1511.390 1228.960 ;
        RECT 1512.510 1228.670 1514.610 1228.960 ;
        RECT 1515.730 1228.670 1517.830 1228.960 ;
        RECT 1518.950 1228.670 1520.590 1228.960 ;
        RECT 1521.710 1228.670 1523.810 1228.960 ;
        RECT 1524.930 1228.670 1526.570 1228.960 ;
        RECT 1527.690 1228.670 1529.790 1228.960 ;
        RECT 1530.910 1228.670 1533.010 1228.960 ;
        RECT 1534.130 1228.670 1535.770 1228.960 ;
        RECT 1536.890 1228.670 1538.990 1228.960 ;
        RECT 1540.110 1228.670 1542.210 1228.960 ;
        RECT 1543.330 1228.670 1544.970 1228.960 ;
        RECT 1546.090 1228.670 1548.190 1228.960 ;
        RECT 1549.310 1228.670 1551.410 1228.960 ;
        RECT 1552.530 1228.670 1554.170 1228.960 ;
        RECT 1555.290 1228.670 1557.390 1228.960 ;
        RECT 1558.510 1228.670 1560.610 1228.960 ;
        RECT 1561.730 1228.670 1563.370 1228.960 ;
        RECT 1564.490 1228.670 1566.590 1228.960 ;
        RECT 1567.710 1228.670 1569.350 1228.960 ;
        RECT 1570.470 1228.670 1572.570 1228.960 ;
        RECT 1573.690 1228.670 1575.790 1228.960 ;
        RECT 1576.910 1228.670 1578.550 1228.960 ;
        RECT 1579.670 1228.670 1581.770 1228.960 ;
        RECT 1582.890 1228.670 1584.990 1228.960 ;
        RECT 1586.110 1228.670 1587.750 1228.960 ;
        RECT 1588.870 1228.670 1590.970 1228.960 ;
        RECT 1592.090 1228.670 1594.190 1228.960 ;
        RECT 1595.310 1228.670 1596.950 1228.960 ;
        RECT 1598.070 1228.670 1600.170 1228.960 ;
        RECT 1601.290 1228.670 1602.930 1228.960 ;
        RECT 1604.050 1228.670 1606.150 1228.960 ;
        RECT 1607.270 1228.670 1609.370 1228.960 ;
        RECT 1610.490 1228.670 1612.130 1228.960 ;
        RECT 1613.250 1228.670 1615.350 1228.960 ;
        RECT 1616.470 1228.670 1618.570 1228.960 ;
        RECT 1619.690 1228.670 1621.330 1228.960 ;
        RECT 1622.450 1228.670 1624.550 1228.960 ;
        RECT 1625.670 1228.670 1627.770 1228.960 ;
        RECT 1628.890 1228.670 1630.530 1228.960 ;
        RECT 1631.650 1228.670 1633.750 1228.960 ;
        RECT 1634.870 1228.670 1636.970 1228.960 ;
        RECT 1638.090 1228.670 1639.730 1228.960 ;
        RECT 1640.850 1228.670 1642.950 1228.960 ;
        RECT 1644.070 1228.670 1645.710 1228.960 ;
        RECT 1646.830 1228.670 1648.930 1228.960 ;
        RECT 1650.050 1228.670 1652.150 1228.960 ;
        RECT 1653.270 1228.670 1654.910 1228.960 ;
        RECT 1656.030 1228.670 1658.130 1228.960 ;
        RECT 1659.250 1228.670 1661.350 1228.960 ;
        RECT 1662.470 1228.670 1664.110 1228.960 ;
        RECT 1665.230 1228.670 1667.330 1228.960 ;
        RECT 1668.450 1228.670 1670.550 1228.960 ;
        RECT 1671.670 1228.670 1673.310 1228.960 ;
        RECT 1674.430 1228.670 1676.530 1228.960 ;
        RECT 1677.650 1228.670 1679.750 1228.960 ;
        RECT 1680.870 1228.670 1682.510 1228.960 ;
        RECT 1683.630 1228.670 1685.730 1228.960 ;
        RECT 1686.850 1228.670 1688.490 1228.960 ;
        RECT 1689.610 1228.670 1691.710 1228.960 ;
        RECT 1692.830 1228.670 1694.930 1228.960 ;
        RECT 1696.050 1228.670 1697.690 1228.960 ;
        RECT 1698.810 1228.670 1700.910 1228.960 ;
        RECT 1702.030 1228.670 1704.130 1228.960 ;
        RECT 1705.250 1228.670 1706.890 1228.960 ;
        RECT 1708.010 1228.670 1710.110 1228.960 ;
        RECT 1711.230 1228.670 1713.330 1228.960 ;
        RECT 1714.450 1228.670 1716.090 1228.960 ;
        RECT 1717.210 1228.670 1719.310 1228.960 ;
        RECT 1720.430 1228.670 1722.530 1228.960 ;
        RECT 1723.650 1228.670 1725.290 1228.960 ;
        RECT 1726.410 1228.670 1728.510 1228.960 ;
        RECT 1729.630 1228.670 1731.270 1228.960 ;
        RECT 1732.390 1228.670 1734.490 1228.960 ;
        RECT 1735.610 1228.670 1737.710 1228.960 ;
        RECT 1738.830 1228.670 1740.470 1228.960 ;
        RECT 1741.590 1228.670 1743.690 1228.960 ;
        RECT 1744.810 1228.670 1746.910 1228.960 ;
        RECT 1748.030 1228.670 1749.670 1228.960 ;
        RECT 1750.790 1228.670 1752.890 1228.960 ;
        RECT 1754.010 1228.670 1756.110 1228.960 ;
        RECT 1757.230 1228.670 1758.870 1228.960 ;
        RECT 1759.990 1228.670 1762.090 1228.960 ;
        RECT 1763.210 1228.670 1764.850 1228.960 ;
        RECT 1765.970 1228.670 1768.070 1228.960 ;
        RECT 1769.190 1228.670 1771.290 1228.960 ;
        RECT 1772.410 1228.670 1774.050 1228.960 ;
        RECT 1775.170 1228.670 1777.270 1228.960 ;
        RECT 1778.390 1228.670 1780.490 1228.960 ;
        RECT 1781.610 1228.670 1783.250 1228.960 ;
        RECT 1784.370 1228.670 1786.470 1228.960 ;
        RECT 1787.590 1228.670 1789.690 1228.960 ;
        RECT 1790.810 1228.670 1792.450 1228.960 ;
        RECT 1793.570 1228.670 1795.670 1228.960 ;
        RECT 1796.790 1228.670 1798.890 1228.960 ;
        RECT 1800.010 1228.670 1801.650 1228.960 ;
        RECT 1802.770 1228.670 1804.870 1228.960 ;
        RECT 1805.990 1228.670 1807.630 1228.960 ;
        RECT 1808.750 1228.670 1810.850 1228.960 ;
        RECT 1811.970 1228.670 1814.070 1228.960 ;
        RECT 1815.190 1228.670 1816.830 1228.960 ;
        RECT 1817.950 1228.670 1820.050 1228.960 ;
        RECT 1821.170 1228.670 1823.270 1228.960 ;
        RECT 1824.390 1228.670 1826.030 1228.960 ;
        RECT 1827.150 1228.670 1829.250 1228.960 ;
        RECT 1830.370 1228.670 1832.470 1228.960 ;
        RECT 1833.590 1228.670 1835.230 1228.960 ;
        RECT 1836.350 1228.670 1838.450 1228.960 ;
        RECT 1839.570 1228.670 1841.670 1228.960 ;
        RECT 1842.790 1228.670 1844.430 1228.960 ;
        RECT 1845.550 1228.670 1847.650 1228.960 ;
        RECT 1848.770 1228.670 1850.410 1228.960 ;
        RECT 1851.530 1228.670 1853.630 1228.960 ;
        RECT 1854.750 1228.670 1856.850 1228.960 ;
        RECT 1857.970 1228.670 1859.610 1228.960 ;
        RECT 1860.730 1228.670 1862.830 1228.960 ;
        RECT 1863.950 1228.670 1866.050 1228.960 ;
        RECT 1867.170 1228.670 1868.810 1228.960 ;
        RECT 1869.930 1228.670 1872.030 1228.960 ;
        RECT 1873.150 1228.670 1875.250 1228.960 ;
        RECT 1876.370 1228.670 1878.010 1228.960 ;
        RECT 1879.130 1228.670 1881.230 1228.960 ;
        RECT 1882.350 1228.670 1884.450 1228.960 ;
        RECT 1885.570 1228.670 1887.210 1228.960 ;
        RECT 1888.330 1228.670 1890.430 1228.960 ;
        RECT 1891.550 1228.670 1893.190 1228.960 ;
        RECT 1894.310 1228.670 1896.410 1228.960 ;
        RECT 1897.530 1228.670 1899.630 1228.960 ;
        RECT 1900.750 1228.670 1902.390 1228.960 ;
        RECT 1903.510 1228.670 1905.610 1228.960 ;
        RECT 1906.730 1228.670 1908.830 1228.960 ;
        RECT 1909.950 1228.670 1911.590 1228.960 ;
        RECT 1912.710 1228.670 1914.810 1228.960 ;
        RECT 1915.930 1228.670 1918.030 1228.960 ;
        RECT 1919.150 1228.670 1920.790 1228.960 ;
        RECT 1921.910 1228.670 1924.010 1228.960 ;
        RECT 1925.130 1228.670 1926.770 1228.960 ;
        RECT 1927.890 1228.670 1929.990 1228.960 ;
        RECT 1931.110 1228.670 1933.210 1228.960 ;
        RECT 1934.330 1228.670 1935.970 1228.960 ;
        RECT 1937.090 1228.670 1939.190 1228.960 ;
        RECT 1940.310 1228.670 1942.410 1228.960 ;
        RECT 1943.530 1228.670 1945.170 1228.960 ;
        RECT 1946.290 1228.670 1948.390 1228.960 ;
        RECT 1949.510 1228.670 1951.610 1228.960 ;
        RECT 1952.730 1228.670 1954.370 1228.960 ;
        RECT 1955.490 1228.670 1957.590 1228.960 ;
        RECT 1958.710 1228.670 1960.810 1228.960 ;
        RECT 1961.930 1228.670 1963.570 1228.960 ;
        RECT 1964.690 1228.670 1966.790 1228.960 ;
        RECT 1967.910 1228.670 1969.550 1228.960 ;
        RECT 1970.670 1228.670 1972.770 1228.960 ;
        RECT 1973.890 1228.670 1975.990 1228.960 ;
        RECT 1977.110 1228.670 1978.750 1228.960 ;
        RECT 1979.870 1228.670 1981.970 1228.960 ;
        RECT 1983.090 1228.670 1985.190 1228.960 ;
        RECT 1986.310 1228.670 1987.950 1228.960 ;
        RECT 1989.070 1228.670 1991.170 1228.960 ;
        RECT 1992.290 1228.670 1994.390 1228.960 ;
        RECT 1995.510 1228.670 1997.150 1228.960 ;
        RECT 1998.270 1228.670 2000.370 1228.960 ;
        RECT 2001.490 1228.670 2003.590 1228.960 ;
        RECT 2004.710 1228.670 2006.350 1228.960 ;
        RECT 2007.470 1228.670 2009.570 1228.960 ;
        RECT 2010.690 1228.670 2012.330 1228.960 ;
        RECT 2013.450 1228.670 2015.550 1228.960 ;
        RECT 2016.670 1228.670 2018.770 1228.960 ;
        RECT 2019.890 1228.670 2021.530 1228.960 ;
        RECT 2022.650 1228.670 2024.750 1228.960 ;
        RECT 2025.870 1228.670 2027.970 1228.960 ;
        RECT 2029.090 1228.670 2030.730 1228.960 ;
        RECT 2031.850 1228.670 2033.950 1228.960 ;
        RECT 2035.070 1228.670 2037.170 1228.960 ;
        RECT 2038.290 1228.670 2039.930 1228.960 ;
        RECT 2041.050 1228.670 2043.150 1228.960 ;
        RECT 2044.270 1228.670 2046.370 1228.960 ;
        RECT 2047.490 1228.670 2049.130 1228.960 ;
        RECT 2050.250 1228.670 2052.350 1228.960 ;
        RECT 2053.470 1228.670 2055.110 1228.960 ;
        RECT 2056.230 1228.670 2058.330 1228.960 ;
        RECT 2059.450 1228.670 2061.550 1228.960 ;
        RECT 2062.670 1228.670 2064.310 1228.960 ;
        RECT 2065.430 1228.670 2067.530 1228.960 ;
        RECT 2068.650 1228.670 2070.750 1228.960 ;
        RECT 2071.870 1228.670 2073.510 1228.960 ;
        RECT 2074.630 1228.670 2076.730 1228.960 ;
        RECT 2077.850 1228.670 2079.950 1228.960 ;
        RECT 2081.070 1228.670 2082.710 1228.960 ;
        RECT 2083.830 1228.670 2085.930 1228.960 ;
        RECT 2087.050 1228.670 2088.690 1228.960 ;
        RECT 2089.810 1228.670 2091.910 1228.960 ;
        RECT 2093.030 1228.670 2095.130 1228.960 ;
        RECT 2096.250 1228.670 2097.890 1228.960 ;
        RECT 2099.010 1228.670 2101.110 1228.960 ;
        RECT 2102.230 1228.670 2104.330 1228.960 ;
        RECT 2105.450 1228.670 2107.090 1228.960 ;
        RECT 2108.210 1228.670 2110.310 1228.960 ;
        RECT 2111.430 1228.670 2113.530 1228.960 ;
        RECT 2114.650 1228.670 2116.290 1228.960 ;
        RECT 2117.410 1228.670 2119.510 1228.960 ;
        RECT 2120.630 1228.670 2122.730 1228.960 ;
        RECT 2123.850 1228.670 2125.490 1228.960 ;
        RECT 2126.610 1228.670 2128.710 1228.960 ;
        RECT 2129.830 1228.670 2131.470 1228.960 ;
        RECT 2132.590 1228.670 2134.690 1228.960 ;
        RECT 2135.810 1228.670 2137.910 1228.960 ;
        RECT 2139.030 1228.670 2140.670 1228.960 ;
        RECT 2141.790 1228.670 2143.890 1228.960 ;
        RECT 2145.010 1228.670 2147.110 1228.960 ;
        RECT 2148.230 1228.670 2149.870 1228.960 ;
        RECT 2150.990 1228.670 2153.090 1228.960 ;
        RECT 2154.210 1228.670 2156.310 1228.960 ;
        RECT 2157.430 1228.670 2159.070 1228.960 ;
        RECT 2160.190 1228.670 2162.290 1228.960 ;
        RECT 2163.410 1228.670 2165.510 1228.960 ;
        RECT 2166.630 1228.670 2168.270 1228.960 ;
        RECT 2169.390 1228.670 2171.490 1228.960 ;
        RECT 2172.610 1228.670 2174.250 1228.960 ;
        RECT 2175.370 1228.670 2177.470 1228.960 ;
        RECT 2178.590 1228.670 2180.690 1228.960 ;
        RECT 2181.810 1228.670 2183.450 1228.960 ;
        RECT 2184.570 1228.670 2186.670 1228.960 ;
        RECT 2187.790 1228.670 2189.890 1228.960 ;
        RECT 2191.010 1228.670 2192.650 1228.960 ;
        RECT 2193.770 1228.670 2195.870 1228.960 ;
        RECT 2196.990 1228.670 2199.090 1228.960 ;
        RECT 2200.210 1228.670 2201.850 1228.960 ;
        RECT 2202.970 1228.670 2205.070 1228.960 ;
        RECT 2206.190 1228.670 2208.290 1228.960 ;
        RECT 2209.410 1228.670 2211.050 1228.960 ;
        RECT 2212.170 1228.670 2214.270 1228.960 ;
        RECT 2215.390 1228.670 2217.030 1228.960 ;
        RECT 2218.150 1228.670 2220.250 1228.960 ;
        RECT 2221.370 1228.670 2223.470 1228.960 ;
        RECT 2224.590 1228.670 2226.230 1228.960 ;
        RECT 2227.350 1228.670 2229.450 1228.960 ;
        RECT 2230.570 1228.670 2232.670 1228.960 ;
        RECT 2233.790 1228.670 2235.430 1228.960 ;
        RECT 2236.550 1228.670 2238.650 1228.960 ;
        RECT 2239.770 1228.670 2241.870 1228.960 ;
      LAYER met2 ;
        RECT 2248.130 1219.680 2248.690 1228.680 ;
      LAYER met3 ;
        RECT 743.960 2537.140 752.960 2538.340 ;
        RECT 743.960 2162.460 752.960 2163.660 ;
        RECT 743.960 1787.100 752.960 1788.300 ;
        RECT 743.960 1412.420 752.960 1413.620 ;
      LAYER met3 ;
        RECT 771.000 1236.395 2231.800 2713.685 ;
      LAYER met3 ;
        RECT 2246.960 1975.460 2255.960 1976.660 ;
      LAYER met4 ;
        RECT 771.000 1236.320 2231.800 2713.760 ;
      LAYER met5 ;
        RECT 755.480 1328.760 2244.040 2708.980 ;
      LAYER met5 ;
        RECT 755.480 1290.465 2244.040 1292.065 ;
        RECT 755.480 1252.170 2244.040 1253.770 ;
  END
END user_project_wrapper
END LIBRARY

