magic
tech sky130A
magscale 1 2
timestamp 1606969352
<< checkpaint >>
rect -1260 -1260 14029 16173
<< viali >>
rect 4353 12257 4387 12291
rect 4537 12257 4571 12291
rect 5733 12257 5767 12291
rect 7573 12257 7607 12291
rect 8493 12257 8527 12291
rect 8677 12257 8711 12291
rect 10241 12257 10275 12291
rect 5549 12189 5583 12223
rect 6929 12189 6963 12223
rect 4629 12121 4663 12155
rect 8769 12121 8803 12155
rect 5917 12053 5951 12087
rect 10425 12053 10459 12087
rect 6837 11713 6871 11747
rect 3249 11645 3283 11679
rect 3433 11645 3467 11679
rect 4353 11645 4387 11679
rect 4629 11645 4663 11679
rect 4721 11645 4755 11679
rect 5641 11645 5675 11679
rect 5825 11645 5859 11679
rect 7021 11645 7055 11679
rect 8309 11645 8343 11679
rect 9321 11645 9355 11679
rect 9505 11645 9539 11679
rect 8125 11577 8159 11611
rect 8493 11577 8527 11611
rect 3249 11509 3283 11543
rect 5641 11509 5675 11543
rect 7205 11509 7239 11543
rect 9413 11509 9447 11543
rect 7849 11305 7883 11339
rect 9781 11305 9815 11339
rect 3157 11237 3191 11271
rect 2881 11169 2915 11203
rect 3065 11169 3099 11203
rect 4353 11169 4387 11203
rect 7297 11169 7331 11203
rect 7665 11169 7699 11203
rect 9689 11169 9723 11203
rect 9965 11169 9999 11203
rect 4077 11101 4111 11135
rect 5733 11101 5767 11135
rect 7757 11101 7791 11135
rect 8125 10761 8159 10795
rect 2237 10625 2271 10659
rect 3525 10625 3559 10659
rect 1869 10557 1903 10591
rect 2145 10557 2179 10591
rect 3249 10557 3283 10591
rect 3433 10557 3467 10591
rect 4445 10557 4479 10591
rect 4537 10557 4571 10591
rect 5641 10557 5675 10591
rect 5825 10557 5859 10591
rect 8125 10557 8159 10591
rect 8217 10557 8251 10591
rect 9229 10557 9263 10591
rect 9413 10557 9447 10591
rect 4721 10489 4755 10523
rect 6837 10489 6871 10523
rect 7021 10489 7055 10523
rect 7205 10489 7239 10523
rect 5641 10421 5675 10455
rect 9321 10421 9355 10455
rect 1869 10217 1903 10251
rect 6193 10217 6227 10251
rect 7481 10217 7515 10251
rect 8769 10217 8803 10251
rect 5181 10149 5215 10183
rect 6009 10149 6043 10183
rect 7297 10149 7331 10183
rect 1685 10081 1719 10115
rect 1869 10081 1903 10115
rect 2881 10081 2915 10115
rect 3065 10081 3099 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 7757 10081 7791 10115
rect 8585 10081 8619 10115
rect 9689 10081 9723 10115
rect 9965 10081 9999 10115
rect 3157 10013 3191 10047
rect 10057 10013 10091 10047
rect 6377 9945 6411 9979
rect 6193 9877 6227 9911
rect 7481 9877 7515 9911
rect 8769 9673 8803 9707
rect 7297 9605 7331 9639
rect 2329 9537 2363 9571
rect 2513 9469 2547 9503
rect 4353 9469 4387 9503
rect 4537 9469 4571 9503
rect 5457 9469 5491 9503
rect 5641 9469 5675 9503
rect 6929 9469 6963 9503
rect 8401 9469 8435 9503
rect 8585 9469 8619 9503
rect 9689 9401 9723 9435
rect 9873 9401 9907 9435
rect 10057 9401 10091 9435
rect 2697 9333 2731 9367
rect 4353 9333 4387 9367
rect 5825 9333 5859 9367
rect 1593 9061 1627 9095
rect 1961 9061 1995 9095
rect 3157 9061 3191 9095
rect 1777 8993 1811 9027
rect 2881 8993 2915 9027
rect 3065 8993 3099 9027
rect 4633 8993 4667 9027
rect 6561 8993 6595 9027
rect 7573 8993 7607 9027
rect 7665 8993 7699 9027
rect 9689 8993 9723 9027
rect 9873 8993 9907 9027
rect 4445 8925 4479 8959
rect 5733 8925 5767 8959
rect 6285 8925 6319 8959
rect 6745 8925 6779 8959
rect 4813 8789 4847 8823
rect 9781 8789 9815 8823
rect 3433 8585 3467 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 3801 8517 3835 8551
rect 8493 8517 8527 8551
rect 3525 8449 3559 8483
rect 5273 8449 5307 8483
rect 9229 8449 9263 8483
rect 10149 8449 10183 8483
rect 1501 8381 1535 8415
rect 3433 8381 3467 8415
rect 5365 8381 5399 8415
rect 5733 8381 5767 8415
rect 5917 8381 5951 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7297 8381 7331 8415
rect 7573 8381 7607 8415
rect 8769 8381 8803 8415
rect 10057 8381 10091 8415
rect 2145 8313 2179 8347
rect 4721 8313 4755 8347
rect 8677 8313 8711 8347
rect 6929 8245 6963 8279
rect 4261 8041 4295 8075
rect 8401 8041 8435 8075
rect 2973 7973 3007 8007
rect 9689 7973 9723 8007
rect 10241 7973 10275 8007
rect 1685 7905 1719 7939
rect 1869 7905 1903 7939
rect 2789 7905 2823 7939
rect 3157 7905 3191 7939
rect 4261 7905 4295 7939
rect 4445 7905 4479 7939
rect 4721 7905 4755 7939
rect 4813 7905 4847 7939
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 6653 7905 6687 7939
rect 7297 7905 7331 7939
rect 8125 7905 8159 7939
rect 8401 7905 8435 7939
rect 9873 7905 9907 7939
rect 5825 7837 5859 7871
rect 6929 7837 6963 7871
rect 8585 7837 8619 7871
rect 1869 7769 1903 7803
rect 5549 7497 5583 7531
rect 6929 7429 6963 7463
rect 2605 7361 2639 7395
rect 3157 7361 3191 7395
rect 7481 7361 7515 7395
rect 2513 7293 2547 7327
rect 2789 7293 2823 7327
rect 4169 7293 4203 7327
rect 4445 7293 4479 7327
rect 7403 7293 7437 7327
rect 7849 7293 7883 7327
rect 7941 7293 7975 7327
rect 8861 7293 8895 7327
rect 8953 7293 8987 7327
rect 9137 7293 9171 7327
rect 9321 7157 9355 7191
rect 2421 6817 2455 6851
rect 2881 6817 2915 6851
rect 3157 6817 3191 6851
rect 4353 6817 4387 6851
rect 4813 6817 4847 6851
rect 6101 6817 6135 6851
rect 6285 6817 6319 6851
rect 6469 6817 6503 6851
rect 6837 6817 6871 6851
rect 7021 6817 7055 6851
rect 8033 6817 8067 6851
rect 9873 6817 9907 6851
rect 5641 6749 5675 6783
rect 7941 6749 7975 6783
rect 10149 6749 10183 6783
rect 2237 6409 2271 6443
rect 2421 6409 2455 6443
rect 4077 6273 4111 6307
rect 5917 6273 5951 6307
rect 8769 6273 8803 6307
rect 3433 6205 3467 6239
rect 5457 6205 5491 6239
rect 5733 6205 5767 6239
rect 6929 6205 6963 6239
rect 9229 6205 9263 6239
rect 9413 6205 9447 6239
rect 9781 6205 9815 6239
rect 9965 6205 9999 6239
rect 2053 6137 2087 6171
rect 4905 6137 4939 6171
rect 7573 6137 7607 6171
rect 2237 6069 2271 6103
rect 1869 5865 1903 5899
rect 2789 5797 2823 5831
rect 1685 5729 1719 5763
rect 1869 5729 1903 5763
rect 2973 5729 3007 5763
rect 7021 5729 7055 5763
rect 8125 5729 8159 5763
rect 8309 5729 8343 5763
rect 8769 5729 8803 5763
rect 9873 5729 9907 5763
rect 4077 5661 4111 5695
rect 4353 5661 4387 5695
rect 8401 5661 8435 5695
rect 3065 5525 3099 5559
rect 5641 5525 5675 5559
rect 7021 5525 7055 5559
rect 9965 5525 9999 5559
rect 7113 5321 7147 5355
rect 10241 5321 10275 5355
rect 2881 5185 2915 5219
rect 2605 5117 2639 5151
rect 2697 5117 2731 5151
rect 3893 5117 3927 5151
rect 5181 5117 5215 5151
rect 6929 5117 6963 5151
rect 8585 5117 8619 5151
rect 10149 5117 10183 5151
rect 3709 5049 3743 5083
rect 4261 5049 4295 5083
rect 5733 5049 5767 5083
rect 8401 5049 8435 5083
rect 9965 5049 9999 5083
rect 8677 4981 8711 5015
rect 7481 4777 7515 4811
rect 1777 4709 1811 4743
rect 1961 4709 1995 4743
rect 6285 4709 6319 4743
rect 10057 4709 10091 4743
rect 1593 4641 1627 4675
rect 2881 4641 2915 4675
rect 3065 4641 3099 4675
rect 4721 4641 4755 4675
rect 4905 4641 4939 4675
rect 5917 4641 5951 4675
rect 7389 4641 7423 4675
rect 7665 4641 7699 4675
rect 7849 4641 7883 4675
rect 9689 4641 9723 4675
rect 9873 4641 9907 4675
rect 3157 4573 3191 4607
rect 4905 4505 4939 4539
rect 3433 4097 3467 4131
rect 5457 4097 5491 4131
rect 8769 4097 8803 4131
rect 1409 4029 1443 4063
rect 3065 4029 3099 4063
rect 3249 4029 3283 4063
rect 4353 4029 4387 4063
rect 4537 4029 4571 4063
rect 5641 4029 5675 4063
rect 6837 4029 6871 4063
rect 7389 4029 7423 4063
rect 9781 4029 9815 4063
rect 9873 4029 9907 4063
rect 4629 3961 4663 3995
rect 8401 3961 8435 3995
rect 8585 3961 8619 3995
rect 10057 3961 10091 3995
rect 1593 3893 1627 3927
rect 5825 3893 5859 3927
rect 7113 3893 7147 3927
rect 5181 3689 5215 3723
rect 6653 3689 6687 3723
rect 2329 3553 2363 3587
rect 4077 3553 4111 3587
rect 5181 3553 5215 3587
rect 5365 3553 5399 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 8217 3553 8251 3587
rect 8493 3553 8527 3587
rect 9781 3553 9815 3587
rect 9873 3553 9907 3587
rect 10057 3553 10091 3587
rect 8585 3485 8619 3519
rect 4261 3417 4295 3451
rect 2513 3349 2547 3383
rect 6285 3349 6319 3383
rect 4445 3145 4479 3179
rect 8401 3145 8435 3179
rect 10241 3145 10275 3179
rect 5825 3077 5859 3111
rect 7205 3077 7239 3111
rect 8861 3009 8895 3043
rect 3249 2941 3283 2975
rect 4445 2941 4479 2975
rect 4629 2941 4663 2975
rect 5549 2941 5583 2975
rect 5733 2941 5767 2975
rect 8769 2941 8803 2975
rect 9137 2941 9171 2975
rect 9321 2941 9355 2975
rect 10149 2941 10183 2975
rect 10425 2941 10459 2975
rect 6837 2873 6871 2907
rect 7021 2873 7055 2907
rect 3433 2805 3467 2839
rect 4721 2601 4755 2635
rect 8861 2533 8895 2567
rect 9965 2533 9999 2567
rect 10149 2533 10183 2567
rect 2881 2465 2915 2499
rect 4537 2465 4571 2499
rect 4721 2465 4755 2499
rect 5641 2465 5675 2499
rect 5825 2465 5859 2499
rect 7021 2465 7055 2499
rect 7205 2465 7239 2499
rect 7297 2465 7331 2499
rect 8769 2465 8803 2499
rect 9781 2465 9815 2499
rect 5917 2329 5951 2363
rect 3065 2261 3099 2295
<< metal1 >>
rect 1104 12538 11592 12560
rect 1104 12486 4478 12538
rect 4530 12486 4542 12538
rect 4594 12486 4606 12538
rect 4658 12486 4670 12538
rect 4722 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 11592 12538
rect 1104 12464 11592 12486
rect 5626 12316 5632 12368
rect 5684 12356 5690 12368
rect 5684 12328 8524 12356
rect 5684 12316 5690 12328
rect 4338 12288 4344 12300
rect 4299 12260 4344 12288
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4540 12220 4568 12251
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 4948 12260 5733 12288
rect 4948 12248 4954 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 7561 12291 7619 12297
rect 5960 12260 7144 12288
rect 5960 12248 5966 12260
rect 4304 12192 4568 12220
rect 5537 12223 5595 12229
rect 4304 12180 4310 12192
rect 5537 12189 5549 12223
rect 5583 12220 5595 12223
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 5583 12192 6929 12220
rect 5583 12189 5595 12192
rect 5537 12183 5595 12189
rect 6917 12189 6929 12192
rect 6963 12220 6975 12223
rect 7006 12220 7012 12232
rect 6963 12192 7012 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7116 12220 7144 12260
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 7742 12288 7748 12300
rect 7607 12260 7748 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 8496 12297 8524 12328
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12257 8539 12291
rect 8481 12251 8539 12257
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10686 12288 10692 12300
rect 10275 12260 10692 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 8680 12220 8708 12251
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 7116 12192 8708 12220
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4617 12155 4675 12161
rect 4617 12152 4629 12155
rect 4212 12124 4629 12152
rect 4212 12112 4218 12124
rect 4617 12121 4629 12124
rect 4663 12152 4675 12155
rect 4663 12124 7236 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 7098 12084 7104 12096
rect 5951 12056 7104 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7208 12084 7236 12124
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 8757 12155 8815 12161
rect 8757 12152 8769 12155
rect 7616 12124 8769 12152
rect 7616 12112 7622 12124
rect 8757 12121 8769 12124
rect 8803 12121 8815 12155
rect 8757 12115 8815 12121
rect 7742 12084 7748 12096
rect 7208 12056 7748 12084
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 9640 12056 10425 12084
rect 9640 12044 9646 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10413 12047 10471 12053
rect 1104 11994 11592 12016
rect 1104 11942 2730 11994
rect 2782 11942 2794 11994
rect 2846 11942 2858 11994
rect 2910 11942 2922 11994
rect 2974 11942 6226 11994
rect 6278 11942 6290 11994
rect 6342 11942 6354 11994
rect 6406 11942 6418 11994
rect 6470 11942 9722 11994
rect 9774 11942 9786 11994
rect 9838 11942 9850 11994
rect 9902 11942 9914 11994
rect 9966 11942 11592 11994
rect 1104 11920 11592 11942
rect 6914 11880 6920 11892
rect 5736 11852 6920 11880
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 4062 11744 4068 11756
rect 2096 11716 4068 11744
rect 2096 11704 2102 11716
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3510 11676 3516 11688
rect 3467 11648 3516 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3252 11608 3280 11639
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 4338 11676 4344 11688
rect 3936 11648 4344 11676
rect 3936 11636 3942 11648
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 5074 11676 5080 11688
rect 4755 11648 5080 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 3694 11608 3700 11620
rect 3252 11580 3700 11608
rect 3694 11568 3700 11580
rect 3752 11568 3758 11620
rect 4632 11608 4660 11639
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 5736 11676 5764 11852
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7466 11812 7472 11824
rect 5828 11784 7472 11812
rect 5828 11685 5856 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6604 11716 6837 11744
rect 6604 11704 6610 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 9766 11744 9772 11756
rect 6825 11707 6883 11713
rect 6932 11716 9772 11744
rect 5675 11648 5764 11676
rect 5813 11679 5871 11685
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 5813 11645 5825 11679
rect 5859 11645 5871 11679
rect 5813 11639 5871 11645
rect 6932 11608 6960 11716
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 4632 11580 6960 11608
rect 7024 11552 7052 11639
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 8297 11679 8355 11685
rect 8297 11676 8309 11679
rect 7156 11648 8309 11676
rect 7156 11636 7162 11648
rect 8297 11645 8309 11648
rect 8343 11645 8355 11679
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 8297 11639 8355 11645
rect 8588 11648 9321 11676
rect 7834 11568 7840 11620
rect 7892 11608 7898 11620
rect 8113 11611 8171 11617
rect 8113 11608 8125 11611
rect 7892 11580 8125 11608
rect 7892 11568 7898 11580
rect 8113 11577 8125 11580
rect 8159 11577 8171 11611
rect 8478 11608 8484 11620
rect 8439 11580 8484 11608
rect 8113 11571 8171 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 3234 11540 3240 11552
rect 3195 11512 3240 11540
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 4948 11512 5641 11540
rect 4948 11500 4954 11512
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 7006 11500 7012 11552
rect 7064 11500 7070 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 7156 11512 7205 11540
rect 7156 11500 7162 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 7193 11503 7251 11509
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 8588 11540 8616 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9508 11608 9536 11639
rect 8996 11580 9536 11608
rect 8996 11568 9002 11580
rect 7800 11512 8616 11540
rect 7800 11500 7806 11512
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 8720 11512 9413 11540
rect 8720 11500 8726 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 1104 11450 11592 11472
rect 1104 11398 4478 11450
rect 4530 11398 4542 11450
rect 4594 11398 4606 11450
rect 4658 11398 4670 11450
rect 4722 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 11592 11450
rect 1104 11376 11592 11398
rect 4338 11336 4344 11348
rect 3160 11308 4344 11336
rect 3160 11277 3188 11308
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 9766 11336 9772 11348
rect 9727 11308 9772 11336
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 3145 11271 3203 11277
rect 3145 11237 3157 11271
rect 3191 11237 3203 11271
rect 3145 11231 3203 11237
rect 5074 11228 5080 11280
rect 5132 11268 5138 11280
rect 5132 11240 9720 11268
rect 5132 11228 5138 11240
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11169 2927 11203
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 2869 11163 2927 11169
rect 2884 11132 2912 11163
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 3476 11172 4353 11200
rect 3476 11160 3482 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 9692 11209 9720 11240
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 7064 11172 7297 11200
rect 7064 11160 7070 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 9677 11203 9735 11209
rect 7699 11172 8800 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 3142 11132 3148 11144
rect 2884 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 4062 11132 4068 11144
rect 4023 11104 4068 11132
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6730 11132 6736 11144
rect 5767 11104 6736 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11132 7803 11135
rect 8386 11132 8392 11144
rect 7791 11104 8392 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 5552 11036 6132 11064
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 5552 10996 5580 11036
rect 3936 10968 5580 10996
rect 6104 10996 6132 11036
rect 8772 11008 8800 11172
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10042 11200 10048 11212
rect 9999 11172 10048 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 8570 10996 8576 11008
rect 6104 10968 8576 10996
rect 3936 10956 3942 10968
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8754 10996 8760 11008
rect 8667 10968 8760 10996
rect 8754 10956 8760 10968
rect 8812 10996 8818 11008
rect 10594 10996 10600 11008
rect 8812 10968 10600 10996
rect 8812 10956 8818 10968
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 1104 10906 11592 10928
rect 1104 10854 2730 10906
rect 2782 10854 2794 10906
rect 2846 10854 2858 10906
rect 2910 10854 2922 10906
rect 2974 10854 6226 10906
rect 6278 10854 6290 10906
rect 6342 10854 6354 10906
rect 6406 10854 6418 10906
rect 6470 10854 9722 10906
rect 9774 10854 9786 10906
rect 9838 10854 9850 10906
rect 9902 10854 9914 10906
rect 9966 10854 11592 10906
rect 1104 10832 11592 10854
rect 4154 10792 4160 10804
rect 2792 10764 4160 10792
rect 2792 10736 2820 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7524 10764 8125 10792
rect 7524 10752 7530 10764
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8113 10755 8171 10761
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 9214 10792 9220 10804
rect 8628 10764 9220 10792
rect 8628 10752 8634 10764
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 2774 10684 2780 10736
rect 2832 10684 2838 10736
rect 6914 10724 6920 10736
rect 3252 10696 6920 10724
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 3050 10656 3056 10668
rect 2271 10628 3056 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 1854 10588 1860 10600
rect 1815 10560 1860 10588
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2590 10588 2596 10600
rect 2179 10560 2596 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3252 10597 3280 10696
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 10318 10724 10324 10736
rect 8128 10696 10324 10724
rect 3513 10659 3571 10665
rect 3513 10625 3525 10659
rect 3559 10656 3571 10659
rect 7926 10656 7932 10668
rect 3559 10628 7932 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10588 3479 10591
rect 3602 10588 3608 10600
rect 3467 10560 3608 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4430 10588 4436 10600
rect 4391 10560 4436 10588
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10557 4583 10591
rect 5626 10588 5632 10600
rect 5587 10560 5632 10588
rect 4525 10551 4583 10557
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 4540 10520 4568 10551
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 7098 10588 7104 10600
rect 5859 10560 7104 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 8128 10597 8156 10696
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 10042 10656 10048 10668
rect 8352 10628 10048 10656
rect 8352 10616 8358 10628
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10557 8171 10591
rect 8113 10551 8171 10557
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 8386 10588 8392 10600
rect 8251 10560 8392 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 8386 10548 8392 10560
rect 8444 10588 8450 10600
rect 9214 10588 9220 10600
rect 8444 10560 9076 10588
rect 9175 10560 9220 10588
rect 8444 10548 8450 10560
rect 4212 10492 4568 10520
rect 4709 10523 4767 10529
rect 4212 10480 4218 10492
rect 4709 10489 4721 10523
rect 4755 10520 4767 10523
rect 5902 10520 5908 10532
rect 4755 10492 5908 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4724 10452 4752 10483
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 6825 10523 6883 10529
rect 6825 10520 6837 10523
rect 6788 10492 6837 10520
rect 6788 10480 6794 10492
rect 6825 10489 6837 10492
rect 6871 10489 6883 10523
rect 7006 10520 7012 10532
rect 6967 10492 7012 10520
rect 6825 10483 6883 10489
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7193 10523 7251 10529
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 8294 10520 8300 10532
rect 7239 10492 8300 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 9048 10520 9076 10560
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9398 10588 9404 10600
rect 9359 10560 9404 10588
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 10502 10520 10508 10532
rect 9048 10492 10508 10520
rect 10502 10480 10508 10492
rect 10560 10520 10566 10532
rect 11974 10520 11980 10532
rect 10560 10492 11980 10520
rect 10560 10480 10566 10492
rect 11974 10480 11980 10492
rect 12032 10480 12038 10532
rect 4120 10424 4752 10452
rect 4120 10412 4126 10424
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5132 10424 5641 10452
rect 5132 10412 5138 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 6052 10424 9321 10452
rect 6052 10412 6058 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 9309 10415 9367 10421
rect 1104 10362 11592 10384
rect 1104 10310 4478 10362
rect 4530 10310 4542 10362
rect 4594 10310 4606 10362
rect 4658 10310 4670 10362
rect 4722 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 11592 10362
rect 1104 10288 11592 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 4246 10248 4252 10260
rect 1903 10220 4252 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 5776 10220 6193 10248
rect 5776 10208 5782 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 7466 10248 7472 10260
rect 7427 10220 7472 10248
rect 6181 10211 6239 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 9306 10248 9312 10260
rect 8803 10220 9312 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 4890 10180 4896 10192
rect 3068 10152 4896 10180
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10081 1731 10115
rect 1673 10075 1731 10081
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 2958 10112 2964 10124
rect 2915 10084 2964 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 1688 9976 1716 10075
rect 1872 10044 1900 10075
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3068 10121 3096 10152
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 5169 10183 5227 10189
rect 5169 10149 5181 10183
rect 5215 10180 5227 10183
rect 5626 10180 5632 10192
rect 5215 10152 5632 10180
rect 5215 10149 5227 10152
rect 5169 10143 5227 10149
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 5997 10183 6055 10189
rect 5997 10149 6009 10183
rect 6043 10149 6055 10183
rect 5997 10143 6055 10149
rect 7285 10183 7343 10189
rect 7285 10149 7297 10183
rect 7331 10149 7343 10183
rect 7285 10143 7343 10149
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10081 3111 10115
rect 4798 10112 4804 10124
rect 4759 10084 4804 10112
rect 3053 10075 3111 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5258 10072 5264 10124
rect 5316 10112 5322 10124
rect 6012 10112 6040 10143
rect 5316 10084 6040 10112
rect 7300 10112 7328 10143
rect 7466 10112 7472 10124
rect 7300 10084 7472 10112
rect 5316 10072 5322 10084
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 7708 10084 7757 10112
rect 7708 10072 7714 10084
rect 7745 10081 7757 10084
rect 7791 10081 7803 10115
rect 8570 10112 8576 10124
rect 8531 10084 8576 10112
rect 7745 10075 7803 10081
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9364 10084 9689 10112
rect 9364 10072 9370 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10112 10011 10115
rect 10134 10112 10140 10124
rect 9999 10084 10140 10112
rect 9999 10081 10011 10084
rect 9953 10075 10011 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 2774 10044 2780 10056
rect 1872 10016 2780 10044
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 9398 10044 9404 10056
rect 3191 10016 9404 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10594 10044 10600 10056
rect 10091 10016 10600 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 4246 9976 4252 9988
rect 1688 9948 4252 9976
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 6365 9979 6423 9985
rect 6365 9945 6377 9979
rect 6411 9976 6423 9979
rect 6411 9948 9444 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 9416 9920 9444 9948
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 5994 9908 6000 9920
rect 3108 9880 6000 9908
rect 3108 9868 3114 9880
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 6144 9880 6193 9908
rect 6144 9868 6150 9880
rect 6181 9877 6193 9880
rect 6227 9877 6239 9911
rect 6181 9871 6239 9877
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 8386 9908 8392 9920
rect 7515 9880 8392 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9398 9868 9404 9920
rect 9456 9868 9462 9920
rect 1104 9818 11592 9840
rect 1104 9766 2730 9818
rect 2782 9766 2794 9818
rect 2846 9766 2858 9818
rect 2910 9766 2922 9818
rect 2974 9766 6226 9818
rect 6278 9766 6290 9818
rect 6342 9766 6354 9818
rect 6406 9766 6418 9818
rect 6470 9766 9722 9818
rect 9774 9766 9786 9818
rect 9838 9766 9850 9818
rect 9902 9766 9914 9818
rect 9966 9766 11592 9818
rect 1104 9744 11592 9766
rect 658 9664 664 9716
rect 716 9704 722 9716
rect 2498 9704 2504 9716
rect 716 9676 2504 9704
rect 716 9664 722 9676
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 8386 9704 8392 9716
rect 3660 9676 8392 9704
rect 3660 9664 3666 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 8757 9707 8815 9713
rect 8757 9704 8769 9707
rect 8628 9676 8769 9704
rect 8628 9664 8634 9676
rect 8757 9673 8769 9676
rect 8803 9673 8815 9707
rect 8757 9667 8815 9673
rect 9122 9664 9128 9716
rect 9180 9704 9186 9716
rect 10042 9704 10048 9716
rect 9180 9676 10048 9704
rect 9180 9664 9186 9676
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 5074 9636 5080 9648
rect 4356 9608 5080 9636
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 3510 9568 3516 9580
rect 2363 9540 3516 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9500 2559 9503
rect 2590 9500 2596 9512
rect 2547 9472 2596 9500
rect 2547 9469 2559 9472
rect 2501 9463 2559 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 4356 9509 4384 9608
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 7282 9636 7288 9648
rect 5684 9608 6960 9636
rect 7243 9608 7288 9636
rect 5684 9596 5690 9608
rect 6638 9568 6644 9580
rect 4540 9540 6644 9568
rect 4540 9509 4568 9540
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9469 4583 9503
rect 5442 9500 5448 9512
rect 5403 9472 5448 9500
rect 4525 9463 4583 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 6932 9509 6960 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5592 9472 5641 9500
rect 5592 9460 5598 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9469 6975 9503
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 6917 9463 6975 9469
rect 7024 9472 8401 9500
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 7024 9432 7052 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 10410 9500 10416 9512
rect 8619 9472 10416 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 2004 9404 7052 9432
rect 2004 9392 2010 9404
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 9456 9404 9689 9432
rect 9456 9392 9462 9404
rect 9677 9401 9689 9404
rect 9723 9401 9735 9435
rect 9677 9395 9735 9401
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9401 9919 9435
rect 10042 9432 10048 9444
rect 9955 9404 10048 9432
rect 9861 9395 9919 9401
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 2685 9367 2743 9373
rect 2685 9364 2697 9367
rect 1636 9336 2697 9364
rect 1636 9324 1642 9336
rect 2685 9333 2697 9336
rect 2731 9364 2743 9367
rect 3418 9364 3424 9376
rect 2731 9336 3424 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 4338 9364 4344 9376
rect 4299 9336 4344 9364
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 9876 9364 9904 9395
rect 10042 9392 10048 9404
rect 10100 9432 10106 9444
rect 10870 9432 10876 9444
rect 10100 9404 10876 9432
rect 10100 9392 10106 9404
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10226 9364 10232 9376
rect 7432 9336 10232 9364
rect 7432 9324 7438 9336
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 1104 9274 11592 9296
rect 1104 9222 4478 9274
rect 4530 9222 4542 9274
rect 4594 9222 4606 9274
rect 4658 9222 4670 9274
rect 4722 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 11592 9274
rect 1104 9200 11592 9222
rect 6546 9160 6552 9172
rect 4540 9132 6552 9160
rect 1578 9092 1584 9104
rect 1539 9064 1584 9092
rect 1578 9052 1584 9064
rect 1636 9052 1642 9104
rect 1946 9092 1952 9104
rect 1907 9064 1952 9092
rect 1946 9052 1952 9064
rect 2004 9052 2010 9104
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 4154 9092 4160 9104
rect 3191 9064 4160 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 4540 9036 4568 9132
rect 6546 9120 6552 9132
rect 6604 9160 6610 9172
rect 8938 9160 8944 9172
rect 6604 9132 8944 9160
rect 6604 9120 6610 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5132 9064 7696 9092
rect 5132 9052 5138 9064
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 8993 1823 9027
rect 2866 9024 2872 9036
rect 2827 8996 2872 9024
rect 1765 8987 1823 8993
rect 1780 8888 1808 8987
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 8993 3111 9027
rect 3053 8987 3111 8993
rect 3068 8956 3096 8987
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 4522 9024 4528 9036
rect 3752 8996 4528 9024
rect 3752 8984 3758 8996
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 4614 8984 4620 9036
rect 4672 9033 4678 9036
rect 4672 9024 4679 9033
rect 6546 9024 6552 9036
rect 4672 8996 4717 9024
rect 6507 8996 6552 9024
rect 4672 8987 4679 8996
rect 4672 8984 4678 8987
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7668 9033 7696 9064
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 6972 8996 7573 9024
rect 6972 8984 6978 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 7800 8996 9689 9024
rect 7800 8984 7806 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 4062 8956 4068 8968
rect 3068 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4430 8956 4436 8968
rect 4391 8928 4436 8956
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5626 8888 5632 8900
rect 1780 8860 5632 8888
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 5736 8888 5764 8919
rect 5994 8916 6000 8968
rect 6052 8956 6058 8968
rect 6273 8959 6331 8965
rect 6273 8956 6285 8959
rect 6052 8928 6285 8956
rect 6052 8916 6058 8928
rect 6273 8925 6285 8928
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7190 8956 7196 8968
rect 6779 8928 7196 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7190 8916 7196 8928
rect 7248 8956 7254 8968
rect 7834 8956 7840 8968
rect 7248 8928 7840 8956
rect 7248 8916 7254 8928
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 9876 8956 9904 8987
rect 8076 8928 9904 8956
rect 8076 8916 8082 8928
rect 10042 8888 10048 8900
rect 5736 8860 10048 8888
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 4338 8820 4344 8832
rect 1728 8792 4344 8820
rect 1728 8780 1734 8792
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5644 8820 5672 8848
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 5644 8792 9781 8820
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 1104 8730 11592 8752
rect 1104 8678 2730 8730
rect 2782 8678 2794 8730
rect 2846 8678 2858 8730
rect 2910 8678 2922 8730
rect 2974 8678 6226 8730
rect 6278 8678 6290 8730
rect 6342 8678 6354 8730
rect 6406 8678 6418 8730
rect 6470 8678 9722 8730
rect 9774 8678 9786 8730
rect 9838 8678 9850 8730
rect 9902 8678 9914 8730
rect 9966 8678 11592 8730
rect 1104 8656 11592 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 2372 8588 3433 8616
rect 2372 8576 2378 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 4856 8588 10057 8616
rect 4856 8576 4862 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10045 8579 10103 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 3789 8551 3847 8557
rect 3789 8548 3801 8551
rect 3660 8520 3801 8548
rect 3660 8508 3666 8520
rect 3789 8517 3801 8520
rect 3835 8548 3847 8551
rect 3878 8548 3884 8560
rect 3835 8520 3884 8548
rect 3835 8517 3847 8520
rect 3789 8511 3847 8517
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4430 8548 4436 8560
rect 4120 8520 4436 8548
rect 4120 8508 4126 8520
rect 4430 8508 4436 8520
rect 4488 8548 4494 8560
rect 4982 8548 4988 8560
rect 4488 8520 4988 8548
rect 4488 8508 4494 8520
rect 4982 8508 4988 8520
rect 5040 8548 5046 8560
rect 5040 8520 6592 8548
rect 5040 8508 5046 8520
rect 6564 8492 6592 8520
rect 7098 8508 7104 8560
rect 7156 8548 7162 8560
rect 7834 8548 7840 8560
rect 7156 8520 7840 8548
rect 7156 8508 7162 8520
rect 2498 8440 2504 8492
rect 2556 8480 2562 8492
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 2556 8452 3525 8480
rect 2556 8440 2562 8452
rect 3513 8449 3525 8452
rect 3559 8480 3571 8483
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 3559 8452 5273 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 7190 8480 7196 8492
rect 6656 8452 7196 8480
rect 1486 8412 1492 8424
rect 1447 8384 1492 8412
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 4154 8412 4160 8424
rect 3467 8384 4160 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 5353 8415 5411 8421
rect 5353 8381 5365 8415
rect 5399 8412 5411 8415
rect 5399 8384 5672 8412
rect 5399 8381 5411 8384
rect 5353 8375 5411 8381
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 2590 8344 2596 8356
rect 2179 8316 2596 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 2590 8304 2596 8316
rect 2648 8304 2654 8356
rect 4709 8347 4767 8353
rect 4709 8313 4721 8347
rect 4755 8344 4767 8347
rect 4890 8344 4896 8356
rect 4755 8316 4896 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 4798 8276 4804 8288
rect 2832 8248 4804 8276
rect 2832 8236 2838 8248
rect 4798 8236 4804 8248
rect 4856 8276 4862 8288
rect 5074 8276 5080 8288
rect 4856 8248 5080 8276
rect 4856 8236 4862 8248
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5644 8276 5672 8384
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 5905 8415 5963 8421
rect 5776 8384 5821 8412
rect 5776 8372 5782 8384
rect 5905 8381 5917 8415
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 5920 8344 5948 8375
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 6656 8412 6684 8452
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 6822 8412 6828 8424
rect 6512 8384 6684 8412
rect 6783 8384 6828 8412
rect 6512 8372 6518 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7098 8412 7104 8424
rect 7059 8384 7104 8412
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7300 8421 7328 8520
rect 7834 8508 7840 8520
rect 7892 8508 7898 8560
rect 8481 8551 8539 8557
rect 8481 8517 8493 8551
rect 8527 8548 8539 8551
rect 9306 8548 9312 8560
rect 8527 8520 9312 8548
rect 8527 8517 8539 8520
rect 8481 8511 8539 8517
rect 9306 8508 9312 8520
rect 9364 8508 9370 8560
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 9674 8548 9680 8560
rect 9456 8520 9680 8548
rect 9456 8508 9462 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 7432 8452 9229 8480
rect 7432 8440 7438 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10226 8480 10232 8492
rect 10183 8452 10232 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8381 7343 8415
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7285 8375 7343 8381
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 7668 8384 8769 8412
rect 6086 8344 6092 8356
rect 5920 8316 6092 8344
rect 6086 8304 6092 8316
rect 6144 8344 6150 8356
rect 6144 8316 7144 8344
rect 6144 8304 6150 8316
rect 6917 8279 6975 8285
rect 6917 8276 6929 8279
rect 5644 8248 6929 8276
rect 6917 8245 6929 8248
rect 6963 8245 6975 8279
rect 7116 8276 7144 8316
rect 7190 8304 7196 8356
rect 7248 8344 7254 8356
rect 7668 8344 7696 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 10042 8412 10048 8424
rect 10003 8384 10048 8412
rect 8757 8375 8815 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 8018 8344 8024 8356
rect 7248 8316 7696 8344
rect 7760 8316 8024 8344
rect 7248 8304 7254 8316
rect 7558 8276 7564 8288
rect 7116 8248 7564 8276
rect 6917 8239 6975 8245
rect 7558 8236 7564 8248
rect 7616 8276 7622 8288
rect 7760 8276 7788 8316
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8665 8347 8723 8353
rect 8665 8313 8677 8347
rect 8711 8344 8723 8347
rect 8846 8344 8852 8356
rect 8711 8316 8852 8344
rect 8711 8313 8723 8316
rect 8665 8307 8723 8313
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 7616 8248 7788 8276
rect 7616 8236 7622 8248
rect 1104 8186 11592 8208
rect 1104 8134 4478 8186
rect 4530 8134 4542 8186
rect 4594 8134 4606 8186
rect 4658 8134 4670 8186
rect 4722 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 11592 8186
rect 1104 8112 11592 8134
rect 4062 8072 4068 8084
rect 2976 8044 4068 8072
rect 2976 8013 3004 8044
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4212 8044 4261 8072
rect 4212 8032 4218 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 6178 8072 6184 8084
rect 4249 8035 4307 8041
rect 4356 8044 6184 8072
rect 2961 8007 3019 8013
rect 2961 7973 2973 8007
rect 3007 7973 3019 8007
rect 2961 7967 3019 7973
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7905 1915 7939
rect 1857 7899 1915 7905
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 2866 7936 2872 7948
rect 2823 7908 2872 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 1872 7868 1900 7899
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 4062 7936 4068 7948
rect 3191 7908 4068 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4246 7936 4252 7948
rect 4159 7908 4252 7936
rect 4246 7896 4252 7908
rect 4304 7936 4310 7948
rect 4356 7936 4384 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 6696 8044 8401 8072
rect 6696 8032 6702 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 4724 7976 6776 8004
rect 4304 7908 4384 7936
rect 4433 7939 4491 7945
rect 4304 7896 4310 7908
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4614 7936 4620 7948
rect 4479 7908 4620 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4724 7945 4752 7976
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 1872 7840 3372 7868
rect 1857 7803 1915 7809
rect 1857 7769 1869 7803
rect 1903 7800 1915 7803
rect 2774 7800 2780 7812
rect 1903 7772 2780 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 2774 7760 2780 7772
rect 2832 7760 2838 7812
rect 3344 7732 3372 7840
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 4816 7868 4844 7899
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 5684 7908 6285 7936
rect 5684 7896 5690 7908
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 6454 7936 6460 7948
rect 6415 7908 6460 7936
rect 6273 7899 6331 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6604 7908 6653 7936
rect 6604 7896 6610 7908
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6748 7936 6776 7976
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 9677 8007 9735 8013
rect 9677 8004 9689 8007
rect 7064 7976 9689 8004
rect 7064 7964 7070 7976
rect 9677 7973 9689 7976
rect 9723 7973 9735 8007
rect 9677 7967 9735 7973
rect 10229 8007 10287 8013
rect 10229 7973 10241 8007
rect 10275 8004 10287 8007
rect 10686 8004 10692 8016
rect 10275 7976 10692 8004
rect 10275 7973 10287 7976
rect 10229 7967 10287 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 7282 7936 7288 7948
rect 6748 7908 7052 7936
rect 7243 7908 7288 7936
rect 6641 7899 6699 7905
rect 3476 7840 4844 7868
rect 5813 7871 5871 7877
rect 3476 7828 3482 7840
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5902 7868 5908 7880
rect 5859 7840 5908 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6236 7840 6929 7868
rect 6236 7828 6242 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 7024 7868 7052 7908
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 8110 7936 8116 7948
rect 8071 7908 8116 7936
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8938 7936 8944 7948
rect 8435 7908 8944 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 10410 7936 10416 7948
rect 9907 7908 10416 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 8478 7868 8484 7880
rect 7024 7840 8484 7868
rect 6917 7831 6975 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 4246 7760 4252 7812
rect 4304 7800 4310 7812
rect 7466 7800 7472 7812
rect 4304 7772 7472 7800
rect 4304 7760 4310 7772
rect 7466 7760 7472 7772
rect 7524 7800 7530 7812
rect 8588 7800 8616 7831
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9876 7868 9904 7899
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 9732 7840 9904 7868
rect 9732 7828 9738 7840
rect 7524 7772 8616 7800
rect 7524 7760 7530 7772
rect 7650 7732 7656 7744
rect 3344 7704 7656 7732
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 1104 7642 11592 7664
rect 1104 7590 2730 7642
rect 2782 7590 2794 7642
rect 2846 7590 2858 7642
rect 2910 7590 2922 7642
rect 2974 7590 6226 7642
rect 6278 7590 6290 7642
rect 6342 7590 6354 7642
rect 6406 7590 6418 7642
rect 6470 7590 9722 7642
rect 9774 7590 9786 7642
rect 9838 7590 9850 7642
rect 9902 7590 9914 7642
rect 9966 7590 11592 7642
rect 1104 7568 11592 7590
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 4396 7500 5549 7528
rect 4396 7488 4402 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 9490 7528 9496 7540
rect 5960 7500 9496 7528
rect 5960 7488 5966 7500
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 6917 7463 6975 7469
rect 6917 7429 6929 7463
rect 6963 7460 6975 7463
rect 7282 7460 7288 7472
rect 6963 7432 7288 7460
rect 6963 7429 6975 7432
rect 6917 7423 6975 7429
rect 7282 7420 7288 7432
rect 7340 7420 7346 7472
rect 7558 7460 7564 7472
rect 7484 7432 7564 7460
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2464 7364 2605 7392
rect 2464 7352 2470 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 2593 7355 2651 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 7484 7401 7512 7432
rect 7558 7420 7564 7432
rect 7616 7420 7622 7472
rect 10594 7460 10600 7472
rect 7852 7432 10600 7460
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2516 7256 2544 7287
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2740 7296 2789 7324
rect 2740 7284 2746 7296
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 2777 7287 2835 7293
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 4028 7296 4169 7324
rect 4028 7284 4034 7296
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4157 7287 4215 7293
rect 4264 7296 4445 7324
rect 3326 7256 3332 7268
rect 2516 7228 3332 7256
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 4264 7256 4292 7296
rect 4433 7293 4445 7296
rect 4479 7324 4491 7327
rect 5626 7324 5632 7336
rect 4479 7296 5632 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 7852 7333 7880 7432
rect 10594 7420 10600 7432
rect 10652 7420 10658 7472
rect 7391 7327 7449 7333
rect 7391 7324 7403 7327
rect 6604 7296 7403 7324
rect 6604 7284 6610 7296
rect 7391 7293 7403 7296
rect 7437 7293 7449 7327
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7391 7287 7449 7293
rect 7668 7296 7849 7324
rect 3844 7228 4292 7256
rect 3844 7216 3850 7228
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 7668 7256 7696 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 7944 7256 7972 7287
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8720 7296 8861 7324
rect 8720 7284 8726 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9122 7324 9128 7336
rect 8996 7296 9041 7324
rect 9083 7296 9128 7324
rect 8996 7284 9002 7296
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 7248 7228 7696 7256
rect 7760 7228 7972 7256
rect 7248 7216 7254 7228
rect 7760 7200 7788 7228
rect 7742 7148 7748 7200
rect 7800 7148 7806 7200
rect 9306 7188 9312 7200
rect 9267 7160 9312 7188
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 1104 7098 11592 7120
rect 1104 7046 4478 7098
rect 4530 7046 4542 7098
rect 4594 7046 4606 7098
rect 4658 7046 4670 7098
rect 4722 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 11592 7098
rect 1104 7024 11592 7046
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 8662 6984 8668 6996
rect 5408 6956 8668 6984
rect 5408 6944 5414 6956
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 4890 6916 4896 6928
rect 2424 6888 4896 6916
rect 2424 6857 2452 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2556 6820 2881 6848
rect 2556 6808 2562 6820
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 3108 6820 3157 6848
rect 3108 6808 3114 6820
rect 3145 6817 3157 6820
rect 3191 6848 3203 6851
rect 4338 6848 4344 6860
rect 3191 6820 3740 6848
rect 4299 6820 4344 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3712 6780 3740 6820
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 4764 6820 4813 6848
rect 4764 6808 4770 6820
rect 4801 6817 4813 6820
rect 4847 6848 4859 6851
rect 5074 6848 5080 6860
rect 4847 6820 5080 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5442 6848 5448 6860
rect 5184 6820 5448 6848
rect 5184 6780 5212 6820
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 5500 6820 5948 6848
rect 5500 6808 5506 6820
rect 3712 6752 5212 6780
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5920 6780 5948 6820
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 6052 6820 6101 6848
rect 6052 6808 6058 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6089 6811 6147 6817
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 6236 6820 6285 6848
rect 6236 6808 6242 6820
rect 6273 6817 6285 6820
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6817 6515 6851
rect 6822 6848 6828 6860
rect 6783 6820 6828 6848
rect 6457 6811 6515 6817
rect 6472 6780 6500 6811
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 7006 6848 7012 6860
rect 6967 6820 7012 6848
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7156 6820 8033 6848
rect 7156 6808 7162 6820
rect 8021 6817 8033 6820
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10226 6848 10232 6860
rect 9907 6820 10232 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 7024 6780 7052 6808
rect 5920 6752 6500 6780
rect 6840 6752 7052 6780
rect 5629 6743 5687 6749
rect 5644 6712 5672 6743
rect 6840 6724 6868 6752
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7708 6752 7941 6780
rect 7708 6740 7714 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 7929 6743 7987 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 5902 6712 5908 6724
rect 5644 6684 5908 6712
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 6822 6672 6828 6724
rect 6880 6672 6886 6724
rect 10686 6712 10692 6724
rect 6932 6684 10692 6712
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 6932 6644 6960 6684
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 2372 6616 6960 6644
rect 2372 6604 2378 6616
rect 1104 6554 11592 6576
rect 1104 6502 2730 6554
rect 2782 6502 2794 6554
rect 2846 6502 2858 6554
rect 2910 6502 2922 6554
rect 2974 6502 6226 6554
rect 6278 6502 6290 6554
rect 6342 6502 6354 6554
rect 6406 6502 6418 6554
rect 6470 6502 9722 6554
rect 9774 6502 9786 6554
rect 9838 6502 9850 6554
rect 9902 6502 9914 6554
rect 9966 6502 11592 6554
rect 1104 6480 11592 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6409 2283 6443
rect 2225 6403 2283 6409
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 8938 6440 8944 6452
rect 2455 6412 8944 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 2240 6372 2268 6403
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 3786 6372 3792 6384
rect 2240 6344 3792 6372
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 3988 6344 8800 6372
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 2464 6208 3433 6236
rect 2464 6196 2470 6208
rect 3421 6205 3433 6208
rect 3467 6236 3479 6239
rect 3988 6236 4016 6344
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 5350 6304 5356 6316
rect 4111 6276 5356 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 5592 6276 5917 6304
rect 5592 6264 5598 6276
rect 5905 6273 5917 6276
rect 5951 6304 5963 6307
rect 6822 6304 6828 6316
rect 5951 6276 6828 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 8772 6313 8800 6344
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 9858 6304 9864 6316
rect 8757 6267 8815 6273
rect 9416 6276 9864 6304
rect 3467 6208 4016 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 4212 6208 5457 6236
rect 4212 6196 4218 6208
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6270 6236 6276 6248
rect 5767 6208 6276 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6205 6975 6239
rect 9214 6236 9220 6248
rect 9175 6208 9220 6236
rect 6917 6199 6975 6205
rect 2041 6171 2099 6177
rect 2041 6137 2053 6171
rect 2087 6168 2099 6171
rect 4706 6168 4712 6180
rect 2087 6140 4712 6168
rect 2087 6137 2099 6140
rect 2041 6131 2099 6137
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 4893 6171 4951 6177
rect 4893 6137 4905 6171
rect 4939 6168 4951 6171
rect 6086 6168 6092 6180
rect 4939 6140 6092 6168
rect 4939 6137 4951 6140
rect 4893 6131 4951 6137
rect 6086 6128 6092 6140
rect 6144 6128 6150 6180
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 4798 6100 4804 6112
rect 2271 6072 4804 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6730 6100 6736 6112
rect 5592 6072 6736 6100
rect 5592 6060 5598 6072
rect 6730 6060 6736 6072
rect 6788 6100 6794 6112
rect 6932 6100 6960 6199
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9416 6245 9444 6276
rect 9858 6264 9864 6276
rect 9916 6304 9922 6316
rect 10134 6304 10140 6316
rect 9916 6276 10140 6304
rect 9916 6264 9922 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9548 6208 9781 6236
rect 9548 6196 9554 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10042 6236 10048 6248
rect 9999 6208 10048 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 7466 6128 7472 6180
rect 7524 6168 7530 6180
rect 7561 6171 7619 6177
rect 7561 6168 7573 6171
rect 7524 6140 7573 6168
rect 7524 6128 7530 6140
rect 7561 6137 7573 6140
rect 7607 6137 7619 6171
rect 7561 6131 7619 6137
rect 6788 6072 6960 6100
rect 6788 6060 6794 6072
rect 1104 6010 11592 6032
rect 1104 5958 4478 6010
rect 4530 5958 4542 6010
rect 4594 5958 4606 6010
rect 4658 5958 4670 6010
rect 4722 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 11592 6010
rect 1104 5936 11592 5958
rect 1857 5899 1915 5905
rect 1857 5865 1869 5899
rect 1903 5896 1915 5899
rect 2498 5896 2504 5908
rect 1903 5868 2504 5896
rect 1903 5865 1915 5868
rect 1857 5859 1915 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 7834 5896 7840 5908
rect 2792 5868 7840 5896
rect 1762 5828 1768 5840
rect 1675 5800 1768 5828
rect 1688 5769 1716 5800
rect 1762 5788 1768 5800
rect 1820 5828 1826 5840
rect 2792 5837 2820 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 2777 5831 2835 5837
rect 1820 5800 1992 5828
rect 1820 5788 1826 5800
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 1964 5760 1992 5800
rect 2777 5797 2789 5831
rect 2823 5797 2835 5831
rect 3050 5828 3056 5840
rect 2777 5791 2835 5797
rect 2884 5800 3056 5828
rect 2884 5760 2912 5800
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 1964 5732 2912 5760
rect 2961 5763 3019 5769
rect 1857 5723 1915 5729
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 5994 5760 6000 5772
rect 3007 5732 6000 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 1872 5692 1900 5723
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 7006 5760 7012 5772
rect 6696 5732 7012 5760
rect 6696 5720 6702 5732
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 8113 5763 8171 5769
rect 8113 5760 8125 5763
rect 7892 5732 8125 5760
rect 7892 5720 7898 5732
rect 8113 5729 8125 5732
rect 8159 5729 8171 5763
rect 8294 5760 8300 5772
rect 8255 5732 8300 5760
rect 8113 5723 8171 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8754 5760 8760 5772
rect 8715 5732 8760 5760
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9858 5760 9864 5772
rect 9819 5732 9864 5760
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 3050 5692 3056 5704
rect 1872 5664 3056 5692
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 4028 5664 4077 5692
rect 4028 5652 4034 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4065 5655 4123 5661
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 7190 5624 7196 5636
rect 6788 5596 7196 5624
rect 6788 5584 6794 5596
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5556 3111 5559
rect 5350 5556 5356 5568
rect 3099 5528 5356 5556
rect 3099 5525 3111 5528
rect 3053 5519 3111 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5500 5528 5641 5556
rect 5500 5516 5506 5528
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 5629 5519 5687 5525
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 7006 5556 7012 5568
rect 5776 5528 7012 5556
rect 5776 5516 5782 5528
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 9953 5559 10011 5565
rect 9953 5525 9965 5559
rect 9999 5556 10011 5559
rect 10042 5556 10048 5568
rect 9999 5528 10048 5556
rect 9999 5525 10011 5528
rect 9953 5519 10011 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 1104 5466 11592 5488
rect 1104 5414 2730 5466
rect 2782 5414 2794 5466
rect 2846 5414 2858 5466
rect 2910 5414 2922 5466
rect 2974 5414 6226 5466
rect 6278 5414 6290 5466
rect 6342 5414 6354 5466
rect 6406 5414 6418 5466
rect 6470 5414 9722 5466
rect 9774 5414 9786 5466
rect 9838 5414 9850 5466
rect 9902 5414 9914 5466
rect 9966 5414 11592 5466
rect 1104 5392 11592 5414
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 6972 5324 7113 5352
rect 6972 5312 6978 5324
rect 7101 5321 7113 5324
rect 7147 5352 7159 5355
rect 7190 5352 7196 5364
rect 7147 5324 7196 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 10226 5352 10232 5364
rect 10187 5324 10232 5352
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 7650 5284 7656 5296
rect 2700 5256 7656 5284
rect 2700 5216 2728 5256
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 2608 5188 2728 5216
rect 2869 5219 2927 5225
rect 2608 5157 2636 5188
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 3050 5216 3056 5228
rect 2915 5188 3056 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 9306 5216 9312 5228
rect 3344 5188 9312 5216
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 3344 5148 3372 5188
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 2731 5120 3372 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3476 5120 3893 5148
rect 3476 5108 3482 5120
rect 3881 5117 3893 5120
rect 3927 5148 3939 5151
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 3927 5120 5181 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 5169 5117 5181 5120
rect 5215 5148 5227 5151
rect 5442 5148 5448 5160
rect 5215 5120 5448 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6052 5120 6929 5148
rect 6052 5108 6058 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 8570 5148 8576 5160
rect 8531 5120 8576 5148
rect 6917 5111 6975 5117
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 10134 5148 10140 5160
rect 10095 5120 10140 5148
rect 10134 5108 10140 5120
rect 10192 5108 10198 5160
rect 3697 5083 3755 5089
rect 3697 5049 3709 5083
rect 3743 5049 3755 5083
rect 3697 5043 3755 5049
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5080 4307 5083
rect 5626 5080 5632 5092
rect 4295 5052 5632 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 3712 5012 3740 5043
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 5718 5040 5724 5092
rect 5776 5080 5782 5092
rect 6638 5080 6644 5092
rect 5776 5052 6644 5080
rect 5776 5040 5782 5052
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 7466 5040 7472 5092
rect 7524 5080 7530 5092
rect 8294 5080 8300 5092
rect 7524 5052 8300 5080
rect 7524 5040 7530 5052
rect 8294 5040 8300 5052
rect 8352 5080 8358 5092
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 8352 5052 8401 5080
rect 8352 5040 8358 5052
rect 8389 5049 8401 5052
rect 8435 5049 8447 5083
rect 8389 5043 8447 5049
rect 9953 5083 10011 5089
rect 9953 5049 9965 5083
rect 9999 5080 10011 5083
rect 10686 5080 10692 5092
rect 9999 5052 10692 5080
rect 9999 5049 10011 5052
rect 9953 5043 10011 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 7834 5012 7840 5024
rect 3712 4984 7840 5012
rect 7834 4972 7840 4984
rect 7892 5012 7898 5024
rect 8665 5015 8723 5021
rect 8665 5012 8677 5015
rect 7892 4984 8677 5012
rect 7892 4972 7898 4984
rect 8665 4981 8677 4984
rect 8711 4981 8723 5015
rect 8665 4975 8723 4981
rect 1104 4922 11592 4944
rect 1104 4870 4478 4922
rect 4530 4870 4542 4922
rect 4594 4870 4606 4922
rect 4658 4870 4670 4922
rect 4722 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 11592 4922
rect 1104 4848 11592 4870
rect 7466 4808 7472 4820
rect 1964 4780 7328 4808
rect 7427 4780 7472 4808
rect 1762 4740 1768 4752
rect 1723 4712 1768 4740
rect 1762 4700 1768 4712
rect 1820 4700 1826 4752
rect 1964 4749 1992 4780
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4709 2007 4743
rect 4154 4740 4160 4752
rect 1949 4703 2007 4709
rect 2884 4712 4160 4740
rect 2884 4681 2912 4712
rect 4154 4700 4160 4712
rect 4212 4740 4218 4752
rect 4982 4740 4988 4752
rect 4212 4712 4988 4740
rect 4212 4700 4218 4712
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 5718 4740 5724 4752
rect 5184 4712 5724 4740
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4672 1639 4675
rect 2869 4675 2927 4681
rect 2869 4672 2881 4675
rect 1627 4644 2881 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 2869 4641 2881 4644
rect 2915 4641 2927 4675
rect 3050 4672 3056 4684
rect 3011 4644 3056 4672
rect 2869 4635 2927 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 4706 4672 4712 4684
rect 4667 4644 4712 4672
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4856 4644 4905 4672
rect 4856 4632 4862 4644
rect 4893 4641 4905 4644
rect 4939 4672 4951 4675
rect 5184 4672 5212 4712
rect 5718 4700 5724 4712
rect 5776 4700 5782 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6273 4743 6331 4749
rect 6273 4740 6285 4743
rect 6052 4712 6285 4740
rect 6052 4700 6058 4712
rect 6273 4709 6285 4712
rect 6319 4709 6331 4743
rect 7300 4740 7328 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 8846 4740 8852 4752
rect 7300 4712 8852 4740
rect 6273 4703 6331 4709
rect 4939 4644 5212 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 5684 4644 5917 4672
rect 5684 4632 5690 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7852 4681 7880 4712
rect 8846 4700 8852 4712
rect 8904 4700 8910 4752
rect 10045 4743 10103 4749
rect 10045 4709 10057 4743
rect 10091 4740 10103 4743
rect 10318 4740 10324 4752
rect 10091 4712 10324 4740
rect 10091 4709 10103 4712
rect 10045 4703 10103 4709
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6880 4644 7389 4672
rect 6880 4632 6886 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4641 7895 4675
rect 9674 4672 9680 4684
rect 9635 4644 9680 4672
rect 7837 4635 7895 4641
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 5718 4604 5724 4616
rect 3191 4576 5724 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7668 4604 7696 4635
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4641 9919 4675
rect 9861 4635 9919 4641
rect 6972 4576 7696 4604
rect 6972 4564 6978 4576
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 9876 4604 9904 4635
rect 8352 4576 9904 4604
rect 8352 4564 8358 4576
rect 4893 4539 4951 4545
rect 4893 4505 4905 4539
rect 4939 4536 4951 4539
rect 7558 4536 7564 4548
rect 4939 4508 7564 4536
rect 4939 4505 4951 4508
rect 4893 4499 4951 4505
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 1104 4378 11592 4400
rect 1104 4326 2730 4378
rect 2782 4326 2794 4378
rect 2846 4326 2858 4378
rect 2910 4326 2922 4378
rect 2974 4326 6226 4378
rect 6278 4326 6290 4378
rect 6342 4326 6354 4378
rect 6406 4326 6418 4378
rect 6470 4326 9722 4378
rect 9774 4326 9786 4378
rect 9838 4326 9850 4378
rect 9902 4326 9914 4378
rect 9966 4326 11592 4378
rect 1104 4304 11592 4326
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5074 4264 5080 4276
rect 4764 4236 5080 4264
rect 4764 4224 4770 4236
rect 5074 4224 5080 4236
rect 5132 4264 5138 4276
rect 8570 4264 8576 4276
rect 5132 4236 8576 4264
rect 5132 4224 5138 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3694 4128 3700 4140
rect 3467 4100 3700 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 4798 4128 4804 4140
rect 4356 4100 4804 4128
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 2590 4060 2596 4072
rect 1443 4032 2596 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4029 3111 4063
rect 3234 4060 3240 4072
rect 3195 4032 3240 4060
rect 3053 4023 3111 4029
rect 3068 3992 3096 4023
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 4356 4069 4384 4100
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5408 4100 5457 4128
rect 5408 4088 5414 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 8202 4128 8208 4140
rect 6052 4100 8208 4128
rect 6052 4088 6058 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4128 8815 4131
rect 9582 4128 9588 4140
rect 8803 4100 9588 4128
rect 8803 4097 8815 4100
rect 8757 4091 8815 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10042 4128 10048 4140
rect 9784 4100 10048 4128
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4060 4583 4063
rect 5166 4060 5172 4072
rect 4571 4032 5172 4060
rect 4571 4029 4583 4032
rect 4525 4023 4583 4029
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6638 4060 6644 4072
rect 5675 4032 6644 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 6822 4060 6828 4072
rect 6783 4032 6828 4060
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7374 4060 7380 4072
rect 7335 4032 7380 4060
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 9122 4060 9128 4072
rect 7484 4032 9128 4060
rect 3602 3992 3608 4004
rect 3068 3964 3608 3992
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 4617 3995 4675 4001
rect 4617 3961 4629 3995
rect 4663 3992 4675 3995
rect 7484 3992 7512 4032
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9784 4069 9812 4100
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 4663 3964 7512 3992
rect 8389 3995 8447 4001
rect 4663 3961 4675 3964
rect 4617 3955 4675 3961
rect 8389 3961 8401 3995
rect 8435 3961 8447 3995
rect 8570 3992 8576 4004
rect 8531 3964 8576 3992
rect 8389 3955 8447 3961
rect 658 3884 664 3936
rect 716 3924 722 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 716 3896 1593 3924
rect 716 3884 722 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 4856 3896 5825 3924
rect 4856 3884 4862 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 7098 3924 7104 3936
rect 7059 3896 7104 3924
rect 5813 3887 5871 3893
rect 7098 3884 7104 3896
rect 7156 3924 7162 3936
rect 7558 3924 7564 3936
rect 7156 3896 7564 3924
rect 7156 3884 7162 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 8404 3924 8432 3955
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 9876 3992 9904 4023
rect 10042 3992 10048 4004
rect 9640 3964 9904 3992
rect 10003 3964 10048 3992
rect 9640 3952 9646 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10410 3924 10416 3936
rect 8404 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 1104 3834 11592 3856
rect 1104 3782 4478 3834
rect 4530 3782 4542 3834
rect 4594 3782 4606 3834
rect 4658 3782 4670 3834
rect 4722 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 11592 3834
rect 1104 3760 11592 3782
rect 5166 3720 5172 3732
rect 5127 3692 5172 3720
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 10042 3720 10048 3732
rect 7800 3692 10048 3720
rect 7800 3680 7806 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 5442 3652 5448 3664
rect 4396 3624 5448 3652
rect 4396 3612 4402 3624
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3584 2375 3587
rect 3970 3584 3976 3596
rect 2363 3556 3976 3584
rect 2363 3553 2375 3556
rect 2317 3547 2375 3553
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4798 3584 4804 3596
rect 4111 3556 4804 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5184 3593 5212 3624
rect 5442 3612 5448 3624
rect 5500 3652 5506 3664
rect 8570 3652 8576 3664
rect 5500 3624 8576 3652
rect 5500 3612 5506 3624
rect 8570 3612 8576 3624
rect 8628 3612 8634 3664
rect 10226 3652 10232 3664
rect 9784 3624 10232 3652
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3553 5227 3587
rect 5169 3547 5227 3553
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3584 5411 3587
rect 5994 3584 6000 3596
rect 5399 3556 6000 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 6144 3556 6285 3584
rect 6144 3544 6150 3556
rect 6273 3553 6285 3556
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 7190 3584 7196 3596
rect 6503 3556 7196 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 8662 3584 8668 3596
rect 8527 3556 8668 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 4430 3476 4436 3528
rect 4488 3516 4494 3528
rect 7742 3516 7748 3528
rect 4488 3488 7748 3516
rect 4488 3476 4494 3488
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 4249 3451 4307 3457
rect 4249 3417 4261 3451
rect 4295 3448 4307 3451
rect 6086 3448 6092 3460
rect 4295 3420 6092 3448
rect 4295 3417 4307 3420
rect 4249 3411 4307 3417
rect 6086 3408 6092 3420
rect 6144 3448 6150 3460
rect 8220 3448 8248 3547
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 9784 3593 9812 3624
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10502 3584 10508 3596
rect 10091 3556 10508 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 9876 3516 9904 3547
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 8619 3488 9904 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 6144 3420 8248 3448
rect 6144 3408 6150 3420
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2501 3383 2559 3389
rect 2501 3380 2513 3383
rect 2096 3352 2513 3380
rect 2096 3340 2102 3352
rect 2501 3349 2513 3352
rect 2547 3349 2559 3383
rect 2501 3343 2559 3349
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6273 3383 6331 3389
rect 6273 3380 6285 3383
rect 5868 3352 6285 3380
rect 5868 3340 5874 3352
rect 6273 3349 6285 3352
rect 6319 3349 6331 3383
rect 6273 3343 6331 3349
rect 1104 3290 11592 3312
rect 1104 3238 2730 3290
rect 2782 3238 2794 3290
rect 2846 3238 2858 3290
rect 2910 3238 2922 3290
rect 2974 3238 6226 3290
rect 6278 3238 6290 3290
rect 6342 3238 6354 3290
rect 6406 3238 6418 3290
rect 6470 3238 9722 3290
rect 9774 3238 9786 3290
rect 9838 3238 9850 3290
rect 9902 3238 9914 3290
rect 9966 3238 11592 3290
rect 1104 3216 11592 3238
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 3384 3148 4445 3176
rect 3384 3136 3390 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 6730 3176 6736 3188
rect 4433 3139 4491 3145
rect 4632 3148 6736 3176
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2941 3295 2975
rect 4430 2972 4436 2984
rect 4391 2944 4436 2972
rect 3237 2935 3295 2941
rect 3252 2904 3280 2935
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4632 2981 4660 3148
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 7834 3176 7840 3188
rect 6932 3148 7840 3176
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 6546 3108 6552 3120
rect 5859 3080 6552 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 6638 3068 6644 3120
rect 6696 3108 6702 3120
rect 6932 3108 6960 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8754 3176 8760 3188
rect 8435 3148 8760 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 10226 3176 10232 3188
rect 10187 3148 10232 3176
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 6696 3080 6960 3108
rect 7193 3111 7251 3117
rect 6696 3068 6702 3080
rect 7193 3077 7205 3111
rect 7239 3108 7251 3111
rect 8294 3108 8300 3120
rect 7239 3080 8300 3108
rect 7239 3077 7251 3080
rect 7193 3071 7251 3077
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 10134 3108 10140 3120
rect 8772 3080 10140 3108
rect 8772 3040 8800 3080
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 4816 3012 8800 3040
rect 8849 3043 8907 3049
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2941 4675 2975
rect 4617 2935 4675 2941
rect 4816 2904 4844 3012
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 10594 3040 10600 3052
rect 8895 3012 10600 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 5500 2944 5549 2972
rect 5500 2932 5506 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 5721 2975 5779 2981
rect 5721 2972 5733 2975
rect 5684 2944 5733 2972
rect 5684 2932 5690 2944
rect 5721 2941 5733 2944
rect 5767 2941 5779 2975
rect 5902 2972 5908 2984
rect 5815 2944 5908 2972
rect 5721 2935 5779 2941
rect 3252 2876 4844 2904
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 5828 2904 5856 2944
rect 5902 2932 5908 2944
rect 5960 2972 5966 2984
rect 8754 2972 8760 2984
rect 5960 2944 7236 2972
rect 8715 2944 8760 2972
rect 5960 2932 5966 2944
rect 4948 2876 5856 2904
rect 4948 2864 4954 2876
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 6825 2907 6883 2913
rect 6825 2904 6837 2907
rect 6696 2876 6837 2904
rect 6696 2864 6702 2876
rect 6825 2873 6837 2876
rect 6871 2873 6883 2907
rect 7006 2904 7012 2916
rect 6967 2876 7012 2904
rect 6825 2867 6883 2873
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7208 2904 7236 2944
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8864 2944 9137 2972
rect 8864 2904 8892 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 10137 2975 10195 2981
rect 10137 2972 10149 2975
rect 9355 2944 10149 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 10137 2941 10149 2944
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 11974 2972 11980 2984
rect 10459 2944 11980 2972
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 7208 2876 8892 2904
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9324 2904 9352 2935
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 9088 2876 9352 2904
rect 9088 2864 9094 2876
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 8754 2836 8760 2848
rect 3467 2808 8760 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 1104 2746 11592 2768
rect 1104 2694 4478 2746
rect 4530 2694 4542 2746
rect 4594 2694 4606 2746
rect 4658 2694 4670 2746
rect 4722 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 11592 2746
rect 1104 2672 11592 2694
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 6822 2632 6828 2644
rect 4755 2604 6828 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 6932 2604 7972 2632
rect 6932 2564 6960 2604
rect 7650 2564 7656 2576
rect 2884 2536 6960 2564
rect 7024 2536 7656 2564
rect 2884 2505 2912 2536
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 2869 2459 2927 2465
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 4724 2428 4752 2459
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 4856 2468 5641 2496
rect 4856 2456 4862 2468
rect 5629 2465 5641 2468
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 7024 2505 7052 2536
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 5776 2468 5825 2496
rect 5776 2456 5782 2468
rect 5813 2465 5825 2468
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7190 2496 7196 2508
rect 7151 2468 7196 2496
rect 7009 2459 7067 2465
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 7340 2468 7385 2496
rect 7340 2456 7346 2468
rect 7466 2428 7472 2440
rect 4724 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7944 2428 7972 2604
rect 8849 2567 8907 2573
rect 8849 2533 8861 2567
rect 8895 2564 8907 2567
rect 9030 2564 9036 2576
rect 8895 2536 9036 2564
rect 8895 2533 8907 2536
rect 8849 2527 8907 2533
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9180 2536 9965 2564
rect 9180 2524 9186 2536
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 10134 2564 10140 2576
rect 10095 2536 10140 2564
rect 9953 2527 10011 2533
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 8754 2496 8760 2508
rect 8715 2468 8760 2496
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10870 2496 10876 2508
rect 9815 2468 10876 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 9784 2428 9812 2459
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 7944 2400 9812 2428
rect 4982 2320 4988 2372
rect 5040 2360 5046 2372
rect 5905 2363 5963 2369
rect 5905 2360 5917 2363
rect 5040 2332 5917 2360
rect 5040 2320 5046 2332
rect 5905 2329 5917 2332
rect 5951 2329 5963 2363
rect 5905 2323 5963 2329
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 7742 2292 7748 2304
rect 3099 2264 7748 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 1104 2202 11592 2224
rect 1104 2150 2730 2202
rect 2782 2150 2794 2202
rect 2846 2150 2858 2202
rect 2910 2150 2922 2202
rect 2974 2150 6226 2202
rect 6278 2150 6290 2202
rect 6342 2150 6354 2202
rect 6406 2150 6418 2202
rect 6470 2150 9722 2202
rect 9774 2150 9786 2202
rect 9838 2150 9850 2202
rect 9902 2150 9914 2202
rect 9966 2150 11592 2202
rect 1104 2128 11592 2150
rect 4522 2048 4528 2100
rect 4580 2088 4586 2100
rect 7558 2088 7564 2100
rect 4580 2060 7564 2088
rect 4580 2048 4586 2060
rect 7558 2048 7564 2060
rect 7616 2048 7622 2100
<< via1 >>
rect 4478 12486 4530 12538
rect 4542 12486 4594 12538
rect 4606 12486 4658 12538
rect 4670 12486 4722 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 5632 12316 5684 12368
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 4252 12180 4304 12232
rect 4896 12248 4948 12300
rect 5908 12248 5960 12300
rect 7012 12180 7064 12232
rect 7748 12248 7800 12300
rect 10692 12248 10744 12300
rect 4160 12112 4212 12164
rect 7104 12044 7156 12096
rect 7564 12112 7616 12164
rect 7748 12044 7800 12096
rect 9588 12044 9640 12096
rect 2730 11942 2782 11994
rect 2794 11942 2846 11994
rect 2858 11942 2910 11994
rect 2922 11942 2974 11994
rect 6226 11942 6278 11994
rect 6290 11942 6342 11994
rect 6354 11942 6406 11994
rect 6418 11942 6470 11994
rect 9722 11942 9774 11994
rect 9786 11942 9838 11994
rect 9850 11942 9902 11994
rect 9914 11942 9966 11994
rect 2044 11704 2096 11756
rect 4068 11704 4120 11756
rect 3516 11636 3568 11688
rect 3884 11636 3936 11688
rect 4344 11679 4396 11688
rect 4344 11645 4353 11679
rect 4353 11645 4387 11679
rect 4387 11645 4396 11679
rect 4344 11636 4396 11645
rect 3700 11568 3752 11620
rect 5080 11636 5132 11688
rect 6920 11840 6972 11892
rect 7472 11772 7524 11824
rect 6552 11704 6604 11756
rect 9772 11704 9824 11756
rect 7104 11636 7156 11688
rect 7840 11568 7892 11620
rect 8484 11611 8536 11620
rect 8484 11577 8493 11611
rect 8493 11577 8527 11611
rect 8527 11577 8536 11611
rect 8484 11568 8536 11577
rect 3240 11543 3292 11552
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 4896 11500 4948 11552
rect 7012 11500 7064 11552
rect 7104 11500 7156 11552
rect 7748 11500 7800 11552
rect 8944 11568 8996 11620
rect 8668 11500 8720 11552
rect 4478 11398 4530 11450
rect 4542 11398 4594 11450
rect 4606 11398 4658 11450
rect 4670 11398 4722 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 4344 11296 4396 11348
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 5080 11228 5132 11280
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 3424 11160 3476 11212
rect 7012 11160 7064 11212
rect 3148 11092 3200 11144
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 6736 11092 6788 11144
rect 8392 11092 8444 11144
rect 3884 10956 3936 11008
rect 10048 11160 10100 11212
rect 8576 10956 8628 11008
rect 8760 10956 8812 11008
rect 10600 10956 10652 11008
rect 2730 10854 2782 10906
rect 2794 10854 2846 10906
rect 2858 10854 2910 10906
rect 2922 10854 2974 10906
rect 6226 10854 6278 10906
rect 6290 10854 6342 10906
rect 6354 10854 6406 10906
rect 6418 10854 6470 10906
rect 9722 10854 9774 10906
rect 9786 10854 9838 10906
rect 9850 10854 9902 10906
rect 9914 10854 9966 10906
rect 4160 10752 4212 10804
rect 7472 10752 7524 10804
rect 8576 10752 8628 10804
rect 9220 10752 9272 10804
rect 2780 10684 2832 10736
rect 3056 10616 3108 10668
rect 1860 10591 1912 10600
rect 1860 10557 1869 10591
rect 1869 10557 1903 10591
rect 1903 10557 1912 10591
rect 1860 10548 1912 10557
rect 2596 10548 2648 10600
rect 6920 10684 6972 10736
rect 7932 10616 7984 10668
rect 3608 10548 3660 10600
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 5632 10591 5684 10600
rect 4160 10480 4212 10532
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 7104 10548 7156 10600
rect 10324 10684 10376 10736
rect 8300 10616 8352 10668
rect 10048 10616 10100 10668
rect 8392 10548 8444 10600
rect 9220 10591 9272 10600
rect 4068 10412 4120 10464
rect 5908 10480 5960 10532
rect 6736 10480 6788 10532
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 8300 10480 8352 10532
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10508 10480 10560 10532
rect 11980 10480 12032 10532
rect 5080 10412 5132 10464
rect 6000 10412 6052 10464
rect 4478 10310 4530 10362
rect 4542 10310 4594 10362
rect 4606 10310 4658 10362
rect 4670 10310 4722 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 4252 10208 4304 10260
rect 5724 10208 5776 10260
rect 7472 10251 7524 10260
rect 7472 10217 7481 10251
rect 7481 10217 7515 10251
rect 7515 10217 7524 10251
rect 7472 10208 7524 10217
rect 9312 10208 9364 10260
rect 2964 10072 3016 10124
rect 4896 10140 4948 10192
rect 5632 10140 5684 10192
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5264 10072 5316 10124
rect 7472 10072 7524 10124
rect 7656 10072 7708 10124
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 9312 10072 9364 10124
rect 10140 10072 10192 10124
rect 2780 10004 2832 10056
rect 9404 10004 9456 10056
rect 10600 10004 10652 10056
rect 4252 9936 4304 9988
rect 3056 9868 3108 9920
rect 6000 9868 6052 9920
rect 6092 9868 6144 9920
rect 8392 9868 8444 9920
rect 9404 9868 9456 9920
rect 2730 9766 2782 9818
rect 2794 9766 2846 9818
rect 2858 9766 2910 9818
rect 2922 9766 2974 9818
rect 6226 9766 6278 9818
rect 6290 9766 6342 9818
rect 6354 9766 6406 9818
rect 6418 9766 6470 9818
rect 9722 9766 9774 9818
rect 9786 9766 9838 9818
rect 9850 9766 9902 9818
rect 9914 9766 9966 9818
rect 664 9664 716 9716
rect 2504 9664 2556 9716
rect 3608 9664 3660 9716
rect 8392 9664 8444 9716
rect 8576 9664 8628 9716
rect 9128 9664 9180 9716
rect 10048 9664 10100 9716
rect 3516 9528 3568 9580
rect 2596 9460 2648 9512
rect 5080 9596 5132 9648
rect 5632 9596 5684 9648
rect 7288 9639 7340 9648
rect 6644 9528 6696 9580
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 5540 9460 5592 9512
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 1952 9392 2004 9444
rect 10416 9460 10468 9512
rect 9404 9392 9456 9444
rect 10048 9435 10100 9444
rect 1584 9324 1636 9376
rect 3424 9324 3476 9376
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 7380 9324 7432 9376
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 10876 9392 10928 9444
rect 10232 9324 10284 9376
rect 4478 9222 4530 9274
rect 4542 9222 4594 9274
rect 4606 9222 4658 9274
rect 4670 9222 4722 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 1584 9095 1636 9104
rect 1584 9061 1593 9095
rect 1593 9061 1627 9095
rect 1627 9061 1636 9095
rect 1584 9052 1636 9061
rect 1952 9095 2004 9104
rect 1952 9061 1961 9095
rect 1961 9061 1995 9095
rect 1995 9061 2004 9095
rect 1952 9052 2004 9061
rect 4160 9052 4212 9104
rect 6552 9120 6604 9172
rect 8944 9120 8996 9172
rect 5080 9052 5132 9104
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 3700 8984 3752 9036
rect 4528 8984 4580 9036
rect 4620 9027 4672 9036
rect 4620 8993 4633 9027
rect 4633 8993 4667 9027
rect 4667 8993 4672 9027
rect 6552 9027 6604 9036
rect 4620 8984 4672 8993
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 6920 8984 6972 9036
rect 7748 8984 7800 9036
rect 4068 8916 4120 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 5632 8848 5684 8900
rect 6000 8916 6052 8968
rect 7196 8916 7248 8968
rect 7840 8916 7892 8968
rect 8024 8916 8076 8968
rect 10048 8848 10100 8900
rect 1676 8780 1728 8832
rect 4344 8780 4396 8832
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 2730 8678 2782 8730
rect 2794 8678 2846 8730
rect 2858 8678 2910 8730
rect 2922 8678 2974 8730
rect 6226 8678 6278 8730
rect 6290 8678 6342 8730
rect 6354 8678 6406 8730
rect 6418 8678 6470 8730
rect 9722 8678 9774 8730
rect 9786 8678 9838 8730
rect 9850 8678 9902 8730
rect 9914 8678 9966 8730
rect 2320 8576 2372 8628
rect 4804 8576 4856 8628
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 3608 8508 3660 8560
rect 3884 8508 3936 8560
rect 4068 8508 4120 8560
rect 4436 8508 4488 8560
rect 4988 8508 5040 8560
rect 7104 8508 7156 8560
rect 2504 8440 2556 8492
rect 6552 8440 6604 8492
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 4160 8372 4212 8424
rect 2596 8304 2648 8356
rect 4896 8304 4948 8356
rect 2780 8236 2832 8288
rect 4804 8236 4856 8288
rect 5080 8236 5132 8288
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 6460 8372 6512 8424
rect 7196 8440 7248 8492
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 7840 8508 7892 8560
rect 9312 8508 9364 8560
rect 9404 8508 9456 8560
rect 9680 8508 9732 8560
rect 7380 8440 7432 8492
rect 10232 8440 10284 8492
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 6092 8304 6144 8356
rect 7196 8304 7248 8356
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 7564 8236 7616 8288
rect 8024 8304 8076 8356
rect 8852 8304 8904 8356
rect 4478 8134 4530 8186
rect 4542 8134 4594 8186
rect 4606 8134 4658 8186
rect 4670 8134 4722 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 4068 8032 4120 8084
rect 4160 8032 4212 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 2872 7896 2924 7948
rect 4068 7896 4120 7948
rect 4252 7939 4304 7948
rect 4252 7905 4261 7939
rect 4261 7905 4295 7939
rect 4295 7905 4304 7939
rect 6184 8032 6236 8084
rect 6644 8032 6696 8084
rect 4252 7896 4304 7905
rect 4620 7896 4672 7948
rect 2780 7760 2832 7812
rect 3424 7828 3476 7880
rect 5632 7896 5684 7948
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 6552 7896 6604 7948
rect 7012 7964 7064 8016
rect 10692 7964 10744 8016
rect 7288 7939 7340 7948
rect 5908 7828 5960 7880
rect 6184 7828 6236 7880
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 8944 7896 8996 7948
rect 8484 7828 8536 7880
rect 4252 7760 4304 7812
rect 7472 7760 7524 7812
rect 9680 7828 9732 7880
rect 10416 7896 10468 7948
rect 7656 7692 7708 7744
rect 2730 7590 2782 7642
rect 2794 7590 2846 7642
rect 2858 7590 2910 7642
rect 2922 7590 2974 7642
rect 6226 7590 6278 7642
rect 6290 7590 6342 7642
rect 6354 7590 6406 7642
rect 6418 7590 6470 7642
rect 9722 7590 9774 7642
rect 9786 7590 9838 7642
rect 9850 7590 9902 7642
rect 9914 7590 9966 7642
rect 4344 7488 4396 7540
rect 5908 7488 5960 7540
rect 9496 7488 9548 7540
rect 7288 7420 7340 7472
rect 2412 7352 2464 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 7564 7420 7616 7472
rect 2688 7284 2740 7336
rect 3976 7284 4028 7336
rect 3332 7216 3384 7268
rect 3792 7216 3844 7268
rect 5632 7284 5684 7336
rect 6552 7284 6604 7336
rect 10600 7420 10652 7472
rect 7196 7216 7248 7268
rect 8668 7284 8720 7336
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 9128 7327 9180 7336
rect 8944 7284 8996 7293
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 7748 7148 7800 7200
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 4478 7046 4530 7098
rect 4542 7046 4594 7098
rect 4606 7046 4658 7098
rect 4670 7046 4722 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 5356 6944 5408 6996
rect 8668 6944 8720 6996
rect 4896 6876 4948 6928
rect 2504 6808 2556 6860
rect 3056 6808 3108 6860
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 4712 6808 4764 6860
rect 5080 6808 5132 6860
rect 5448 6808 5500 6860
rect 6000 6808 6052 6860
rect 6184 6808 6236 6860
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 7104 6808 7156 6860
rect 10232 6808 10284 6860
rect 7656 6740 7708 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 5908 6672 5960 6724
rect 6828 6672 6880 6724
rect 2320 6604 2372 6656
rect 10692 6672 10744 6724
rect 2730 6502 2782 6554
rect 2794 6502 2846 6554
rect 2858 6502 2910 6554
rect 2922 6502 2974 6554
rect 6226 6502 6278 6554
rect 6290 6502 6342 6554
rect 6354 6502 6406 6554
rect 6418 6502 6470 6554
rect 9722 6502 9774 6554
rect 9786 6502 9838 6554
rect 9850 6502 9902 6554
rect 9914 6502 9966 6554
rect 8944 6400 8996 6452
rect 3792 6332 3844 6384
rect 2412 6196 2464 6248
rect 5356 6264 5408 6316
rect 5540 6264 5592 6316
rect 6828 6264 6880 6316
rect 4160 6196 4212 6248
rect 6276 6196 6328 6248
rect 9220 6239 9272 6248
rect 4712 6128 4764 6180
rect 6092 6128 6144 6180
rect 4804 6060 4856 6112
rect 5540 6060 5592 6112
rect 6736 6060 6788 6112
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 9864 6264 9916 6316
rect 10140 6264 10192 6316
rect 9496 6196 9548 6248
rect 10048 6196 10100 6248
rect 7472 6128 7524 6180
rect 4478 5958 4530 6010
rect 4542 5958 4594 6010
rect 4606 5958 4658 6010
rect 4670 5958 4722 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 2504 5856 2556 5908
rect 1768 5788 1820 5840
rect 7840 5856 7892 5908
rect 3056 5788 3108 5840
rect 6000 5720 6052 5772
rect 6644 5720 6696 5772
rect 7012 5763 7064 5772
rect 7012 5729 7021 5763
rect 7021 5729 7055 5763
rect 7055 5729 7064 5763
rect 7012 5720 7064 5729
rect 7840 5720 7892 5772
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 8760 5763 8812 5772
rect 8760 5729 8769 5763
rect 8769 5729 8803 5763
rect 8803 5729 8812 5763
rect 8760 5720 8812 5729
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 3056 5652 3108 5704
rect 3976 5652 4028 5704
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 6736 5584 6788 5636
rect 7196 5584 7248 5636
rect 5356 5516 5408 5568
rect 5448 5516 5500 5568
rect 5724 5516 5776 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 10048 5516 10100 5568
rect 2730 5414 2782 5466
rect 2794 5414 2846 5466
rect 2858 5414 2910 5466
rect 2922 5414 2974 5466
rect 6226 5414 6278 5466
rect 6290 5414 6342 5466
rect 6354 5414 6406 5466
rect 6418 5414 6470 5466
rect 9722 5414 9774 5466
rect 9786 5414 9838 5466
rect 9850 5414 9902 5466
rect 9914 5414 9966 5466
rect 6920 5312 6972 5364
rect 7196 5312 7248 5364
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 7656 5244 7708 5296
rect 3056 5176 3108 5228
rect 9312 5176 9364 5228
rect 3424 5108 3476 5160
rect 5448 5108 5500 5160
rect 6000 5108 6052 5160
rect 8576 5151 8628 5160
rect 8576 5117 8585 5151
rect 8585 5117 8619 5151
rect 8619 5117 8628 5151
rect 8576 5108 8628 5117
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 5632 5040 5684 5092
rect 5724 5083 5776 5092
rect 5724 5049 5733 5083
rect 5733 5049 5767 5083
rect 5767 5049 5776 5083
rect 5724 5040 5776 5049
rect 6644 5040 6696 5092
rect 7472 5040 7524 5092
rect 8300 5040 8352 5092
rect 10692 5040 10744 5092
rect 7840 4972 7892 5024
rect 4478 4870 4530 4922
rect 4542 4870 4594 4922
rect 4606 4870 4658 4922
rect 4670 4870 4722 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 7472 4811 7524 4820
rect 1768 4743 1820 4752
rect 1768 4709 1777 4743
rect 1777 4709 1811 4743
rect 1811 4709 1820 4743
rect 1768 4700 1820 4709
rect 4160 4700 4212 4752
rect 4988 4700 5040 4752
rect 3056 4675 3108 4684
rect 3056 4641 3065 4675
rect 3065 4641 3099 4675
rect 3099 4641 3108 4675
rect 3056 4632 3108 4641
rect 4712 4675 4764 4684
rect 4712 4641 4721 4675
rect 4721 4641 4755 4675
rect 4755 4641 4764 4675
rect 4712 4632 4764 4641
rect 4804 4632 4856 4684
rect 5724 4700 5776 4752
rect 6000 4700 6052 4752
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 5632 4632 5684 4684
rect 6828 4632 6880 4684
rect 8852 4700 8904 4752
rect 10324 4700 10376 4752
rect 9680 4675 9732 4684
rect 5724 4564 5776 4616
rect 6920 4564 6972 4616
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 8300 4564 8352 4616
rect 7564 4496 7616 4548
rect 2730 4326 2782 4378
rect 2794 4326 2846 4378
rect 2858 4326 2910 4378
rect 2922 4326 2974 4378
rect 6226 4326 6278 4378
rect 6290 4326 6342 4378
rect 6354 4326 6406 4378
rect 6418 4326 6470 4378
rect 9722 4326 9774 4378
rect 9786 4326 9838 4378
rect 9850 4326 9902 4378
rect 9914 4326 9966 4378
rect 4712 4224 4764 4276
rect 5080 4224 5132 4276
rect 8576 4224 8628 4276
rect 3700 4088 3752 4140
rect 2596 4020 2648 4072
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 4804 4088 4856 4140
rect 5356 4088 5408 4140
rect 6000 4088 6052 4140
rect 8208 4088 8260 4140
rect 9588 4088 9640 4140
rect 5172 4020 5224 4072
rect 6644 4020 6696 4072
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 7380 4063 7432 4072
rect 7380 4029 7389 4063
rect 7389 4029 7423 4063
rect 7423 4029 7432 4063
rect 7380 4020 7432 4029
rect 3608 3952 3660 4004
rect 9128 4020 9180 4072
rect 10048 4088 10100 4140
rect 8576 3995 8628 4004
rect 664 3884 716 3936
rect 4804 3884 4856 3936
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 7564 3884 7616 3936
rect 8576 3961 8585 3995
rect 8585 3961 8619 3995
rect 8619 3961 8628 3995
rect 8576 3952 8628 3961
rect 9588 3952 9640 4004
rect 10048 3995 10100 4004
rect 10048 3961 10057 3995
rect 10057 3961 10091 3995
rect 10091 3961 10100 3995
rect 10048 3952 10100 3961
rect 10416 3884 10468 3936
rect 4478 3782 4530 3834
rect 4542 3782 4594 3834
rect 4606 3782 4658 3834
rect 4670 3782 4722 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 7748 3680 7800 3732
rect 10048 3680 10100 3732
rect 4344 3612 4396 3664
rect 3976 3544 4028 3596
rect 4804 3544 4856 3596
rect 5448 3612 5500 3664
rect 8576 3612 8628 3664
rect 6000 3544 6052 3596
rect 6092 3544 6144 3596
rect 7196 3544 7248 3596
rect 4436 3476 4488 3528
rect 7748 3476 7800 3528
rect 6092 3408 6144 3460
rect 8668 3544 8720 3596
rect 10232 3612 10284 3664
rect 10508 3544 10560 3596
rect 2044 3340 2096 3392
rect 5816 3340 5868 3392
rect 2730 3238 2782 3290
rect 2794 3238 2846 3290
rect 2858 3238 2910 3290
rect 2922 3238 2974 3290
rect 6226 3238 6278 3290
rect 6290 3238 6342 3290
rect 6354 3238 6406 3290
rect 6418 3238 6470 3290
rect 9722 3238 9774 3290
rect 9786 3238 9838 3290
rect 9850 3238 9902 3290
rect 9914 3238 9966 3290
rect 3332 3136 3384 3188
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 6736 3136 6788 3188
rect 6552 3068 6604 3120
rect 6644 3068 6696 3120
rect 7840 3136 7892 3188
rect 8760 3136 8812 3188
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 8300 3068 8352 3120
rect 10140 3068 10192 3120
rect 10600 3000 10652 3052
rect 5448 2932 5500 2984
rect 5632 2932 5684 2984
rect 4896 2864 4948 2916
rect 5908 2932 5960 2984
rect 8760 2975 8812 2984
rect 6644 2864 6696 2916
rect 7012 2907 7064 2916
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7012 2864 7064 2873
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 9036 2864 9088 2916
rect 11980 2932 12032 2984
rect 8760 2796 8812 2848
rect 4478 2694 4530 2746
rect 4542 2694 4594 2746
rect 4606 2694 4658 2746
rect 4670 2694 4722 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 6828 2592 6880 2644
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 4804 2456 4856 2508
rect 5724 2456 5776 2508
rect 7656 2524 7708 2576
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 7472 2388 7524 2440
rect 9036 2524 9088 2576
rect 9128 2524 9180 2576
rect 10140 2567 10192 2576
rect 10140 2533 10149 2567
rect 10149 2533 10183 2567
rect 10183 2533 10192 2567
rect 10140 2524 10192 2533
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 10876 2456 10928 2508
rect 4988 2320 5040 2372
rect 7748 2252 7800 2304
rect 2730 2150 2782 2202
rect 2794 2150 2846 2202
rect 2858 2150 2910 2202
rect 2922 2150 2974 2202
rect 6226 2150 6278 2202
rect 6290 2150 6342 2202
rect 6354 2150 6406 2202
rect 6418 2150 6470 2202
rect 9722 2150 9774 2202
rect 9786 2150 9838 2202
rect 9850 2150 9902 2202
rect 9914 2150 9966 2202
rect 4528 2048 4580 2100
rect 7564 2048 7616 2100
<< metal2 >>
rect 662 14113 718 14913
rect 2042 14113 2098 14913
rect 3422 14113 3478 14913
rect 4894 14113 4950 14913
rect 6274 14113 6330 14913
rect 7746 14113 7802 14913
rect 9126 14113 9182 14913
rect 10598 14113 10654 14913
rect 11978 14113 12034 14913
rect 676 9722 704 14113
rect 2056 11762 2084 14113
rect 2704 11996 3000 12016
rect 2760 11994 2784 11996
rect 2840 11994 2864 11996
rect 2920 11994 2944 11996
rect 2782 11942 2784 11994
rect 2846 11942 2858 11994
rect 2920 11942 2922 11994
rect 2760 11940 2784 11942
rect 2840 11940 2864 11942
rect 2920 11940 2944 11942
rect 2704 11920 3000 11940
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 1858 11248 1914 11257
rect 1858 11183 1914 11192
rect 3056 11212 3108 11218
rect 1872 10606 1900 11183
rect 3056 11154 3108 11160
rect 2704 10908 3000 10928
rect 2760 10906 2784 10908
rect 2840 10906 2864 10908
rect 2920 10906 2944 10908
rect 2782 10854 2784 10906
rect 2846 10854 2858 10906
rect 2920 10854 2922 10906
rect 2760 10852 2784 10854
rect 2840 10852 2864 10854
rect 2920 10852 2944 10854
rect 2704 10832 3000 10852
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 664 9716 716 9722
rect 664 9658 716 9664
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9110 1624 9318
rect 1964 9110 1992 9386
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1676 8832 1728 8838
rect 1490 8800 1546 8809
rect 1676 8774 1728 8780
rect 1490 8735 1546 8744
rect 1504 8430 1532 8735
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1688 7954 1716 8774
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 2332 6662 2360 8570
rect 2516 8498 2544 9658
rect 2608 9518 2636 10542
rect 2792 10062 2820 10678
rect 3068 10674 3096 11154
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2976 10010 3004 10066
rect 2976 9982 3096 10010
rect 3068 9926 3096 9982
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2704 9820 3000 9840
rect 2760 9818 2784 9820
rect 2840 9818 2864 9820
rect 2920 9818 2944 9820
rect 2782 9766 2784 9818
rect 2846 9766 2858 9818
rect 2920 9766 2922 9818
rect 2760 9764 2784 9766
rect 2840 9764 2864 9766
rect 2920 9764 2944 9766
rect 2704 9744 3000 9764
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6225 2360 6598
rect 2424 6254 2452 7346
rect 2516 7290 2544 8434
rect 2608 8362 2636 9454
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2884 8945 2912 8978
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 2704 8732 3000 8752
rect 2760 8730 2784 8732
rect 2840 8730 2864 8732
rect 2920 8730 2944 8732
rect 2782 8678 2784 8730
rect 2846 8678 2858 8730
rect 2920 8678 2922 8730
rect 2760 8676 2784 8678
rect 2840 8676 2864 8678
rect 2920 8676 2944 8678
rect 2704 8656 3000 8676
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2608 7460 2636 8298
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7818 2820 8230
rect 3068 8106 3096 9862
rect 2884 8078 3096 8106
rect 2884 7954 2912 8078
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2704 7644 3000 7664
rect 2760 7642 2784 7644
rect 2840 7642 2864 7644
rect 2920 7642 2944 7644
rect 2782 7590 2784 7642
rect 2846 7590 2858 7642
rect 2920 7590 2922 7642
rect 2760 7588 2784 7590
rect 2840 7588 2864 7590
rect 2920 7588 2944 7590
rect 2704 7568 3000 7588
rect 2608 7432 2728 7460
rect 2700 7342 2728 7432
rect 3160 7410 3188 11086
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2688 7336 2740 7342
rect 2516 7262 2636 7290
rect 2688 7278 2740 7284
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2412 6248 2464 6254
rect 2318 6216 2374 6225
rect 2412 6190 2464 6196
rect 2318 6151 2374 6160
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1780 4758 1808 5782
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 664 3936 716 3942
rect 664 3878 716 3884
rect 676 800 704 3878
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 800 2084 3334
rect 2424 1329 2452 6190
rect 2516 5914 2544 6802
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2608 4078 2636 7262
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2704 6556 3000 6576
rect 2760 6554 2784 6556
rect 2840 6554 2864 6556
rect 2920 6554 2944 6556
rect 2782 6502 2784 6554
rect 2846 6502 2858 6554
rect 2920 6502 2922 6554
rect 2760 6500 2784 6502
rect 2840 6500 2864 6502
rect 2920 6500 2944 6502
rect 2704 6480 3000 6500
rect 3068 5846 3096 6802
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2704 5468 3000 5488
rect 2760 5466 2784 5468
rect 2840 5466 2864 5468
rect 2920 5466 2944 5468
rect 2782 5414 2784 5466
rect 2846 5414 2858 5466
rect 2920 5414 2922 5466
rect 2760 5412 2784 5414
rect 2840 5412 2864 5414
rect 2920 5412 2944 5414
rect 2704 5392 3000 5412
rect 3068 5234 3096 5646
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2704 4380 3000 4400
rect 2760 4378 2784 4380
rect 2840 4378 2864 4380
rect 2920 4378 2944 4380
rect 2782 4326 2784 4378
rect 2846 4326 2858 4378
rect 2920 4326 2922 4378
rect 2760 4324 2784 4326
rect 2840 4324 2864 4326
rect 2920 4324 2944 4326
rect 2704 4304 3000 4324
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2704 3292 3000 3312
rect 2760 3290 2784 3292
rect 2840 3290 2864 3292
rect 2920 3290 2944 3292
rect 2782 3238 2784 3290
rect 2846 3238 2858 3290
rect 2920 3238 2922 3290
rect 2760 3236 2784 3238
rect 2840 3236 2864 3238
rect 2920 3236 2944 3238
rect 2704 3216 3000 3236
rect 3068 2553 3096 4626
rect 3252 4078 3280 11494
rect 3436 11218 3464 14113
rect 3606 13696 3662 13705
rect 3606 13631 3662 13640
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3528 11064 3556 11630
rect 3436 11036 3556 11064
rect 3436 9382 3464 11036
rect 3620 10996 3648 13631
rect 4452 12540 4748 12560
rect 4508 12538 4532 12540
rect 4588 12538 4612 12540
rect 4668 12538 4692 12540
rect 4530 12486 4532 12538
rect 4594 12486 4606 12538
rect 4668 12486 4670 12538
rect 4508 12484 4532 12486
rect 4588 12484 4612 12486
rect 4668 12484 4692 12486
rect 4452 12464 4748 12484
rect 4908 12306 4936 14113
rect 6288 12594 6316 14113
rect 6288 12566 6500 12594
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3528 10968 3648 10996
rect 3528 9586 3556 10968
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 9722 3648 10542
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 7886 3464 9318
rect 3712 9042 3740 11562
rect 3896 11014 3924 11630
rect 4080 11150 4108 11698
rect 4068 11144 4120 11150
rect 3988 11104 4068 11132
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3344 3777 3372 7210
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3330 3768 3386 3777
rect 3330 3703 3386 3712
rect 3344 3194 3372 3703
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3054 2544 3110 2553
rect 3054 2479 3110 2488
rect 2704 2204 3000 2224
rect 2760 2202 2784 2204
rect 2840 2202 2864 2204
rect 2920 2202 2944 2204
rect 2782 2150 2784 2202
rect 2846 2150 2858 2202
rect 2920 2150 2922 2202
rect 2760 2148 2784 2150
rect 2840 2148 2864 2150
rect 2920 2148 2944 2150
rect 2704 2128 3000 2148
rect 2410 1320 2466 1329
rect 2410 1255 2466 1264
rect 3436 800 3464 5102
rect 3620 4010 3648 8502
rect 3712 4146 3740 8978
rect 3896 8566 3924 10950
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3988 7342 4016 11104
rect 4068 11086 4120 11092
rect 4172 10810 4200 12106
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 8974 4108 10406
rect 4172 9110 4200 10474
rect 4264 10266 4292 12174
rect 4356 11694 4384 12242
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4452 11452 4748 11472
rect 4508 11450 4532 11452
rect 4588 11450 4612 11452
rect 4668 11450 4692 11452
rect 4530 11398 4532 11450
rect 4594 11398 4606 11450
rect 4668 11398 4670 11450
rect 4508 11396 4532 11398
rect 4588 11396 4612 11398
rect 4668 11396 4692 11398
rect 4452 11376 4748 11396
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4356 10146 4384 11290
rect 4436 10600 4488 10606
rect 4488 10560 4844 10588
rect 4436 10542 4488 10548
rect 4452 10364 4748 10384
rect 4508 10362 4532 10364
rect 4588 10362 4612 10364
rect 4668 10362 4692 10364
rect 4530 10310 4532 10362
rect 4594 10310 4606 10362
rect 4668 10310 4670 10362
rect 4508 10308 4532 10310
rect 4588 10308 4612 10310
rect 4668 10308 4692 10310
rect 4452 10288 4748 10308
rect 4264 10118 4384 10146
rect 4816 10130 4844 10560
rect 4908 10198 4936 11494
rect 5092 11286 5120 11630
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5092 10554 5120 11222
rect 5644 10606 5672 12310
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5000 10526 5120 10554
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4804 10124 4856 10130
rect 4264 9994 4292 10118
rect 4804 10066 4856 10072
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4080 8090 4108 8502
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4172 8090 4200 8366
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4264 7954 4292 9930
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 8838 4384 9318
rect 4452 9276 4748 9296
rect 4508 9274 4532 9276
rect 4588 9274 4612 9276
rect 4668 9274 4692 9276
rect 4530 9222 4532 9274
rect 4594 9222 4606 9274
rect 4668 9222 4670 9274
rect 4508 9220 4532 9222
rect 4588 9220 4612 9222
rect 4668 9220 4692 9222
rect 4452 9200 4748 9220
rect 4528 9036 4580 9042
rect 4620 9036 4672 9042
rect 4580 8996 4620 9024
rect 4528 8978 4580 8984
rect 4620 8978 4672 8984
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4816 8922 4844 10066
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4448 8566 4476 8910
rect 4816 8894 4936 8922
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8634 4844 8774
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4908 8362 4936 8894
rect 5000 8566 5028 10526
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 10130 5120 10406
rect 5644 10198 5672 10542
rect 5920 10538 5948 12242
rect 6472 12084 6500 12566
rect 7760 12306 7788 14113
rect 7948 12540 8244 12560
rect 8004 12538 8028 12540
rect 8084 12538 8108 12540
rect 8164 12538 8188 12540
rect 8026 12486 8028 12538
rect 8090 12486 8102 12538
rect 8164 12486 8166 12538
rect 8004 12484 8028 12486
rect 8084 12484 8108 12486
rect 8164 12484 8188 12486
rect 7948 12464 8244 12484
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6472 12056 6592 12084
rect 6200 11996 6496 12016
rect 6256 11994 6280 11996
rect 6336 11994 6360 11996
rect 6416 11994 6440 11996
rect 6278 11942 6280 11994
rect 6342 11942 6354 11994
rect 6416 11942 6418 11994
rect 6256 11940 6280 11942
rect 6336 11940 6360 11942
rect 6416 11940 6440 11942
rect 6200 11920 6496 11940
rect 6564 11762 6592 12056
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6200 10908 6496 10928
rect 6256 10906 6280 10908
rect 6336 10906 6360 10908
rect 6416 10906 6440 10908
rect 6278 10854 6280 10906
rect 6342 10854 6354 10906
rect 6416 10854 6418 10906
rect 6256 10852 6280 10854
rect 6336 10852 6360 10854
rect 6416 10852 6440 10854
rect 6200 10832 6496 10852
rect 6748 10538 6776 11086
rect 6932 10742 6960 11834
rect 7024 11558 7052 12174
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11694 7144 12038
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7024 11218 7052 11494
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5092 9110 5120 9590
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4452 8188 4748 8208
rect 4508 8186 4532 8188
rect 4588 8186 4612 8188
rect 4668 8186 4692 8188
rect 4530 8134 4532 8186
rect 4594 8134 4606 8186
rect 4668 8134 4670 8186
rect 4508 8132 4532 8134
rect 4588 8132 4612 8134
rect 4668 8132 4692 8134
rect 4452 8112 4748 8132
rect 4816 7970 4844 8230
rect 4632 7954 4844 7970
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4620 7948 4844 7954
rect 4672 7942 4844 7948
rect 4620 7890 4672 7896
rect 4080 7698 4108 7890
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4264 7698 4292 7754
rect 4080 7670 4292 7698
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 6390 3832 7210
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3988 5710 4016 7278
rect 4356 6866 4384 7482
rect 4452 7100 4748 7120
rect 4508 7098 4532 7100
rect 4588 7098 4612 7100
rect 4668 7098 4692 7100
rect 4530 7046 4532 7098
rect 4594 7046 4606 7098
rect 4668 7046 4670 7098
rect 4508 7044 4532 7046
rect 4588 7044 4612 7046
rect 4668 7044 4692 7046
rect 4452 7024 4748 7044
rect 4908 6934 4936 8298
rect 5092 8294 5120 9046
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3988 3602 4016 5646
rect 4172 4758 4200 6190
rect 4356 5710 4384 6802
rect 4724 6186 4752 6802
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4452 6012 4748 6032
rect 4508 6010 4532 6012
rect 4588 6010 4612 6012
rect 4668 6010 4692 6012
rect 4530 5958 4532 6010
rect 4594 5958 4606 6010
rect 4668 5958 4670 6010
rect 4508 5956 4532 5958
rect 4588 5956 4612 5958
rect 4668 5956 4692 5958
rect 4452 5936 4748 5956
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4356 3670 4384 5646
rect 4452 4924 4748 4944
rect 4508 4922 4532 4924
rect 4588 4922 4612 4924
rect 4668 4922 4692 4924
rect 4530 4870 4532 4922
rect 4594 4870 4606 4922
rect 4668 4870 4670 4922
rect 4508 4868 4532 4870
rect 4588 4868 4612 4870
rect 4668 4868 4692 4870
rect 4452 4848 4748 4868
rect 4816 4690 4844 6054
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4724 4282 4752 4626
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4816 4146 4844 4626
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4452 3836 4748 3856
rect 4508 3834 4532 3836
rect 4588 3834 4612 3836
rect 4668 3834 4692 3836
rect 4530 3782 4532 3834
rect 4594 3782 4606 3834
rect 4668 3782 4670 3834
rect 4508 3780 4532 3782
rect 4588 3780 4612 3782
rect 4668 3780 4692 3782
rect 4452 3760 4748 3780
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4816 3602 4844 3878
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4436 3528 4488 3534
rect 4908 3482 4936 6870
rect 5080 6860 5132 6866
rect 5276 6848 5304 10066
rect 5644 9738 5672 10134
rect 5552 9710 5672 9738
rect 5552 9518 5580 9710
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5132 6820 5304 6848
rect 5080 6802 5132 6808
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4436 3470 4488 3476
rect 4448 2990 4476 3470
rect 4816 3454 4936 3482
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4452 2748 4748 2768
rect 4508 2746 4532 2748
rect 4588 2746 4612 2748
rect 4668 2746 4692 2748
rect 4530 2694 4532 2746
rect 4594 2694 4606 2746
rect 4668 2694 4670 2746
rect 4508 2692 4532 2694
rect 4588 2692 4612 2694
rect 4668 2692 4692 2694
rect 4452 2672 4748 2692
rect 4816 2514 4844 3454
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4540 2106 4568 2450
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 4908 800 4936 2858
rect 5000 2378 5028 4694
rect 5092 4282 5120 6802
rect 5368 6322 5396 6938
rect 5460 6866 5488 9454
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5552 6322 5580 9454
rect 5644 8906 5672 9590
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 7954 5672 8842
rect 5736 8430 5764 10202
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5644 6202 5672 7278
rect 5552 6174 5672 6202
rect 5552 6118 5580 6174
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5368 4146 5396 5510
rect 5460 5166 5488 5510
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5552 4570 5580 6054
rect 5736 5574 5764 8366
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5644 4690 5672 5034
rect 5736 4758 5764 5034
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5724 4616 5776 4622
rect 5552 4542 5672 4570
rect 5724 4558 5776 4564
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5184 3738 5212 4014
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5460 2990 5488 3606
rect 5644 2990 5672 4542
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5736 2514 5764 4558
rect 5828 3398 5856 9318
rect 5920 7970 5948 10474
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 9926 6040 10406
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6012 8974 6040 9862
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6104 8362 6132 9862
rect 6200 9820 6496 9840
rect 6256 9818 6280 9820
rect 6336 9818 6360 9820
rect 6416 9818 6440 9820
rect 6278 9766 6280 9818
rect 6342 9766 6354 9818
rect 6416 9766 6418 9818
rect 6256 9764 6280 9766
rect 6336 9764 6360 9766
rect 6416 9764 6440 9766
rect 6200 9744 6496 9764
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6564 9042 6592 9114
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6200 8732 6496 8752
rect 6256 8730 6280 8732
rect 6336 8730 6360 8732
rect 6416 8730 6440 8732
rect 6278 8678 6280 8730
rect 6342 8678 6354 8730
rect 6416 8678 6418 8730
rect 6256 8676 6280 8678
rect 6336 8676 6360 8678
rect 6416 8676 6440 8678
rect 6200 8656 6496 8676
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5920 7942 6132 7970
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7546 5948 7822
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6104 6848 6132 7942
rect 6196 7886 6224 8026
rect 6472 7993 6500 8366
rect 6458 7984 6514 7993
rect 6564 7954 6592 8434
rect 6656 8090 6684 9522
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6458 7919 6460 7928
rect 6512 7919 6514 7928
rect 6552 7948 6604 7954
rect 6460 7890 6512 7896
rect 6552 7890 6604 7896
rect 6184 7880 6236 7886
rect 6472 7859 6500 7890
rect 6184 7822 6236 7828
rect 6200 7644 6496 7664
rect 6256 7642 6280 7644
rect 6336 7642 6360 7644
rect 6416 7642 6440 7644
rect 6278 7590 6280 7642
rect 6342 7590 6354 7642
rect 6416 7590 6418 7642
rect 6256 7588 6280 7590
rect 6336 7588 6360 7590
rect 6416 7588 6440 7590
rect 6200 7568 6496 7588
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6184 6860 6236 6866
rect 6104 6820 6184 6848
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5920 2990 5948 6666
rect 6012 5778 6040 6802
rect 6104 6338 6132 6820
rect 6184 6802 6236 6808
rect 6200 6556 6496 6576
rect 6256 6554 6280 6556
rect 6336 6554 6360 6556
rect 6416 6554 6440 6556
rect 6278 6502 6280 6554
rect 6342 6502 6354 6554
rect 6416 6502 6418 6554
rect 6256 6500 6280 6502
rect 6336 6500 6360 6502
rect 6416 6500 6440 6502
rect 6200 6480 6496 6500
rect 6104 6310 6316 6338
rect 6288 6254 6316 6310
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6012 5166 6040 5714
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6012 4758 6040 5102
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6012 3602 6040 4082
rect 6104 3602 6132 6122
rect 6288 5681 6316 6190
rect 6274 5672 6330 5681
rect 6274 5607 6330 5616
rect 6200 5468 6496 5488
rect 6256 5466 6280 5468
rect 6336 5466 6360 5468
rect 6416 5466 6440 5468
rect 6278 5414 6280 5466
rect 6342 5414 6354 5466
rect 6416 5414 6418 5466
rect 6256 5412 6280 5414
rect 6336 5412 6360 5414
rect 6416 5412 6440 5414
rect 6200 5392 6496 5412
rect 6200 4380 6496 4400
rect 6256 4378 6280 4380
rect 6336 4378 6360 4380
rect 6416 4378 6440 4380
rect 6278 4326 6280 4378
rect 6342 4326 6354 4378
rect 6416 4326 6418 4378
rect 6256 4324 6280 4326
rect 6336 4324 6360 4326
rect 6416 4324 6440 4326
rect 6200 4304 6496 4324
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 6104 1986 6132 3402
rect 6200 3292 6496 3312
rect 6256 3290 6280 3292
rect 6336 3290 6360 3292
rect 6416 3290 6440 3292
rect 6278 3238 6280 3290
rect 6342 3238 6354 3290
rect 6416 3238 6418 3290
rect 6256 3236 6280 3238
rect 6336 3236 6360 3238
rect 6416 3236 6440 3238
rect 6200 3216 6496 3236
rect 6564 3126 6592 7278
rect 6748 6118 6776 10474
rect 6932 9042 6960 10678
rect 7116 10606 7144 11494
rect 7484 10810 7512 11766
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6826 8936 6882 8945
rect 6826 8871 6882 8880
rect 6840 8430 6868 8871
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 6866 6868 8366
rect 7024 8106 7052 10474
rect 7116 8566 7144 10542
rect 7484 10266 7512 10746
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 9330 7328 9590
rect 7380 9376 7432 9382
rect 7300 9324 7380 9330
rect 7300 9318 7432 9324
rect 7300 9302 7420 9318
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7208 8498 7236 8910
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6932 8078 7052 8106
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6932 6746 6960 8078
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7024 6866 7052 7958
rect 7116 6866 7144 8366
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7208 7460 7236 8298
rect 7300 7954 7328 9302
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7288 7472 7340 7478
rect 7208 7432 7288 7460
rect 7288 7414 7340 7420
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 6828 6724 6880 6730
rect 6932 6718 7052 6746
rect 6828 6666 6880 6672
rect 6840 6440 6868 6666
rect 6840 6412 6960 6440
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6656 5098 6684 5714
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6656 3738 6684 4014
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3194 6776 5578
rect 6840 4690 6868 6258
rect 6932 5370 6960 6412
rect 7024 5778 7052 6718
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6932 4622 6960 5199
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6656 2922 6684 3062
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6840 2650 6868 4014
rect 7024 2922 7052 5510
rect 7116 3942 7144 6802
rect 7208 5642 7236 7210
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7208 3602 7236 5306
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7300 3482 7328 7414
rect 7392 4078 7420 8434
rect 7484 7818 7512 10066
rect 7576 8430 7604 12106
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11558 7788 12038
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7576 7698 7604 8230
rect 7668 7750 7696 10066
rect 7760 9160 7788 11494
rect 7852 11354 7880 11562
rect 7948 11452 8244 11472
rect 8004 11450 8028 11452
rect 8084 11450 8108 11452
rect 8164 11450 8188 11452
rect 8026 11398 8028 11450
rect 8090 11398 8102 11450
rect 8164 11398 8166 11450
rect 8004 11396 8028 11398
rect 8084 11396 8108 11398
rect 8164 11396 8188 11398
rect 7948 11376 8244 11396
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 7932 10668 7984 10674
rect 8300 10668 8352 10674
rect 7984 10628 8300 10656
rect 7932 10610 7984 10616
rect 8300 10610 8352 10616
rect 8404 10606 8432 11086
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 7948 10364 8244 10384
rect 8004 10362 8028 10364
rect 8084 10362 8108 10364
rect 8164 10362 8188 10364
rect 8026 10310 8028 10362
rect 8090 10310 8102 10362
rect 8164 10310 8166 10362
rect 8004 10308 8028 10310
rect 8084 10308 8108 10310
rect 8164 10308 8188 10310
rect 7948 10288 8244 10308
rect 7948 9276 8244 9296
rect 8004 9274 8028 9276
rect 8084 9274 8108 9276
rect 8164 9274 8188 9276
rect 8026 9222 8028 9274
rect 8090 9222 8102 9274
rect 8164 9222 8166 9274
rect 8004 9220 8028 9222
rect 8084 9220 8108 9222
rect 8164 9220 8188 9222
rect 7948 9200 8244 9220
rect 7760 9132 7880 9160
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7484 7670 7604 7698
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7484 6186 7512 7670
rect 7564 7472 7616 7478
rect 7760 7460 7788 8978
rect 7852 8974 7880 9132
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7616 7432 7788 7460
rect 7564 7414 7616 7420
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7484 5098 7512 6122
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7208 3454 7328 3482
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7208 2514 7236 3454
rect 7286 2544 7342 2553
rect 7196 2508 7248 2514
rect 7286 2479 7288 2488
rect 7196 2450 7248 2456
rect 7340 2479 7342 2488
rect 7288 2450 7340 2456
rect 7484 2446 7512 4762
rect 7576 4554 7604 7414
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 5302 7696 6734
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 6200 2204 6496 2224
rect 6256 2202 6280 2204
rect 6336 2202 6360 2204
rect 6416 2202 6440 2204
rect 6278 2150 6280 2202
rect 6342 2150 6354 2202
rect 6416 2150 6418 2202
rect 6256 2148 6280 2150
rect 6336 2148 6360 2150
rect 6416 2148 6440 2150
rect 6200 2128 6496 2148
rect 7576 2106 7604 3878
rect 7668 2582 7696 5238
rect 7760 3738 7788 7142
rect 7852 5914 7880 8502
rect 8036 8362 8064 8910
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7948 8188 8244 8208
rect 8004 8186 8028 8188
rect 8084 8186 8108 8188
rect 8164 8186 8188 8188
rect 8026 8134 8028 8186
rect 8090 8134 8102 8186
rect 8164 8134 8166 8186
rect 8004 8132 8028 8134
rect 8084 8132 8108 8134
rect 8164 8132 8188 8134
rect 7948 8112 8244 8132
rect 8114 7984 8170 7993
rect 8114 7919 8116 7928
rect 8168 7919 8170 7928
rect 8116 7890 8168 7896
rect 7948 7100 8244 7120
rect 8004 7098 8028 7100
rect 8084 7098 8108 7100
rect 8164 7098 8188 7100
rect 8026 7046 8028 7098
rect 8090 7046 8102 7098
rect 8164 7046 8166 7098
rect 8004 7044 8028 7046
rect 8084 7044 8108 7046
rect 8164 7044 8188 7046
rect 7948 7024 8244 7044
rect 7948 6012 8244 6032
rect 8004 6010 8028 6012
rect 8084 6010 8108 6012
rect 8164 6010 8188 6012
rect 8026 5958 8028 6010
rect 8090 5958 8102 6010
rect 8164 5958 8166 6010
rect 8004 5956 8028 5958
rect 8084 5956 8108 5958
rect 8164 5956 8188 5958
rect 7948 5936 8244 5956
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8312 5778 8340 10474
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9722 8432 9862
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 7852 5030 7880 5714
rect 8404 5710 8432 9658
rect 8496 8945 8524 11562
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10810 8616 10950
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8588 9722 8616 10066
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8482 8936 8538 8945
rect 8482 8871 8538 8880
rect 8680 7970 8708 11494
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8496 7942 8708 7970
rect 8496 7886 8524 7942
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 7002 8708 7278
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8772 5778 8800 10950
rect 8956 9178 8984 11562
rect 9140 9722 9168 14113
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9232 10606 9260 10746
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9324 10266 9352 13631
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9494 11248 9550 11257
rect 9494 11183 9550 11192
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9324 10130 9352 10202
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9416 10062 9444 10542
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9416 9450 9444 9862
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7760 3534 7788 3674
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7852 3194 7880 4966
rect 7948 4924 8244 4944
rect 8004 4922 8028 4924
rect 8084 4922 8108 4924
rect 8164 4922 8188 4924
rect 8026 4870 8028 4922
rect 8090 4870 8102 4922
rect 8164 4870 8166 4922
rect 8004 4868 8028 4870
rect 8084 4868 8108 4870
rect 8164 4868 8188 4870
rect 7948 4848 8244 4868
rect 8312 4706 8340 5034
rect 8220 4678 8340 4706
rect 8220 4146 8248 4678
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7948 3836 8244 3856
rect 8004 3834 8028 3836
rect 8084 3834 8108 3836
rect 8164 3834 8188 3836
rect 8026 3782 8028 3834
rect 8090 3782 8102 3834
rect 8164 3782 8166 3834
rect 8004 3780 8028 3782
rect 8084 3780 8108 3782
rect 8164 3780 8188 3782
rect 7948 3760 8244 3780
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 8312 3126 8340 4558
rect 8588 4282 8616 5102
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8588 3670 8616 3946
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8680 3074 8708 3538
rect 8772 3194 8800 5714
rect 8864 4758 8892 8298
rect 8956 7954 8984 9114
rect 9416 8566 9444 9386
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 8956 6458 8984 7278
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 9140 4078 9168 7278
rect 9324 7206 9352 8502
rect 9508 7546 9536 11183
rect 9600 8945 9628 12038
rect 9696 11996 9992 12016
rect 9752 11994 9776 11996
rect 9832 11994 9856 11996
rect 9912 11994 9936 11996
rect 9774 11942 9776 11994
rect 9838 11942 9850 11994
rect 9912 11942 9914 11994
rect 9752 11940 9776 11942
rect 9832 11940 9856 11942
rect 9912 11940 9936 11942
rect 9696 11920 9992 11940
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11354 9812 11698
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9696 10908 9992 10928
rect 9752 10906 9776 10908
rect 9832 10906 9856 10908
rect 9912 10906 9936 10908
rect 9774 10854 9776 10906
rect 9838 10854 9850 10906
rect 9912 10854 9914 10906
rect 9752 10852 9776 10854
rect 9832 10852 9856 10854
rect 9912 10852 9936 10854
rect 9696 10832 9992 10852
rect 10060 10674 10088 11154
rect 10612 11014 10640 14113
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9696 9820 9992 9840
rect 9752 9818 9776 9820
rect 9832 9818 9856 9820
rect 9912 9818 9936 9820
rect 9774 9766 9776 9818
rect 9838 9766 9850 9818
rect 9912 9766 9914 9818
rect 9752 9764 9776 9766
rect 9832 9764 9856 9766
rect 9912 9764 9936 9766
rect 9696 9744 9992 9764
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10060 9450 10088 9658
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9586 8936 9642 8945
rect 9586 8871 9642 8880
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9696 8732 9992 8752
rect 9752 8730 9776 8732
rect 9832 8730 9856 8732
rect 9912 8730 9936 8732
rect 9774 8678 9776 8730
rect 9838 8678 9850 8730
rect 9912 8678 9914 8730
rect 9752 8676 9776 8678
rect 9832 8676 9856 8678
rect 9912 8676 9936 8678
rect 9696 8656 9992 8676
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9692 7886 9720 8502
rect 10060 8430 10088 8842
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9696 7644 9992 7664
rect 9752 7642 9776 7644
rect 9832 7642 9856 7644
rect 9912 7642 9936 7644
rect 9774 7590 9776 7642
rect 9838 7590 9850 7642
rect 9912 7590 9914 7642
rect 9752 7588 9776 7590
rect 9832 7588 9856 7590
rect 9912 7588 9936 7590
rect 9696 7568 9992 7588
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8680 3046 8800 3074
rect 8772 2990 8800 3046
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8772 2854 8800 2926
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 7948 2748 8244 2768
rect 8004 2746 8028 2748
rect 8084 2746 8108 2748
rect 8164 2746 8188 2748
rect 8026 2694 8028 2746
rect 8090 2694 8102 2746
rect 8164 2694 8166 2746
rect 8004 2692 8028 2694
rect 8084 2692 8108 2694
rect 8164 2692 8188 2694
rect 7948 2672 8244 2692
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 8772 2514 8800 2790
rect 9048 2582 9076 2858
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 6104 1958 6316 1986
rect 6288 800 6316 1958
rect 7760 800 7788 2246
rect 9140 800 9168 2518
rect 9232 1329 9260 6190
rect 9324 5234 9352 7142
rect 9508 6254 9536 7482
rect 10152 6798 10180 10066
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 8498 10272 9318
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9696 6556 9992 6576
rect 9752 6554 9776 6556
rect 9832 6554 9856 6556
rect 9912 6554 9936 6556
rect 9774 6502 9776 6554
rect 9838 6502 9850 6554
rect 9912 6502 9914 6554
rect 9752 6500 9776 6502
rect 9832 6500 9856 6502
rect 9912 6500 9936 6502
rect 9696 6480 9992 6500
rect 10152 6322 10180 6734
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9876 5778 9904 6258
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10138 6216 10194 6225
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 10060 5574 10088 6190
rect 10138 6151 10194 6160
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9696 5468 9992 5488
rect 9752 5466 9776 5468
rect 9832 5466 9856 5468
rect 9912 5466 9936 5468
rect 9774 5414 9776 5466
rect 9838 5414 9850 5466
rect 9912 5414 9914 5466
rect 9752 5412 9776 5414
rect 9832 5412 9856 5414
rect 9912 5412 9936 5414
rect 9696 5392 9992 5412
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 4570 9720 4626
rect 9600 4542 9720 4570
rect 9600 4146 9628 4542
rect 9696 4380 9992 4400
rect 9752 4378 9776 4380
rect 9832 4378 9856 4380
rect 9912 4378 9936 4380
rect 9774 4326 9776 4378
rect 9838 4326 9850 4378
rect 9912 4326 9914 4378
rect 9752 4324 9776 4326
rect 9832 4324 9856 4326
rect 9912 4324 9936 4326
rect 9696 4304 9992 4324
rect 10060 4146 10088 5510
rect 10152 5166 10180 6151
rect 10244 5370 10272 6802
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10336 4758 10364 10678
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 8634 10456 9454
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9600 3777 9628 3946
rect 9586 3768 9642 3777
rect 10060 3738 10088 3946
rect 10428 3942 10456 7890
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 9586 3703 9642 3712
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 9696 3292 9992 3312
rect 9752 3290 9776 3292
rect 9832 3290 9856 3292
rect 9912 3290 9936 3292
rect 9774 3238 9776 3290
rect 9838 3238 9850 3290
rect 9912 3238 9914 3290
rect 9752 3236 9776 3238
rect 9832 3236 9856 3238
rect 9912 3236 9936 3238
rect 9696 3216 9992 3236
rect 10244 3194 10272 3606
rect 10520 3602 10548 10474
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10612 7478 10640 9998
rect 10704 8022 10732 12242
rect 11992 10538 12020 14113
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10704 6730 10732 7958
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10704 5098 10732 6666
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10152 2582 10180 3062
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 9696 2204 9992 2224
rect 9752 2202 9776 2204
rect 9832 2202 9856 2204
rect 9912 2202 9936 2204
rect 9774 2150 9776 2202
rect 9838 2150 9850 2202
rect 9912 2150 9914 2202
rect 9752 2148 9776 2150
rect 9832 2148 9856 2150
rect 9912 2148 9936 2150
rect 9696 2128 9992 2148
rect 9218 1320 9274 1329
rect 9218 1255 9274 1264
rect 10612 800 10640 2994
rect 10888 2514 10916 9386
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 11992 800 12020 2926
rect 662 0 718 800
rect 2042 0 2098 800
rect 3422 0 3478 800
rect 4894 0 4950 800
rect 6274 0 6330 800
rect 7746 0 7802 800
rect 9126 0 9182 800
rect 10598 0 10654 800
rect 11978 0 12034 800
<< via2 >>
rect 2704 11994 2760 11996
rect 2784 11994 2840 11996
rect 2864 11994 2920 11996
rect 2944 11994 3000 11996
rect 2704 11942 2730 11994
rect 2730 11942 2760 11994
rect 2784 11942 2794 11994
rect 2794 11942 2840 11994
rect 2864 11942 2910 11994
rect 2910 11942 2920 11994
rect 2944 11942 2974 11994
rect 2974 11942 3000 11994
rect 2704 11940 2760 11942
rect 2784 11940 2840 11942
rect 2864 11940 2920 11942
rect 2944 11940 3000 11942
rect 1858 11192 1914 11248
rect 2704 10906 2760 10908
rect 2784 10906 2840 10908
rect 2864 10906 2920 10908
rect 2944 10906 3000 10908
rect 2704 10854 2730 10906
rect 2730 10854 2760 10906
rect 2784 10854 2794 10906
rect 2794 10854 2840 10906
rect 2864 10854 2910 10906
rect 2910 10854 2920 10906
rect 2944 10854 2974 10906
rect 2974 10854 3000 10906
rect 2704 10852 2760 10854
rect 2784 10852 2840 10854
rect 2864 10852 2920 10854
rect 2944 10852 3000 10854
rect 1490 8744 1546 8800
rect 2704 9818 2760 9820
rect 2784 9818 2840 9820
rect 2864 9818 2920 9820
rect 2944 9818 3000 9820
rect 2704 9766 2730 9818
rect 2730 9766 2760 9818
rect 2784 9766 2794 9818
rect 2794 9766 2840 9818
rect 2864 9766 2910 9818
rect 2910 9766 2920 9818
rect 2944 9766 2974 9818
rect 2974 9766 3000 9818
rect 2704 9764 2760 9766
rect 2784 9764 2840 9766
rect 2864 9764 2920 9766
rect 2944 9764 3000 9766
rect 2870 8880 2926 8936
rect 2704 8730 2760 8732
rect 2784 8730 2840 8732
rect 2864 8730 2920 8732
rect 2944 8730 3000 8732
rect 2704 8678 2730 8730
rect 2730 8678 2760 8730
rect 2784 8678 2794 8730
rect 2794 8678 2840 8730
rect 2864 8678 2910 8730
rect 2910 8678 2920 8730
rect 2944 8678 2974 8730
rect 2974 8678 3000 8730
rect 2704 8676 2760 8678
rect 2784 8676 2840 8678
rect 2864 8676 2920 8678
rect 2944 8676 3000 8678
rect 2704 7642 2760 7644
rect 2784 7642 2840 7644
rect 2864 7642 2920 7644
rect 2944 7642 3000 7644
rect 2704 7590 2730 7642
rect 2730 7590 2760 7642
rect 2784 7590 2794 7642
rect 2794 7590 2840 7642
rect 2864 7590 2910 7642
rect 2910 7590 2920 7642
rect 2944 7590 2974 7642
rect 2974 7590 3000 7642
rect 2704 7588 2760 7590
rect 2784 7588 2840 7590
rect 2864 7588 2920 7590
rect 2944 7588 3000 7590
rect 2318 6160 2374 6216
rect 2704 6554 2760 6556
rect 2784 6554 2840 6556
rect 2864 6554 2920 6556
rect 2944 6554 3000 6556
rect 2704 6502 2730 6554
rect 2730 6502 2760 6554
rect 2784 6502 2794 6554
rect 2794 6502 2840 6554
rect 2864 6502 2910 6554
rect 2910 6502 2920 6554
rect 2944 6502 2974 6554
rect 2974 6502 3000 6554
rect 2704 6500 2760 6502
rect 2784 6500 2840 6502
rect 2864 6500 2920 6502
rect 2944 6500 3000 6502
rect 2704 5466 2760 5468
rect 2784 5466 2840 5468
rect 2864 5466 2920 5468
rect 2944 5466 3000 5468
rect 2704 5414 2730 5466
rect 2730 5414 2760 5466
rect 2784 5414 2794 5466
rect 2794 5414 2840 5466
rect 2864 5414 2910 5466
rect 2910 5414 2920 5466
rect 2944 5414 2974 5466
rect 2974 5414 3000 5466
rect 2704 5412 2760 5414
rect 2784 5412 2840 5414
rect 2864 5412 2920 5414
rect 2944 5412 3000 5414
rect 2704 4378 2760 4380
rect 2784 4378 2840 4380
rect 2864 4378 2920 4380
rect 2944 4378 3000 4380
rect 2704 4326 2730 4378
rect 2730 4326 2760 4378
rect 2784 4326 2794 4378
rect 2794 4326 2840 4378
rect 2864 4326 2910 4378
rect 2910 4326 2920 4378
rect 2944 4326 2974 4378
rect 2974 4326 3000 4378
rect 2704 4324 2760 4326
rect 2784 4324 2840 4326
rect 2864 4324 2920 4326
rect 2944 4324 3000 4326
rect 2704 3290 2760 3292
rect 2784 3290 2840 3292
rect 2864 3290 2920 3292
rect 2944 3290 3000 3292
rect 2704 3238 2730 3290
rect 2730 3238 2760 3290
rect 2784 3238 2794 3290
rect 2794 3238 2840 3290
rect 2864 3238 2910 3290
rect 2910 3238 2920 3290
rect 2944 3238 2974 3290
rect 2974 3238 3000 3290
rect 2704 3236 2760 3238
rect 2784 3236 2840 3238
rect 2864 3236 2920 3238
rect 2944 3236 3000 3238
rect 3606 13640 3662 13696
rect 4452 12538 4508 12540
rect 4532 12538 4588 12540
rect 4612 12538 4668 12540
rect 4692 12538 4748 12540
rect 4452 12486 4478 12538
rect 4478 12486 4508 12538
rect 4532 12486 4542 12538
rect 4542 12486 4588 12538
rect 4612 12486 4658 12538
rect 4658 12486 4668 12538
rect 4692 12486 4722 12538
rect 4722 12486 4748 12538
rect 4452 12484 4508 12486
rect 4532 12484 4588 12486
rect 4612 12484 4668 12486
rect 4692 12484 4748 12486
rect 3330 3712 3386 3768
rect 3054 2488 3110 2544
rect 2704 2202 2760 2204
rect 2784 2202 2840 2204
rect 2864 2202 2920 2204
rect 2944 2202 3000 2204
rect 2704 2150 2730 2202
rect 2730 2150 2760 2202
rect 2784 2150 2794 2202
rect 2794 2150 2840 2202
rect 2864 2150 2910 2202
rect 2910 2150 2920 2202
rect 2944 2150 2974 2202
rect 2974 2150 3000 2202
rect 2704 2148 2760 2150
rect 2784 2148 2840 2150
rect 2864 2148 2920 2150
rect 2944 2148 3000 2150
rect 2410 1264 2466 1320
rect 4452 11450 4508 11452
rect 4532 11450 4588 11452
rect 4612 11450 4668 11452
rect 4692 11450 4748 11452
rect 4452 11398 4478 11450
rect 4478 11398 4508 11450
rect 4532 11398 4542 11450
rect 4542 11398 4588 11450
rect 4612 11398 4658 11450
rect 4658 11398 4668 11450
rect 4692 11398 4722 11450
rect 4722 11398 4748 11450
rect 4452 11396 4508 11398
rect 4532 11396 4588 11398
rect 4612 11396 4668 11398
rect 4692 11396 4748 11398
rect 4452 10362 4508 10364
rect 4532 10362 4588 10364
rect 4612 10362 4668 10364
rect 4692 10362 4748 10364
rect 4452 10310 4478 10362
rect 4478 10310 4508 10362
rect 4532 10310 4542 10362
rect 4542 10310 4588 10362
rect 4612 10310 4658 10362
rect 4658 10310 4668 10362
rect 4692 10310 4722 10362
rect 4722 10310 4748 10362
rect 4452 10308 4508 10310
rect 4532 10308 4588 10310
rect 4612 10308 4668 10310
rect 4692 10308 4748 10310
rect 4452 9274 4508 9276
rect 4532 9274 4588 9276
rect 4612 9274 4668 9276
rect 4692 9274 4748 9276
rect 4452 9222 4478 9274
rect 4478 9222 4508 9274
rect 4532 9222 4542 9274
rect 4542 9222 4588 9274
rect 4612 9222 4658 9274
rect 4658 9222 4668 9274
rect 4692 9222 4722 9274
rect 4722 9222 4748 9274
rect 4452 9220 4508 9222
rect 4532 9220 4588 9222
rect 4612 9220 4668 9222
rect 4692 9220 4748 9222
rect 7948 12538 8004 12540
rect 8028 12538 8084 12540
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 7948 12486 7974 12538
rect 7974 12486 8004 12538
rect 8028 12486 8038 12538
rect 8038 12486 8084 12538
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8244 12538
rect 7948 12484 8004 12486
rect 8028 12484 8084 12486
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 6200 11994 6256 11996
rect 6280 11994 6336 11996
rect 6360 11994 6416 11996
rect 6440 11994 6496 11996
rect 6200 11942 6226 11994
rect 6226 11942 6256 11994
rect 6280 11942 6290 11994
rect 6290 11942 6336 11994
rect 6360 11942 6406 11994
rect 6406 11942 6416 11994
rect 6440 11942 6470 11994
rect 6470 11942 6496 11994
rect 6200 11940 6256 11942
rect 6280 11940 6336 11942
rect 6360 11940 6416 11942
rect 6440 11940 6496 11942
rect 6200 10906 6256 10908
rect 6280 10906 6336 10908
rect 6360 10906 6416 10908
rect 6440 10906 6496 10908
rect 6200 10854 6226 10906
rect 6226 10854 6256 10906
rect 6280 10854 6290 10906
rect 6290 10854 6336 10906
rect 6360 10854 6406 10906
rect 6406 10854 6416 10906
rect 6440 10854 6470 10906
rect 6470 10854 6496 10906
rect 6200 10852 6256 10854
rect 6280 10852 6336 10854
rect 6360 10852 6416 10854
rect 6440 10852 6496 10854
rect 4452 8186 4508 8188
rect 4532 8186 4588 8188
rect 4612 8186 4668 8188
rect 4692 8186 4748 8188
rect 4452 8134 4478 8186
rect 4478 8134 4508 8186
rect 4532 8134 4542 8186
rect 4542 8134 4588 8186
rect 4612 8134 4658 8186
rect 4658 8134 4668 8186
rect 4692 8134 4722 8186
rect 4722 8134 4748 8186
rect 4452 8132 4508 8134
rect 4532 8132 4588 8134
rect 4612 8132 4668 8134
rect 4692 8132 4748 8134
rect 4452 7098 4508 7100
rect 4532 7098 4588 7100
rect 4612 7098 4668 7100
rect 4692 7098 4748 7100
rect 4452 7046 4478 7098
rect 4478 7046 4508 7098
rect 4532 7046 4542 7098
rect 4542 7046 4588 7098
rect 4612 7046 4658 7098
rect 4658 7046 4668 7098
rect 4692 7046 4722 7098
rect 4722 7046 4748 7098
rect 4452 7044 4508 7046
rect 4532 7044 4588 7046
rect 4612 7044 4668 7046
rect 4692 7044 4748 7046
rect 4452 6010 4508 6012
rect 4532 6010 4588 6012
rect 4612 6010 4668 6012
rect 4692 6010 4748 6012
rect 4452 5958 4478 6010
rect 4478 5958 4508 6010
rect 4532 5958 4542 6010
rect 4542 5958 4588 6010
rect 4612 5958 4658 6010
rect 4658 5958 4668 6010
rect 4692 5958 4722 6010
rect 4722 5958 4748 6010
rect 4452 5956 4508 5958
rect 4532 5956 4588 5958
rect 4612 5956 4668 5958
rect 4692 5956 4748 5958
rect 4452 4922 4508 4924
rect 4532 4922 4588 4924
rect 4612 4922 4668 4924
rect 4692 4922 4748 4924
rect 4452 4870 4478 4922
rect 4478 4870 4508 4922
rect 4532 4870 4542 4922
rect 4542 4870 4588 4922
rect 4612 4870 4658 4922
rect 4658 4870 4668 4922
rect 4692 4870 4722 4922
rect 4722 4870 4748 4922
rect 4452 4868 4508 4870
rect 4532 4868 4588 4870
rect 4612 4868 4668 4870
rect 4692 4868 4748 4870
rect 4452 3834 4508 3836
rect 4532 3834 4588 3836
rect 4612 3834 4668 3836
rect 4692 3834 4748 3836
rect 4452 3782 4478 3834
rect 4478 3782 4508 3834
rect 4532 3782 4542 3834
rect 4542 3782 4588 3834
rect 4612 3782 4658 3834
rect 4658 3782 4668 3834
rect 4692 3782 4722 3834
rect 4722 3782 4748 3834
rect 4452 3780 4508 3782
rect 4532 3780 4588 3782
rect 4612 3780 4668 3782
rect 4692 3780 4748 3782
rect 4452 2746 4508 2748
rect 4532 2746 4588 2748
rect 4612 2746 4668 2748
rect 4692 2746 4748 2748
rect 4452 2694 4478 2746
rect 4478 2694 4508 2746
rect 4532 2694 4542 2746
rect 4542 2694 4588 2746
rect 4612 2694 4658 2746
rect 4658 2694 4668 2746
rect 4692 2694 4722 2746
rect 4722 2694 4748 2746
rect 4452 2692 4508 2694
rect 4532 2692 4588 2694
rect 4612 2692 4668 2694
rect 4692 2692 4748 2694
rect 6200 9818 6256 9820
rect 6280 9818 6336 9820
rect 6360 9818 6416 9820
rect 6440 9818 6496 9820
rect 6200 9766 6226 9818
rect 6226 9766 6256 9818
rect 6280 9766 6290 9818
rect 6290 9766 6336 9818
rect 6360 9766 6406 9818
rect 6406 9766 6416 9818
rect 6440 9766 6470 9818
rect 6470 9766 6496 9818
rect 6200 9764 6256 9766
rect 6280 9764 6336 9766
rect 6360 9764 6416 9766
rect 6440 9764 6496 9766
rect 6200 8730 6256 8732
rect 6280 8730 6336 8732
rect 6360 8730 6416 8732
rect 6440 8730 6496 8732
rect 6200 8678 6226 8730
rect 6226 8678 6256 8730
rect 6280 8678 6290 8730
rect 6290 8678 6336 8730
rect 6360 8678 6406 8730
rect 6406 8678 6416 8730
rect 6440 8678 6470 8730
rect 6470 8678 6496 8730
rect 6200 8676 6256 8678
rect 6280 8676 6336 8678
rect 6360 8676 6416 8678
rect 6440 8676 6496 8678
rect 6458 7948 6514 7984
rect 6458 7928 6460 7948
rect 6460 7928 6512 7948
rect 6512 7928 6514 7948
rect 6200 7642 6256 7644
rect 6280 7642 6336 7644
rect 6360 7642 6416 7644
rect 6440 7642 6496 7644
rect 6200 7590 6226 7642
rect 6226 7590 6256 7642
rect 6280 7590 6290 7642
rect 6290 7590 6336 7642
rect 6360 7590 6406 7642
rect 6406 7590 6416 7642
rect 6440 7590 6470 7642
rect 6470 7590 6496 7642
rect 6200 7588 6256 7590
rect 6280 7588 6336 7590
rect 6360 7588 6416 7590
rect 6440 7588 6496 7590
rect 6200 6554 6256 6556
rect 6280 6554 6336 6556
rect 6360 6554 6416 6556
rect 6440 6554 6496 6556
rect 6200 6502 6226 6554
rect 6226 6502 6256 6554
rect 6280 6502 6290 6554
rect 6290 6502 6336 6554
rect 6360 6502 6406 6554
rect 6406 6502 6416 6554
rect 6440 6502 6470 6554
rect 6470 6502 6496 6554
rect 6200 6500 6256 6502
rect 6280 6500 6336 6502
rect 6360 6500 6416 6502
rect 6440 6500 6496 6502
rect 6274 5616 6330 5672
rect 6200 5466 6256 5468
rect 6280 5466 6336 5468
rect 6360 5466 6416 5468
rect 6440 5466 6496 5468
rect 6200 5414 6226 5466
rect 6226 5414 6256 5466
rect 6280 5414 6290 5466
rect 6290 5414 6336 5466
rect 6360 5414 6406 5466
rect 6406 5414 6416 5466
rect 6440 5414 6470 5466
rect 6470 5414 6496 5466
rect 6200 5412 6256 5414
rect 6280 5412 6336 5414
rect 6360 5412 6416 5414
rect 6440 5412 6496 5414
rect 6200 4378 6256 4380
rect 6280 4378 6336 4380
rect 6360 4378 6416 4380
rect 6440 4378 6496 4380
rect 6200 4326 6226 4378
rect 6226 4326 6256 4378
rect 6280 4326 6290 4378
rect 6290 4326 6336 4378
rect 6360 4326 6406 4378
rect 6406 4326 6416 4378
rect 6440 4326 6470 4378
rect 6470 4326 6496 4378
rect 6200 4324 6256 4326
rect 6280 4324 6336 4326
rect 6360 4324 6416 4326
rect 6440 4324 6496 4326
rect 6200 3290 6256 3292
rect 6280 3290 6336 3292
rect 6360 3290 6416 3292
rect 6440 3290 6496 3292
rect 6200 3238 6226 3290
rect 6226 3238 6256 3290
rect 6280 3238 6290 3290
rect 6290 3238 6336 3290
rect 6360 3238 6406 3290
rect 6406 3238 6416 3290
rect 6440 3238 6470 3290
rect 6470 3238 6496 3290
rect 6200 3236 6256 3238
rect 6280 3236 6336 3238
rect 6360 3236 6416 3238
rect 6440 3236 6496 3238
rect 6826 8880 6882 8936
rect 6918 5208 6974 5264
rect 7948 11450 8004 11452
rect 8028 11450 8084 11452
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 7948 11398 7974 11450
rect 7974 11398 8004 11450
rect 8028 11398 8038 11450
rect 8038 11398 8084 11450
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8244 11450
rect 7948 11396 8004 11398
rect 8028 11396 8084 11398
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 7948 10362 8004 10364
rect 8028 10362 8084 10364
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 7948 10310 7974 10362
rect 7974 10310 8004 10362
rect 8028 10310 8038 10362
rect 8038 10310 8084 10362
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8244 10362
rect 7948 10308 8004 10310
rect 8028 10308 8084 10310
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 7948 9274 8004 9276
rect 8028 9274 8084 9276
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 7948 9222 7974 9274
rect 7974 9222 8004 9274
rect 8028 9222 8038 9274
rect 8038 9222 8084 9274
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8244 9274
rect 7948 9220 8004 9222
rect 8028 9220 8084 9222
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 7286 2508 7342 2544
rect 7286 2488 7288 2508
rect 7288 2488 7340 2508
rect 7340 2488 7342 2508
rect 6200 2202 6256 2204
rect 6280 2202 6336 2204
rect 6360 2202 6416 2204
rect 6440 2202 6496 2204
rect 6200 2150 6226 2202
rect 6226 2150 6256 2202
rect 6280 2150 6290 2202
rect 6290 2150 6336 2202
rect 6360 2150 6406 2202
rect 6406 2150 6416 2202
rect 6440 2150 6470 2202
rect 6470 2150 6496 2202
rect 6200 2148 6256 2150
rect 6280 2148 6336 2150
rect 6360 2148 6416 2150
rect 6440 2148 6496 2150
rect 7948 8186 8004 8188
rect 8028 8186 8084 8188
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 7948 8134 7974 8186
rect 7974 8134 8004 8186
rect 8028 8134 8038 8186
rect 8038 8134 8084 8186
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8244 8186
rect 7948 8132 8004 8134
rect 8028 8132 8084 8134
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8114 7948 8170 7984
rect 8114 7928 8116 7948
rect 8116 7928 8168 7948
rect 8168 7928 8170 7948
rect 7948 7098 8004 7100
rect 8028 7098 8084 7100
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 7948 7046 7974 7098
rect 7974 7046 8004 7098
rect 8028 7046 8038 7098
rect 8038 7046 8084 7098
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8244 7098
rect 7948 7044 8004 7046
rect 8028 7044 8084 7046
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 7948 6010 8004 6012
rect 8028 6010 8084 6012
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 7948 5958 7974 6010
rect 7974 5958 8004 6010
rect 8028 5958 8038 6010
rect 8038 5958 8084 6010
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8244 6010
rect 7948 5956 8004 5958
rect 8028 5956 8084 5958
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8482 8880 8538 8936
rect 9310 13640 9366 13696
rect 9494 11192 9550 11248
rect 7948 4922 8004 4924
rect 8028 4922 8084 4924
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 7948 4870 7974 4922
rect 7974 4870 8004 4922
rect 8028 4870 8038 4922
rect 8038 4870 8084 4922
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8244 4922
rect 7948 4868 8004 4870
rect 8028 4868 8084 4870
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 7948 3834 8004 3836
rect 8028 3834 8084 3836
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 7948 3782 7974 3834
rect 7974 3782 8004 3834
rect 8028 3782 8038 3834
rect 8038 3782 8084 3834
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8244 3834
rect 7948 3780 8004 3782
rect 8028 3780 8084 3782
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 9696 11994 9752 11996
rect 9776 11994 9832 11996
rect 9856 11994 9912 11996
rect 9936 11994 9992 11996
rect 9696 11942 9722 11994
rect 9722 11942 9752 11994
rect 9776 11942 9786 11994
rect 9786 11942 9832 11994
rect 9856 11942 9902 11994
rect 9902 11942 9912 11994
rect 9936 11942 9966 11994
rect 9966 11942 9992 11994
rect 9696 11940 9752 11942
rect 9776 11940 9832 11942
rect 9856 11940 9912 11942
rect 9936 11940 9992 11942
rect 9696 10906 9752 10908
rect 9776 10906 9832 10908
rect 9856 10906 9912 10908
rect 9936 10906 9992 10908
rect 9696 10854 9722 10906
rect 9722 10854 9752 10906
rect 9776 10854 9786 10906
rect 9786 10854 9832 10906
rect 9856 10854 9902 10906
rect 9902 10854 9912 10906
rect 9936 10854 9966 10906
rect 9966 10854 9992 10906
rect 9696 10852 9752 10854
rect 9776 10852 9832 10854
rect 9856 10852 9912 10854
rect 9936 10852 9992 10854
rect 9696 9818 9752 9820
rect 9776 9818 9832 9820
rect 9856 9818 9912 9820
rect 9936 9818 9992 9820
rect 9696 9766 9722 9818
rect 9722 9766 9752 9818
rect 9776 9766 9786 9818
rect 9786 9766 9832 9818
rect 9856 9766 9902 9818
rect 9902 9766 9912 9818
rect 9936 9766 9966 9818
rect 9966 9766 9992 9818
rect 9696 9764 9752 9766
rect 9776 9764 9832 9766
rect 9856 9764 9912 9766
rect 9936 9764 9992 9766
rect 9586 8880 9642 8936
rect 9696 8730 9752 8732
rect 9776 8730 9832 8732
rect 9856 8730 9912 8732
rect 9936 8730 9992 8732
rect 9696 8678 9722 8730
rect 9722 8678 9752 8730
rect 9776 8678 9786 8730
rect 9786 8678 9832 8730
rect 9856 8678 9902 8730
rect 9902 8678 9912 8730
rect 9936 8678 9966 8730
rect 9966 8678 9992 8730
rect 9696 8676 9752 8678
rect 9776 8676 9832 8678
rect 9856 8676 9912 8678
rect 9936 8676 9992 8678
rect 9696 7642 9752 7644
rect 9776 7642 9832 7644
rect 9856 7642 9912 7644
rect 9936 7642 9992 7644
rect 9696 7590 9722 7642
rect 9722 7590 9752 7642
rect 9776 7590 9786 7642
rect 9786 7590 9832 7642
rect 9856 7590 9902 7642
rect 9902 7590 9912 7642
rect 9936 7590 9966 7642
rect 9966 7590 9992 7642
rect 9696 7588 9752 7590
rect 9776 7588 9832 7590
rect 9856 7588 9912 7590
rect 9936 7588 9992 7590
rect 7948 2746 8004 2748
rect 8028 2746 8084 2748
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 7948 2694 7974 2746
rect 7974 2694 8004 2746
rect 8028 2694 8038 2746
rect 8038 2694 8084 2746
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8244 2746
rect 7948 2692 8004 2694
rect 8028 2692 8084 2694
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 9696 6554 9752 6556
rect 9776 6554 9832 6556
rect 9856 6554 9912 6556
rect 9936 6554 9992 6556
rect 9696 6502 9722 6554
rect 9722 6502 9752 6554
rect 9776 6502 9786 6554
rect 9786 6502 9832 6554
rect 9856 6502 9902 6554
rect 9902 6502 9912 6554
rect 9936 6502 9966 6554
rect 9966 6502 9992 6554
rect 9696 6500 9752 6502
rect 9776 6500 9832 6502
rect 9856 6500 9912 6502
rect 9936 6500 9992 6502
rect 10138 6160 10194 6216
rect 9696 5466 9752 5468
rect 9776 5466 9832 5468
rect 9856 5466 9912 5468
rect 9936 5466 9992 5468
rect 9696 5414 9722 5466
rect 9722 5414 9752 5466
rect 9776 5414 9786 5466
rect 9786 5414 9832 5466
rect 9856 5414 9902 5466
rect 9902 5414 9912 5466
rect 9936 5414 9966 5466
rect 9966 5414 9992 5466
rect 9696 5412 9752 5414
rect 9776 5412 9832 5414
rect 9856 5412 9912 5414
rect 9936 5412 9992 5414
rect 9696 4378 9752 4380
rect 9776 4378 9832 4380
rect 9856 4378 9912 4380
rect 9936 4378 9992 4380
rect 9696 4326 9722 4378
rect 9722 4326 9752 4378
rect 9776 4326 9786 4378
rect 9786 4326 9832 4378
rect 9856 4326 9902 4378
rect 9902 4326 9912 4378
rect 9936 4326 9966 4378
rect 9966 4326 9992 4378
rect 9696 4324 9752 4326
rect 9776 4324 9832 4326
rect 9856 4324 9912 4326
rect 9936 4324 9992 4326
rect 9586 3712 9642 3768
rect 9696 3290 9752 3292
rect 9776 3290 9832 3292
rect 9856 3290 9912 3292
rect 9936 3290 9992 3292
rect 9696 3238 9722 3290
rect 9722 3238 9752 3290
rect 9776 3238 9786 3290
rect 9786 3238 9832 3290
rect 9856 3238 9902 3290
rect 9902 3238 9912 3290
rect 9936 3238 9966 3290
rect 9966 3238 9992 3290
rect 9696 3236 9752 3238
rect 9776 3236 9832 3238
rect 9856 3236 9912 3238
rect 9936 3236 9992 3238
rect 9696 2202 9752 2204
rect 9776 2202 9832 2204
rect 9856 2202 9912 2204
rect 9936 2202 9992 2204
rect 9696 2150 9722 2202
rect 9722 2150 9752 2202
rect 9776 2150 9786 2202
rect 9786 2150 9832 2202
rect 9856 2150 9902 2202
rect 9902 2150 9912 2202
rect 9936 2150 9966 2202
rect 9966 2150 9992 2202
rect 9696 2148 9752 2150
rect 9776 2148 9832 2150
rect 9856 2148 9912 2150
rect 9936 2148 9992 2150
rect 9218 1264 9274 1320
<< metal3 >>
rect 0 13698 800 13728
rect 3601 13698 3667 13701
rect 0 13696 3667 13698
rect 0 13640 3606 13696
rect 3662 13640 3667 13696
rect 0 13638 3667 13640
rect 0 13608 800 13638
rect 3601 13635 3667 13638
rect 9305 13698 9371 13701
rect 11969 13698 12769 13728
rect 9305 13696 12769 13698
rect 9305 13640 9310 13696
rect 9366 13640 12769 13696
rect 9305 13638 12769 13640
rect 9305 13635 9371 13638
rect 11969 13608 12769 13638
rect 4440 12544 4760 12545
rect 4440 12480 4448 12544
rect 4512 12480 4528 12544
rect 4592 12480 4608 12544
rect 4672 12480 4688 12544
rect 4752 12480 4760 12544
rect 4440 12479 4760 12480
rect 7936 12544 8256 12545
rect 7936 12480 7944 12544
rect 8008 12480 8024 12544
rect 8088 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8256 12544
rect 7936 12479 8256 12480
rect 2692 12000 3012 12001
rect 2692 11936 2700 12000
rect 2764 11936 2780 12000
rect 2844 11936 2860 12000
rect 2924 11936 2940 12000
rect 3004 11936 3012 12000
rect 2692 11935 3012 11936
rect 6188 12000 6508 12001
rect 6188 11936 6196 12000
rect 6260 11936 6276 12000
rect 6340 11936 6356 12000
rect 6420 11936 6436 12000
rect 6500 11936 6508 12000
rect 6188 11935 6508 11936
rect 9684 12000 10004 12001
rect 9684 11936 9692 12000
rect 9756 11936 9772 12000
rect 9836 11936 9852 12000
rect 9916 11936 9932 12000
rect 9996 11936 10004 12000
rect 9684 11935 10004 11936
rect 4440 11456 4760 11457
rect 4440 11392 4448 11456
rect 4512 11392 4528 11456
rect 4592 11392 4608 11456
rect 4672 11392 4688 11456
rect 4752 11392 4760 11456
rect 4440 11391 4760 11392
rect 7936 11456 8256 11457
rect 7936 11392 7944 11456
rect 8008 11392 8024 11456
rect 8088 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8256 11456
rect 7936 11391 8256 11392
rect 0 11250 800 11280
rect 1853 11250 1919 11253
rect 0 11248 1919 11250
rect 0 11192 1858 11248
rect 1914 11192 1919 11248
rect 0 11190 1919 11192
rect 0 11160 800 11190
rect 1853 11187 1919 11190
rect 9489 11250 9555 11253
rect 11969 11250 12769 11280
rect 9489 11248 12769 11250
rect 9489 11192 9494 11248
rect 9550 11192 12769 11248
rect 9489 11190 12769 11192
rect 9489 11187 9555 11190
rect 11969 11160 12769 11190
rect 2692 10912 3012 10913
rect 2692 10848 2700 10912
rect 2764 10848 2780 10912
rect 2844 10848 2860 10912
rect 2924 10848 2940 10912
rect 3004 10848 3012 10912
rect 2692 10847 3012 10848
rect 6188 10912 6508 10913
rect 6188 10848 6196 10912
rect 6260 10848 6276 10912
rect 6340 10848 6356 10912
rect 6420 10848 6436 10912
rect 6500 10848 6508 10912
rect 6188 10847 6508 10848
rect 9684 10912 10004 10913
rect 9684 10848 9692 10912
rect 9756 10848 9772 10912
rect 9836 10848 9852 10912
rect 9916 10848 9932 10912
rect 9996 10848 10004 10912
rect 9684 10847 10004 10848
rect 4440 10368 4760 10369
rect 4440 10304 4448 10368
rect 4512 10304 4528 10368
rect 4592 10304 4608 10368
rect 4672 10304 4688 10368
rect 4752 10304 4760 10368
rect 4440 10303 4760 10304
rect 7936 10368 8256 10369
rect 7936 10304 7944 10368
rect 8008 10304 8024 10368
rect 8088 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8256 10368
rect 7936 10303 8256 10304
rect 2692 9824 3012 9825
rect 2692 9760 2700 9824
rect 2764 9760 2780 9824
rect 2844 9760 2860 9824
rect 2924 9760 2940 9824
rect 3004 9760 3012 9824
rect 2692 9759 3012 9760
rect 6188 9824 6508 9825
rect 6188 9760 6196 9824
rect 6260 9760 6276 9824
rect 6340 9760 6356 9824
rect 6420 9760 6436 9824
rect 6500 9760 6508 9824
rect 6188 9759 6508 9760
rect 9684 9824 10004 9825
rect 9684 9760 9692 9824
rect 9756 9760 9772 9824
rect 9836 9760 9852 9824
rect 9916 9760 9932 9824
rect 9996 9760 10004 9824
rect 9684 9759 10004 9760
rect 4440 9280 4760 9281
rect 4440 9216 4448 9280
rect 4512 9216 4528 9280
rect 4592 9216 4608 9280
rect 4672 9216 4688 9280
rect 4752 9216 4760 9280
rect 4440 9215 4760 9216
rect 7936 9280 8256 9281
rect 7936 9216 7944 9280
rect 8008 9216 8024 9280
rect 8088 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8256 9280
rect 7936 9215 8256 9216
rect 2865 8938 2931 8941
rect 6821 8938 6887 8941
rect 8477 8938 8543 8941
rect 2865 8936 8543 8938
rect 2865 8880 2870 8936
rect 2926 8880 6826 8936
rect 6882 8880 8482 8936
rect 8538 8880 8543 8936
rect 2865 8878 8543 8880
rect 2865 8875 2931 8878
rect 6821 8875 6887 8878
rect 8477 8875 8543 8878
rect 9581 8938 9647 8941
rect 9581 8936 10242 8938
rect 9581 8880 9586 8936
rect 9642 8880 10242 8936
rect 9581 8878 10242 8880
rect 9581 8875 9647 8878
rect 0 8802 800 8832
rect 1485 8802 1551 8805
rect 0 8800 1551 8802
rect 0 8744 1490 8800
rect 1546 8744 1551 8800
rect 0 8742 1551 8744
rect 10182 8802 10242 8878
rect 11969 8802 12769 8832
rect 10182 8742 12769 8802
rect 0 8712 800 8742
rect 1485 8739 1551 8742
rect 2692 8736 3012 8737
rect 2692 8672 2700 8736
rect 2764 8672 2780 8736
rect 2844 8672 2860 8736
rect 2924 8672 2940 8736
rect 3004 8672 3012 8736
rect 2692 8671 3012 8672
rect 6188 8736 6508 8737
rect 6188 8672 6196 8736
rect 6260 8672 6276 8736
rect 6340 8672 6356 8736
rect 6420 8672 6436 8736
rect 6500 8672 6508 8736
rect 6188 8671 6508 8672
rect 9684 8736 10004 8737
rect 9684 8672 9692 8736
rect 9756 8672 9772 8736
rect 9836 8672 9852 8736
rect 9916 8672 9932 8736
rect 9996 8672 10004 8736
rect 11969 8712 12769 8742
rect 9684 8671 10004 8672
rect 4440 8192 4760 8193
rect 4440 8128 4448 8192
rect 4512 8128 4528 8192
rect 4592 8128 4608 8192
rect 4672 8128 4688 8192
rect 4752 8128 4760 8192
rect 4440 8127 4760 8128
rect 7936 8192 8256 8193
rect 7936 8128 7944 8192
rect 8008 8128 8024 8192
rect 8088 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8256 8192
rect 7936 8127 8256 8128
rect 6453 7986 6519 7989
rect 8109 7986 8175 7989
rect 6453 7984 8175 7986
rect 6453 7928 6458 7984
rect 6514 7928 8114 7984
rect 8170 7928 8175 7984
rect 6453 7926 8175 7928
rect 6453 7923 6519 7926
rect 8109 7923 8175 7926
rect 2692 7648 3012 7649
rect 2692 7584 2700 7648
rect 2764 7584 2780 7648
rect 2844 7584 2860 7648
rect 2924 7584 2940 7648
rect 3004 7584 3012 7648
rect 2692 7583 3012 7584
rect 6188 7648 6508 7649
rect 6188 7584 6196 7648
rect 6260 7584 6276 7648
rect 6340 7584 6356 7648
rect 6420 7584 6436 7648
rect 6500 7584 6508 7648
rect 6188 7583 6508 7584
rect 9684 7648 10004 7649
rect 9684 7584 9692 7648
rect 9756 7584 9772 7648
rect 9836 7584 9852 7648
rect 9916 7584 9932 7648
rect 9996 7584 10004 7648
rect 9684 7583 10004 7584
rect 4440 7104 4760 7105
rect 4440 7040 4448 7104
rect 4512 7040 4528 7104
rect 4592 7040 4608 7104
rect 4672 7040 4688 7104
rect 4752 7040 4760 7104
rect 4440 7039 4760 7040
rect 7936 7104 8256 7105
rect 7936 7040 7944 7104
rect 8008 7040 8024 7104
rect 8088 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8256 7104
rect 7936 7039 8256 7040
rect 2692 6560 3012 6561
rect 2692 6496 2700 6560
rect 2764 6496 2780 6560
rect 2844 6496 2860 6560
rect 2924 6496 2940 6560
rect 3004 6496 3012 6560
rect 2692 6495 3012 6496
rect 6188 6560 6508 6561
rect 6188 6496 6196 6560
rect 6260 6496 6276 6560
rect 6340 6496 6356 6560
rect 6420 6496 6436 6560
rect 6500 6496 6508 6560
rect 6188 6495 6508 6496
rect 9684 6560 10004 6561
rect 9684 6496 9692 6560
rect 9756 6496 9772 6560
rect 9836 6496 9852 6560
rect 9916 6496 9932 6560
rect 9996 6496 10004 6560
rect 9684 6495 10004 6496
rect 0 6218 800 6248
rect 2313 6218 2379 6221
rect 0 6216 2379 6218
rect 0 6160 2318 6216
rect 2374 6160 2379 6216
rect 0 6158 2379 6160
rect 0 6128 800 6158
rect 2313 6155 2379 6158
rect 10133 6218 10199 6221
rect 11969 6218 12769 6248
rect 10133 6216 12769 6218
rect 10133 6160 10138 6216
rect 10194 6160 12769 6216
rect 10133 6158 12769 6160
rect 10133 6155 10199 6158
rect 11969 6128 12769 6158
rect 4440 6016 4760 6017
rect 4440 5952 4448 6016
rect 4512 5952 4528 6016
rect 4592 5952 4608 6016
rect 4672 5952 4688 6016
rect 4752 5952 4760 6016
rect 4440 5951 4760 5952
rect 7936 6016 8256 6017
rect 7936 5952 7944 6016
rect 8008 5952 8024 6016
rect 8088 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8256 6016
rect 7936 5951 8256 5952
rect 6269 5674 6335 5677
rect 6269 5672 6930 5674
rect 6269 5616 6274 5672
rect 6330 5616 6930 5672
rect 6269 5614 6930 5616
rect 6269 5611 6335 5614
rect 2692 5472 3012 5473
rect 2692 5408 2700 5472
rect 2764 5408 2780 5472
rect 2844 5408 2860 5472
rect 2924 5408 2940 5472
rect 3004 5408 3012 5472
rect 2692 5407 3012 5408
rect 6188 5472 6508 5473
rect 6188 5408 6196 5472
rect 6260 5408 6276 5472
rect 6340 5408 6356 5472
rect 6420 5408 6436 5472
rect 6500 5408 6508 5472
rect 6188 5407 6508 5408
rect 6870 5269 6930 5614
rect 9684 5472 10004 5473
rect 9684 5408 9692 5472
rect 9756 5408 9772 5472
rect 9836 5408 9852 5472
rect 9916 5408 9932 5472
rect 9996 5408 10004 5472
rect 9684 5407 10004 5408
rect 6870 5264 6979 5269
rect 6870 5208 6918 5264
rect 6974 5208 6979 5264
rect 6870 5206 6979 5208
rect 6913 5203 6979 5206
rect 4440 4928 4760 4929
rect 4440 4864 4448 4928
rect 4512 4864 4528 4928
rect 4592 4864 4608 4928
rect 4672 4864 4688 4928
rect 4752 4864 4760 4928
rect 4440 4863 4760 4864
rect 7936 4928 8256 4929
rect 7936 4864 7944 4928
rect 8008 4864 8024 4928
rect 8088 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8256 4928
rect 7936 4863 8256 4864
rect 2692 4384 3012 4385
rect 2692 4320 2700 4384
rect 2764 4320 2780 4384
rect 2844 4320 2860 4384
rect 2924 4320 2940 4384
rect 3004 4320 3012 4384
rect 2692 4319 3012 4320
rect 6188 4384 6508 4385
rect 6188 4320 6196 4384
rect 6260 4320 6276 4384
rect 6340 4320 6356 4384
rect 6420 4320 6436 4384
rect 6500 4320 6508 4384
rect 6188 4319 6508 4320
rect 9684 4384 10004 4385
rect 9684 4320 9692 4384
rect 9756 4320 9772 4384
rect 9836 4320 9852 4384
rect 9916 4320 9932 4384
rect 9996 4320 10004 4384
rect 9684 4319 10004 4320
rect 4440 3840 4760 3841
rect 0 3770 800 3800
rect 4440 3776 4448 3840
rect 4512 3776 4528 3840
rect 4592 3776 4608 3840
rect 4672 3776 4688 3840
rect 4752 3776 4760 3840
rect 4440 3775 4760 3776
rect 7936 3840 8256 3841
rect 7936 3776 7944 3840
rect 8008 3776 8024 3840
rect 8088 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8256 3840
rect 7936 3775 8256 3776
rect 3325 3770 3391 3773
rect 0 3768 3391 3770
rect 0 3712 3330 3768
rect 3386 3712 3391 3768
rect 0 3710 3391 3712
rect 0 3680 800 3710
rect 3325 3707 3391 3710
rect 9581 3770 9647 3773
rect 11969 3770 12769 3800
rect 9581 3768 12769 3770
rect 9581 3712 9586 3768
rect 9642 3712 12769 3768
rect 9581 3710 12769 3712
rect 9581 3707 9647 3710
rect 11969 3680 12769 3710
rect 2692 3296 3012 3297
rect 2692 3232 2700 3296
rect 2764 3232 2780 3296
rect 2844 3232 2860 3296
rect 2924 3232 2940 3296
rect 3004 3232 3012 3296
rect 2692 3231 3012 3232
rect 6188 3296 6508 3297
rect 6188 3232 6196 3296
rect 6260 3232 6276 3296
rect 6340 3232 6356 3296
rect 6420 3232 6436 3296
rect 6500 3232 6508 3296
rect 6188 3231 6508 3232
rect 9684 3296 10004 3297
rect 9684 3232 9692 3296
rect 9756 3232 9772 3296
rect 9836 3232 9852 3296
rect 9916 3232 9932 3296
rect 9996 3232 10004 3296
rect 9684 3231 10004 3232
rect 4440 2752 4760 2753
rect 4440 2688 4448 2752
rect 4512 2688 4528 2752
rect 4592 2688 4608 2752
rect 4672 2688 4688 2752
rect 4752 2688 4760 2752
rect 4440 2687 4760 2688
rect 7936 2752 8256 2753
rect 7936 2688 7944 2752
rect 8008 2688 8024 2752
rect 8088 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8256 2752
rect 7936 2687 8256 2688
rect 3049 2546 3115 2549
rect 7281 2546 7347 2549
rect 3049 2544 7347 2546
rect 3049 2488 3054 2544
rect 3110 2488 7286 2544
rect 7342 2488 7347 2544
rect 3049 2486 7347 2488
rect 3049 2483 3115 2486
rect 7281 2483 7347 2486
rect 2692 2208 3012 2209
rect 2692 2144 2700 2208
rect 2764 2144 2780 2208
rect 2844 2144 2860 2208
rect 2924 2144 2940 2208
rect 3004 2144 3012 2208
rect 2692 2143 3012 2144
rect 6188 2208 6508 2209
rect 6188 2144 6196 2208
rect 6260 2144 6276 2208
rect 6340 2144 6356 2208
rect 6420 2144 6436 2208
rect 6500 2144 6508 2208
rect 6188 2143 6508 2144
rect 9684 2208 10004 2209
rect 9684 2144 9692 2208
rect 9756 2144 9772 2208
rect 9836 2144 9852 2208
rect 9916 2144 9932 2208
rect 9996 2144 10004 2208
rect 9684 2143 10004 2144
rect 0 1322 800 1352
rect 2405 1322 2471 1325
rect 0 1320 2471 1322
rect 0 1264 2410 1320
rect 2466 1264 2471 1320
rect 0 1262 2471 1264
rect 0 1232 800 1262
rect 2405 1259 2471 1262
rect 9213 1322 9279 1325
rect 11969 1322 12769 1352
rect 9213 1320 12769 1322
rect 9213 1264 9218 1320
rect 9274 1264 12769 1320
rect 9213 1262 12769 1264
rect 9213 1259 9279 1262
rect 11969 1232 12769 1262
<< via3 >>
rect 4448 12540 4512 12544
rect 4448 12484 4452 12540
rect 4452 12484 4508 12540
rect 4508 12484 4512 12540
rect 4448 12480 4512 12484
rect 4528 12540 4592 12544
rect 4528 12484 4532 12540
rect 4532 12484 4588 12540
rect 4588 12484 4592 12540
rect 4528 12480 4592 12484
rect 4608 12540 4672 12544
rect 4608 12484 4612 12540
rect 4612 12484 4668 12540
rect 4668 12484 4672 12540
rect 4608 12480 4672 12484
rect 4688 12540 4752 12544
rect 4688 12484 4692 12540
rect 4692 12484 4748 12540
rect 4748 12484 4752 12540
rect 4688 12480 4752 12484
rect 7944 12540 8008 12544
rect 7944 12484 7948 12540
rect 7948 12484 8004 12540
rect 8004 12484 8008 12540
rect 7944 12480 8008 12484
rect 8024 12540 8088 12544
rect 8024 12484 8028 12540
rect 8028 12484 8084 12540
rect 8084 12484 8088 12540
rect 8024 12480 8088 12484
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 2700 11996 2764 12000
rect 2700 11940 2704 11996
rect 2704 11940 2760 11996
rect 2760 11940 2764 11996
rect 2700 11936 2764 11940
rect 2780 11996 2844 12000
rect 2780 11940 2784 11996
rect 2784 11940 2840 11996
rect 2840 11940 2844 11996
rect 2780 11936 2844 11940
rect 2860 11996 2924 12000
rect 2860 11940 2864 11996
rect 2864 11940 2920 11996
rect 2920 11940 2924 11996
rect 2860 11936 2924 11940
rect 2940 11996 3004 12000
rect 2940 11940 2944 11996
rect 2944 11940 3000 11996
rect 3000 11940 3004 11996
rect 2940 11936 3004 11940
rect 6196 11996 6260 12000
rect 6196 11940 6200 11996
rect 6200 11940 6256 11996
rect 6256 11940 6260 11996
rect 6196 11936 6260 11940
rect 6276 11996 6340 12000
rect 6276 11940 6280 11996
rect 6280 11940 6336 11996
rect 6336 11940 6340 11996
rect 6276 11936 6340 11940
rect 6356 11996 6420 12000
rect 6356 11940 6360 11996
rect 6360 11940 6416 11996
rect 6416 11940 6420 11996
rect 6356 11936 6420 11940
rect 6436 11996 6500 12000
rect 6436 11940 6440 11996
rect 6440 11940 6496 11996
rect 6496 11940 6500 11996
rect 6436 11936 6500 11940
rect 9692 11996 9756 12000
rect 9692 11940 9696 11996
rect 9696 11940 9752 11996
rect 9752 11940 9756 11996
rect 9692 11936 9756 11940
rect 9772 11996 9836 12000
rect 9772 11940 9776 11996
rect 9776 11940 9832 11996
rect 9832 11940 9836 11996
rect 9772 11936 9836 11940
rect 9852 11996 9916 12000
rect 9852 11940 9856 11996
rect 9856 11940 9912 11996
rect 9912 11940 9916 11996
rect 9852 11936 9916 11940
rect 9932 11996 9996 12000
rect 9932 11940 9936 11996
rect 9936 11940 9992 11996
rect 9992 11940 9996 11996
rect 9932 11936 9996 11940
rect 4448 11452 4512 11456
rect 4448 11396 4452 11452
rect 4452 11396 4508 11452
rect 4508 11396 4512 11452
rect 4448 11392 4512 11396
rect 4528 11452 4592 11456
rect 4528 11396 4532 11452
rect 4532 11396 4588 11452
rect 4588 11396 4592 11452
rect 4528 11392 4592 11396
rect 4608 11452 4672 11456
rect 4608 11396 4612 11452
rect 4612 11396 4668 11452
rect 4668 11396 4672 11452
rect 4608 11392 4672 11396
rect 4688 11452 4752 11456
rect 4688 11396 4692 11452
rect 4692 11396 4748 11452
rect 4748 11396 4752 11452
rect 4688 11392 4752 11396
rect 7944 11452 8008 11456
rect 7944 11396 7948 11452
rect 7948 11396 8004 11452
rect 8004 11396 8008 11452
rect 7944 11392 8008 11396
rect 8024 11452 8088 11456
rect 8024 11396 8028 11452
rect 8028 11396 8084 11452
rect 8084 11396 8088 11452
rect 8024 11392 8088 11396
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 2700 10908 2764 10912
rect 2700 10852 2704 10908
rect 2704 10852 2760 10908
rect 2760 10852 2764 10908
rect 2700 10848 2764 10852
rect 2780 10908 2844 10912
rect 2780 10852 2784 10908
rect 2784 10852 2840 10908
rect 2840 10852 2844 10908
rect 2780 10848 2844 10852
rect 2860 10908 2924 10912
rect 2860 10852 2864 10908
rect 2864 10852 2920 10908
rect 2920 10852 2924 10908
rect 2860 10848 2924 10852
rect 2940 10908 3004 10912
rect 2940 10852 2944 10908
rect 2944 10852 3000 10908
rect 3000 10852 3004 10908
rect 2940 10848 3004 10852
rect 6196 10908 6260 10912
rect 6196 10852 6200 10908
rect 6200 10852 6256 10908
rect 6256 10852 6260 10908
rect 6196 10848 6260 10852
rect 6276 10908 6340 10912
rect 6276 10852 6280 10908
rect 6280 10852 6336 10908
rect 6336 10852 6340 10908
rect 6276 10848 6340 10852
rect 6356 10908 6420 10912
rect 6356 10852 6360 10908
rect 6360 10852 6416 10908
rect 6416 10852 6420 10908
rect 6356 10848 6420 10852
rect 6436 10908 6500 10912
rect 6436 10852 6440 10908
rect 6440 10852 6496 10908
rect 6496 10852 6500 10908
rect 6436 10848 6500 10852
rect 9692 10908 9756 10912
rect 9692 10852 9696 10908
rect 9696 10852 9752 10908
rect 9752 10852 9756 10908
rect 9692 10848 9756 10852
rect 9772 10908 9836 10912
rect 9772 10852 9776 10908
rect 9776 10852 9832 10908
rect 9832 10852 9836 10908
rect 9772 10848 9836 10852
rect 9852 10908 9916 10912
rect 9852 10852 9856 10908
rect 9856 10852 9912 10908
rect 9912 10852 9916 10908
rect 9852 10848 9916 10852
rect 9932 10908 9996 10912
rect 9932 10852 9936 10908
rect 9936 10852 9992 10908
rect 9992 10852 9996 10908
rect 9932 10848 9996 10852
rect 4448 10364 4512 10368
rect 4448 10308 4452 10364
rect 4452 10308 4508 10364
rect 4508 10308 4512 10364
rect 4448 10304 4512 10308
rect 4528 10364 4592 10368
rect 4528 10308 4532 10364
rect 4532 10308 4588 10364
rect 4588 10308 4592 10364
rect 4528 10304 4592 10308
rect 4608 10364 4672 10368
rect 4608 10308 4612 10364
rect 4612 10308 4668 10364
rect 4668 10308 4672 10364
rect 4608 10304 4672 10308
rect 4688 10364 4752 10368
rect 4688 10308 4692 10364
rect 4692 10308 4748 10364
rect 4748 10308 4752 10364
rect 4688 10304 4752 10308
rect 7944 10364 8008 10368
rect 7944 10308 7948 10364
rect 7948 10308 8004 10364
rect 8004 10308 8008 10364
rect 7944 10304 8008 10308
rect 8024 10364 8088 10368
rect 8024 10308 8028 10364
rect 8028 10308 8084 10364
rect 8084 10308 8088 10364
rect 8024 10304 8088 10308
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 2700 9820 2764 9824
rect 2700 9764 2704 9820
rect 2704 9764 2760 9820
rect 2760 9764 2764 9820
rect 2700 9760 2764 9764
rect 2780 9820 2844 9824
rect 2780 9764 2784 9820
rect 2784 9764 2840 9820
rect 2840 9764 2844 9820
rect 2780 9760 2844 9764
rect 2860 9820 2924 9824
rect 2860 9764 2864 9820
rect 2864 9764 2920 9820
rect 2920 9764 2924 9820
rect 2860 9760 2924 9764
rect 2940 9820 3004 9824
rect 2940 9764 2944 9820
rect 2944 9764 3000 9820
rect 3000 9764 3004 9820
rect 2940 9760 3004 9764
rect 6196 9820 6260 9824
rect 6196 9764 6200 9820
rect 6200 9764 6256 9820
rect 6256 9764 6260 9820
rect 6196 9760 6260 9764
rect 6276 9820 6340 9824
rect 6276 9764 6280 9820
rect 6280 9764 6336 9820
rect 6336 9764 6340 9820
rect 6276 9760 6340 9764
rect 6356 9820 6420 9824
rect 6356 9764 6360 9820
rect 6360 9764 6416 9820
rect 6416 9764 6420 9820
rect 6356 9760 6420 9764
rect 6436 9820 6500 9824
rect 6436 9764 6440 9820
rect 6440 9764 6496 9820
rect 6496 9764 6500 9820
rect 6436 9760 6500 9764
rect 9692 9820 9756 9824
rect 9692 9764 9696 9820
rect 9696 9764 9752 9820
rect 9752 9764 9756 9820
rect 9692 9760 9756 9764
rect 9772 9820 9836 9824
rect 9772 9764 9776 9820
rect 9776 9764 9832 9820
rect 9832 9764 9836 9820
rect 9772 9760 9836 9764
rect 9852 9820 9916 9824
rect 9852 9764 9856 9820
rect 9856 9764 9912 9820
rect 9912 9764 9916 9820
rect 9852 9760 9916 9764
rect 9932 9820 9996 9824
rect 9932 9764 9936 9820
rect 9936 9764 9992 9820
rect 9992 9764 9996 9820
rect 9932 9760 9996 9764
rect 4448 9276 4512 9280
rect 4448 9220 4452 9276
rect 4452 9220 4508 9276
rect 4508 9220 4512 9276
rect 4448 9216 4512 9220
rect 4528 9276 4592 9280
rect 4528 9220 4532 9276
rect 4532 9220 4588 9276
rect 4588 9220 4592 9276
rect 4528 9216 4592 9220
rect 4608 9276 4672 9280
rect 4608 9220 4612 9276
rect 4612 9220 4668 9276
rect 4668 9220 4672 9276
rect 4608 9216 4672 9220
rect 4688 9276 4752 9280
rect 4688 9220 4692 9276
rect 4692 9220 4748 9276
rect 4748 9220 4752 9276
rect 4688 9216 4752 9220
rect 7944 9276 8008 9280
rect 7944 9220 7948 9276
rect 7948 9220 8004 9276
rect 8004 9220 8008 9276
rect 7944 9216 8008 9220
rect 8024 9276 8088 9280
rect 8024 9220 8028 9276
rect 8028 9220 8084 9276
rect 8084 9220 8088 9276
rect 8024 9216 8088 9220
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 2700 8732 2764 8736
rect 2700 8676 2704 8732
rect 2704 8676 2760 8732
rect 2760 8676 2764 8732
rect 2700 8672 2764 8676
rect 2780 8732 2844 8736
rect 2780 8676 2784 8732
rect 2784 8676 2840 8732
rect 2840 8676 2844 8732
rect 2780 8672 2844 8676
rect 2860 8732 2924 8736
rect 2860 8676 2864 8732
rect 2864 8676 2920 8732
rect 2920 8676 2924 8732
rect 2860 8672 2924 8676
rect 2940 8732 3004 8736
rect 2940 8676 2944 8732
rect 2944 8676 3000 8732
rect 3000 8676 3004 8732
rect 2940 8672 3004 8676
rect 6196 8732 6260 8736
rect 6196 8676 6200 8732
rect 6200 8676 6256 8732
rect 6256 8676 6260 8732
rect 6196 8672 6260 8676
rect 6276 8732 6340 8736
rect 6276 8676 6280 8732
rect 6280 8676 6336 8732
rect 6336 8676 6340 8732
rect 6276 8672 6340 8676
rect 6356 8732 6420 8736
rect 6356 8676 6360 8732
rect 6360 8676 6416 8732
rect 6416 8676 6420 8732
rect 6356 8672 6420 8676
rect 6436 8732 6500 8736
rect 6436 8676 6440 8732
rect 6440 8676 6496 8732
rect 6496 8676 6500 8732
rect 6436 8672 6500 8676
rect 9692 8732 9756 8736
rect 9692 8676 9696 8732
rect 9696 8676 9752 8732
rect 9752 8676 9756 8732
rect 9692 8672 9756 8676
rect 9772 8732 9836 8736
rect 9772 8676 9776 8732
rect 9776 8676 9832 8732
rect 9832 8676 9836 8732
rect 9772 8672 9836 8676
rect 9852 8732 9916 8736
rect 9852 8676 9856 8732
rect 9856 8676 9912 8732
rect 9912 8676 9916 8732
rect 9852 8672 9916 8676
rect 9932 8732 9996 8736
rect 9932 8676 9936 8732
rect 9936 8676 9992 8732
rect 9992 8676 9996 8732
rect 9932 8672 9996 8676
rect 4448 8188 4512 8192
rect 4448 8132 4452 8188
rect 4452 8132 4508 8188
rect 4508 8132 4512 8188
rect 4448 8128 4512 8132
rect 4528 8188 4592 8192
rect 4528 8132 4532 8188
rect 4532 8132 4588 8188
rect 4588 8132 4592 8188
rect 4528 8128 4592 8132
rect 4608 8188 4672 8192
rect 4608 8132 4612 8188
rect 4612 8132 4668 8188
rect 4668 8132 4672 8188
rect 4608 8128 4672 8132
rect 4688 8188 4752 8192
rect 4688 8132 4692 8188
rect 4692 8132 4748 8188
rect 4748 8132 4752 8188
rect 4688 8128 4752 8132
rect 7944 8188 8008 8192
rect 7944 8132 7948 8188
rect 7948 8132 8004 8188
rect 8004 8132 8008 8188
rect 7944 8128 8008 8132
rect 8024 8188 8088 8192
rect 8024 8132 8028 8188
rect 8028 8132 8084 8188
rect 8084 8132 8088 8188
rect 8024 8128 8088 8132
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 2700 7644 2764 7648
rect 2700 7588 2704 7644
rect 2704 7588 2760 7644
rect 2760 7588 2764 7644
rect 2700 7584 2764 7588
rect 2780 7644 2844 7648
rect 2780 7588 2784 7644
rect 2784 7588 2840 7644
rect 2840 7588 2844 7644
rect 2780 7584 2844 7588
rect 2860 7644 2924 7648
rect 2860 7588 2864 7644
rect 2864 7588 2920 7644
rect 2920 7588 2924 7644
rect 2860 7584 2924 7588
rect 2940 7644 3004 7648
rect 2940 7588 2944 7644
rect 2944 7588 3000 7644
rect 3000 7588 3004 7644
rect 2940 7584 3004 7588
rect 6196 7644 6260 7648
rect 6196 7588 6200 7644
rect 6200 7588 6256 7644
rect 6256 7588 6260 7644
rect 6196 7584 6260 7588
rect 6276 7644 6340 7648
rect 6276 7588 6280 7644
rect 6280 7588 6336 7644
rect 6336 7588 6340 7644
rect 6276 7584 6340 7588
rect 6356 7644 6420 7648
rect 6356 7588 6360 7644
rect 6360 7588 6416 7644
rect 6416 7588 6420 7644
rect 6356 7584 6420 7588
rect 6436 7644 6500 7648
rect 6436 7588 6440 7644
rect 6440 7588 6496 7644
rect 6496 7588 6500 7644
rect 6436 7584 6500 7588
rect 9692 7644 9756 7648
rect 9692 7588 9696 7644
rect 9696 7588 9752 7644
rect 9752 7588 9756 7644
rect 9692 7584 9756 7588
rect 9772 7644 9836 7648
rect 9772 7588 9776 7644
rect 9776 7588 9832 7644
rect 9832 7588 9836 7644
rect 9772 7584 9836 7588
rect 9852 7644 9916 7648
rect 9852 7588 9856 7644
rect 9856 7588 9912 7644
rect 9912 7588 9916 7644
rect 9852 7584 9916 7588
rect 9932 7644 9996 7648
rect 9932 7588 9936 7644
rect 9936 7588 9992 7644
rect 9992 7588 9996 7644
rect 9932 7584 9996 7588
rect 4448 7100 4512 7104
rect 4448 7044 4452 7100
rect 4452 7044 4508 7100
rect 4508 7044 4512 7100
rect 4448 7040 4512 7044
rect 4528 7100 4592 7104
rect 4528 7044 4532 7100
rect 4532 7044 4588 7100
rect 4588 7044 4592 7100
rect 4528 7040 4592 7044
rect 4608 7100 4672 7104
rect 4608 7044 4612 7100
rect 4612 7044 4668 7100
rect 4668 7044 4672 7100
rect 4608 7040 4672 7044
rect 4688 7100 4752 7104
rect 4688 7044 4692 7100
rect 4692 7044 4748 7100
rect 4748 7044 4752 7100
rect 4688 7040 4752 7044
rect 7944 7100 8008 7104
rect 7944 7044 7948 7100
rect 7948 7044 8004 7100
rect 8004 7044 8008 7100
rect 7944 7040 8008 7044
rect 8024 7100 8088 7104
rect 8024 7044 8028 7100
rect 8028 7044 8084 7100
rect 8084 7044 8088 7100
rect 8024 7040 8088 7044
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 2700 6556 2764 6560
rect 2700 6500 2704 6556
rect 2704 6500 2760 6556
rect 2760 6500 2764 6556
rect 2700 6496 2764 6500
rect 2780 6556 2844 6560
rect 2780 6500 2784 6556
rect 2784 6500 2840 6556
rect 2840 6500 2844 6556
rect 2780 6496 2844 6500
rect 2860 6556 2924 6560
rect 2860 6500 2864 6556
rect 2864 6500 2920 6556
rect 2920 6500 2924 6556
rect 2860 6496 2924 6500
rect 2940 6556 3004 6560
rect 2940 6500 2944 6556
rect 2944 6500 3000 6556
rect 3000 6500 3004 6556
rect 2940 6496 3004 6500
rect 6196 6556 6260 6560
rect 6196 6500 6200 6556
rect 6200 6500 6256 6556
rect 6256 6500 6260 6556
rect 6196 6496 6260 6500
rect 6276 6556 6340 6560
rect 6276 6500 6280 6556
rect 6280 6500 6336 6556
rect 6336 6500 6340 6556
rect 6276 6496 6340 6500
rect 6356 6556 6420 6560
rect 6356 6500 6360 6556
rect 6360 6500 6416 6556
rect 6416 6500 6420 6556
rect 6356 6496 6420 6500
rect 6436 6556 6500 6560
rect 6436 6500 6440 6556
rect 6440 6500 6496 6556
rect 6496 6500 6500 6556
rect 6436 6496 6500 6500
rect 9692 6556 9756 6560
rect 9692 6500 9696 6556
rect 9696 6500 9752 6556
rect 9752 6500 9756 6556
rect 9692 6496 9756 6500
rect 9772 6556 9836 6560
rect 9772 6500 9776 6556
rect 9776 6500 9832 6556
rect 9832 6500 9836 6556
rect 9772 6496 9836 6500
rect 9852 6556 9916 6560
rect 9852 6500 9856 6556
rect 9856 6500 9912 6556
rect 9912 6500 9916 6556
rect 9852 6496 9916 6500
rect 9932 6556 9996 6560
rect 9932 6500 9936 6556
rect 9936 6500 9992 6556
rect 9992 6500 9996 6556
rect 9932 6496 9996 6500
rect 4448 6012 4512 6016
rect 4448 5956 4452 6012
rect 4452 5956 4508 6012
rect 4508 5956 4512 6012
rect 4448 5952 4512 5956
rect 4528 6012 4592 6016
rect 4528 5956 4532 6012
rect 4532 5956 4588 6012
rect 4588 5956 4592 6012
rect 4528 5952 4592 5956
rect 4608 6012 4672 6016
rect 4608 5956 4612 6012
rect 4612 5956 4668 6012
rect 4668 5956 4672 6012
rect 4608 5952 4672 5956
rect 4688 6012 4752 6016
rect 4688 5956 4692 6012
rect 4692 5956 4748 6012
rect 4748 5956 4752 6012
rect 4688 5952 4752 5956
rect 7944 6012 8008 6016
rect 7944 5956 7948 6012
rect 7948 5956 8004 6012
rect 8004 5956 8008 6012
rect 7944 5952 8008 5956
rect 8024 6012 8088 6016
rect 8024 5956 8028 6012
rect 8028 5956 8084 6012
rect 8084 5956 8088 6012
rect 8024 5952 8088 5956
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 2700 5468 2764 5472
rect 2700 5412 2704 5468
rect 2704 5412 2760 5468
rect 2760 5412 2764 5468
rect 2700 5408 2764 5412
rect 2780 5468 2844 5472
rect 2780 5412 2784 5468
rect 2784 5412 2840 5468
rect 2840 5412 2844 5468
rect 2780 5408 2844 5412
rect 2860 5468 2924 5472
rect 2860 5412 2864 5468
rect 2864 5412 2920 5468
rect 2920 5412 2924 5468
rect 2860 5408 2924 5412
rect 2940 5468 3004 5472
rect 2940 5412 2944 5468
rect 2944 5412 3000 5468
rect 3000 5412 3004 5468
rect 2940 5408 3004 5412
rect 6196 5468 6260 5472
rect 6196 5412 6200 5468
rect 6200 5412 6256 5468
rect 6256 5412 6260 5468
rect 6196 5408 6260 5412
rect 6276 5468 6340 5472
rect 6276 5412 6280 5468
rect 6280 5412 6336 5468
rect 6336 5412 6340 5468
rect 6276 5408 6340 5412
rect 6356 5468 6420 5472
rect 6356 5412 6360 5468
rect 6360 5412 6416 5468
rect 6416 5412 6420 5468
rect 6356 5408 6420 5412
rect 6436 5468 6500 5472
rect 6436 5412 6440 5468
rect 6440 5412 6496 5468
rect 6496 5412 6500 5468
rect 6436 5408 6500 5412
rect 9692 5468 9756 5472
rect 9692 5412 9696 5468
rect 9696 5412 9752 5468
rect 9752 5412 9756 5468
rect 9692 5408 9756 5412
rect 9772 5468 9836 5472
rect 9772 5412 9776 5468
rect 9776 5412 9832 5468
rect 9832 5412 9836 5468
rect 9772 5408 9836 5412
rect 9852 5468 9916 5472
rect 9852 5412 9856 5468
rect 9856 5412 9912 5468
rect 9912 5412 9916 5468
rect 9852 5408 9916 5412
rect 9932 5468 9996 5472
rect 9932 5412 9936 5468
rect 9936 5412 9992 5468
rect 9992 5412 9996 5468
rect 9932 5408 9996 5412
rect 4448 4924 4512 4928
rect 4448 4868 4452 4924
rect 4452 4868 4508 4924
rect 4508 4868 4512 4924
rect 4448 4864 4512 4868
rect 4528 4924 4592 4928
rect 4528 4868 4532 4924
rect 4532 4868 4588 4924
rect 4588 4868 4592 4924
rect 4528 4864 4592 4868
rect 4608 4924 4672 4928
rect 4608 4868 4612 4924
rect 4612 4868 4668 4924
rect 4668 4868 4672 4924
rect 4608 4864 4672 4868
rect 4688 4924 4752 4928
rect 4688 4868 4692 4924
rect 4692 4868 4748 4924
rect 4748 4868 4752 4924
rect 4688 4864 4752 4868
rect 7944 4924 8008 4928
rect 7944 4868 7948 4924
rect 7948 4868 8004 4924
rect 8004 4868 8008 4924
rect 7944 4864 8008 4868
rect 8024 4924 8088 4928
rect 8024 4868 8028 4924
rect 8028 4868 8084 4924
rect 8084 4868 8088 4924
rect 8024 4864 8088 4868
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 2700 4380 2764 4384
rect 2700 4324 2704 4380
rect 2704 4324 2760 4380
rect 2760 4324 2764 4380
rect 2700 4320 2764 4324
rect 2780 4380 2844 4384
rect 2780 4324 2784 4380
rect 2784 4324 2840 4380
rect 2840 4324 2844 4380
rect 2780 4320 2844 4324
rect 2860 4380 2924 4384
rect 2860 4324 2864 4380
rect 2864 4324 2920 4380
rect 2920 4324 2924 4380
rect 2860 4320 2924 4324
rect 2940 4380 3004 4384
rect 2940 4324 2944 4380
rect 2944 4324 3000 4380
rect 3000 4324 3004 4380
rect 2940 4320 3004 4324
rect 6196 4380 6260 4384
rect 6196 4324 6200 4380
rect 6200 4324 6256 4380
rect 6256 4324 6260 4380
rect 6196 4320 6260 4324
rect 6276 4380 6340 4384
rect 6276 4324 6280 4380
rect 6280 4324 6336 4380
rect 6336 4324 6340 4380
rect 6276 4320 6340 4324
rect 6356 4380 6420 4384
rect 6356 4324 6360 4380
rect 6360 4324 6416 4380
rect 6416 4324 6420 4380
rect 6356 4320 6420 4324
rect 6436 4380 6500 4384
rect 6436 4324 6440 4380
rect 6440 4324 6496 4380
rect 6496 4324 6500 4380
rect 6436 4320 6500 4324
rect 9692 4380 9756 4384
rect 9692 4324 9696 4380
rect 9696 4324 9752 4380
rect 9752 4324 9756 4380
rect 9692 4320 9756 4324
rect 9772 4380 9836 4384
rect 9772 4324 9776 4380
rect 9776 4324 9832 4380
rect 9832 4324 9836 4380
rect 9772 4320 9836 4324
rect 9852 4380 9916 4384
rect 9852 4324 9856 4380
rect 9856 4324 9912 4380
rect 9912 4324 9916 4380
rect 9852 4320 9916 4324
rect 9932 4380 9996 4384
rect 9932 4324 9936 4380
rect 9936 4324 9992 4380
rect 9992 4324 9996 4380
rect 9932 4320 9996 4324
rect 4448 3836 4512 3840
rect 4448 3780 4452 3836
rect 4452 3780 4508 3836
rect 4508 3780 4512 3836
rect 4448 3776 4512 3780
rect 4528 3836 4592 3840
rect 4528 3780 4532 3836
rect 4532 3780 4588 3836
rect 4588 3780 4592 3836
rect 4528 3776 4592 3780
rect 4608 3836 4672 3840
rect 4608 3780 4612 3836
rect 4612 3780 4668 3836
rect 4668 3780 4672 3836
rect 4608 3776 4672 3780
rect 4688 3836 4752 3840
rect 4688 3780 4692 3836
rect 4692 3780 4748 3836
rect 4748 3780 4752 3836
rect 4688 3776 4752 3780
rect 7944 3836 8008 3840
rect 7944 3780 7948 3836
rect 7948 3780 8004 3836
rect 8004 3780 8008 3836
rect 7944 3776 8008 3780
rect 8024 3836 8088 3840
rect 8024 3780 8028 3836
rect 8028 3780 8084 3836
rect 8084 3780 8088 3836
rect 8024 3776 8088 3780
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 2700 3292 2764 3296
rect 2700 3236 2704 3292
rect 2704 3236 2760 3292
rect 2760 3236 2764 3292
rect 2700 3232 2764 3236
rect 2780 3292 2844 3296
rect 2780 3236 2784 3292
rect 2784 3236 2840 3292
rect 2840 3236 2844 3292
rect 2780 3232 2844 3236
rect 2860 3292 2924 3296
rect 2860 3236 2864 3292
rect 2864 3236 2920 3292
rect 2920 3236 2924 3292
rect 2860 3232 2924 3236
rect 2940 3292 3004 3296
rect 2940 3236 2944 3292
rect 2944 3236 3000 3292
rect 3000 3236 3004 3292
rect 2940 3232 3004 3236
rect 6196 3292 6260 3296
rect 6196 3236 6200 3292
rect 6200 3236 6256 3292
rect 6256 3236 6260 3292
rect 6196 3232 6260 3236
rect 6276 3292 6340 3296
rect 6276 3236 6280 3292
rect 6280 3236 6336 3292
rect 6336 3236 6340 3292
rect 6276 3232 6340 3236
rect 6356 3292 6420 3296
rect 6356 3236 6360 3292
rect 6360 3236 6416 3292
rect 6416 3236 6420 3292
rect 6356 3232 6420 3236
rect 6436 3292 6500 3296
rect 6436 3236 6440 3292
rect 6440 3236 6496 3292
rect 6496 3236 6500 3292
rect 6436 3232 6500 3236
rect 9692 3292 9756 3296
rect 9692 3236 9696 3292
rect 9696 3236 9752 3292
rect 9752 3236 9756 3292
rect 9692 3232 9756 3236
rect 9772 3292 9836 3296
rect 9772 3236 9776 3292
rect 9776 3236 9832 3292
rect 9832 3236 9836 3292
rect 9772 3232 9836 3236
rect 9852 3292 9916 3296
rect 9852 3236 9856 3292
rect 9856 3236 9912 3292
rect 9912 3236 9916 3292
rect 9852 3232 9916 3236
rect 9932 3292 9996 3296
rect 9932 3236 9936 3292
rect 9936 3236 9992 3292
rect 9992 3236 9996 3292
rect 9932 3232 9996 3236
rect 4448 2748 4512 2752
rect 4448 2692 4452 2748
rect 4452 2692 4508 2748
rect 4508 2692 4512 2748
rect 4448 2688 4512 2692
rect 4528 2748 4592 2752
rect 4528 2692 4532 2748
rect 4532 2692 4588 2748
rect 4588 2692 4592 2748
rect 4528 2688 4592 2692
rect 4608 2748 4672 2752
rect 4608 2692 4612 2748
rect 4612 2692 4668 2748
rect 4668 2692 4672 2748
rect 4608 2688 4672 2692
rect 4688 2748 4752 2752
rect 4688 2692 4692 2748
rect 4692 2692 4748 2748
rect 4748 2692 4752 2748
rect 4688 2688 4752 2692
rect 7944 2748 8008 2752
rect 7944 2692 7948 2748
rect 7948 2692 8004 2748
rect 8004 2692 8008 2748
rect 7944 2688 8008 2692
rect 8024 2748 8088 2752
rect 8024 2692 8028 2748
rect 8028 2692 8084 2748
rect 8084 2692 8088 2748
rect 8024 2688 8088 2692
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 2700 2204 2764 2208
rect 2700 2148 2704 2204
rect 2704 2148 2760 2204
rect 2760 2148 2764 2204
rect 2700 2144 2764 2148
rect 2780 2204 2844 2208
rect 2780 2148 2784 2204
rect 2784 2148 2840 2204
rect 2840 2148 2844 2204
rect 2780 2144 2844 2148
rect 2860 2204 2924 2208
rect 2860 2148 2864 2204
rect 2864 2148 2920 2204
rect 2920 2148 2924 2204
rect 2860 2144 2924 2148
rect 2940 2204 3004 2208
rect 2940 2148 2944 2204
rect 2944 2148 3000 2204
rect 3000 2148 3004 2204
rect 2940 2144 3004 2148
rect 6196 2204 6260 2208
rect 6196 2148 6200 2204
rect 6200 2148 6256 2204
rect 6256 2148 6260 2204
rect 6196 2144 6260 2148
rect 6276 2204 6340 2208
rect 6276 2148 6280 2204
rect 6280 2148 6336 2204
rect 6336 2148 6340 2204
rect 6276 2144 6340 2148
rect 6356 2204 6420 2208
rect 6356 2148 6360 2204
rect 6360 2148 6416 2204
rect 6416 2148 6420 2204
rect 6356 2144 6420 2148
rect 6436 2204 6500 2208
rect 6436 2148 6440 2204
rect 6440 2148 6496 2204
rect 6496 2148 6500 2204
rect 6436 2144 6500 2148
rect 9692 2204 9756 2208
rect 9692 2148 9696 2204
rect 9696 2148 9752 2204
rect 9752 2148 9756 2204
rect 9692 2144 9756 2148
rect 9772 2204 9836 2208
rect 9772 2148 9776 2204
rect 9776 2148 9832 2204
rect 9832 2148 9836 2204
rect 9772 2144 9836 2148
rect 9852 2204 9916 2208
rect 9852 2148 9856 2204
rect 9856 2148 9912 2204
rect 9912 2148 9916 2204
rect 9852 2144 9916 2148
rect 9932 2204 9996 2208
rect 9932 2148 9936 2204
rect 9936 2148 9992 2204
rect 9992 2148 9996 2204
rect 9932 2144 9996 2148
<< metal4 >>
rect 2692 12000 3012 12560
rect 2692 11936 2700 12000
rect 2764 11936 2780 12000
rect 2844 11936 2860 12000
rect 2924 11936 2940 12000
rect 3004 11936 3012 12000
rect 2692 10912 3012 11936
rect 2692 10848 2700 10912
rect 2764 10848 2780 10912
rect 2844 10848 2860 10912
rect 2924 10848 2940 10912
rect 3004 10848 3012 10912
rect 2692 9824 3012 10848
rect 2692 9760 2700 9824
rect 2764 9760 2780 9824
rect 2844 9760 2860 9824
rect 2924 9760 2940 9824
rect 3004 9760 3012 9824
rect 2692 8736 3012 9760
rect 2692 8672 2700 8736
rect 2764 8672 2780 8736
rect 2844 8672 2860 8736
rect 2924 8672 2940 8736
rect 3004 8672 3012 8736
rect 2692 7648 3012 8672
rect 2692 7584 2700 7648
rect 2764 7584 2780 7648
rect 2844 7584 2860 7648
rect 2924 7584 2940 7648
rect 3004 7584 3012 7648
rect 2692 6560 3012 7584
rect 2692 6496 2700 6560
rect 2764 6496 2780 6560
rect 2844 6496 2860 6560
rect 2924 6496 2940 6560
rect 3004 6496 3012 6560
rect 2692 5472 3012 6496
rect 2692 5408 2700 5472
rect 2764 5408 2780 5472
rect 2844 5408 2860 5472
rect 2924 5408 2940 5472
rect 3004 5408 3012 5472
rect 2692 4384 3012 5408
rect 2692 4320 2700 4384
rect 2764 4320 2780 4384
rect 2844 4320 2860 4384
rect 2924 4320 2940 4384
rect 3004 4320 3012 4384
rect 2692 3296 3012 4320
rect 2692 3232 2700 3296
rect 2764 3232 2780 3296
rect 2844 3232 2860 3296
rect 2924 3232 2940 3296
rect 3004 3232 3012 3296
rect 2692 2208 3012 3232
rect 2692 2144 2700 2208
rect 2764 2144 2780 2208
rect 2844 2144 2860 2208
rect 2924 2144 2940 2208
rect 3004 2144 3012 2208
rect 2692 2128 3012 2144
rect 4440 12544 4760 12560
rect 4440 12480 4448 12544
rect 4512 12480 4528 12544
rect 4592 12480 4608 12544
rect 4672 12480 4688 12544
rect 4752 12480 4760 12544
rect 4440 11456 4760 12480
rect 4440 11392 4448 11456
rect 4512 11392 4528 11456
rect 4592 11392 4608 11456
rect 4672 11392 4688 11456
rect 4752 11392 4760 11456
rect 4440 10368 4760 11392
rect 4440 10304 4448 10368
rect 4512 10304 4528 10368
rect 4592 10304 4608 10368
rect 4672 10304 4688 10368
rect 4752 10304 4760 10368
rect 4440 9280 4760 10304
rect 4440 9216 4448 9280
rect 4512 9216 4528 9280
rect 4592 9216 4608 9280
rect 4672 9216 4688 9280
rect 4752 9216 4760 9280
rect 4440 8192 4760 9216
rect 4440 8128 4448 8192
rect 4512 8128 4528 8192
rect 4592 8128 4608 8192
rect 4672 8128 4688 8192
rect 4752 8128 4760 8192
rect 4440 7104 4760 8128
rect 4440 7040 4448 7104
rect 4512 7040 4528 7104
rect 4592 7040 4608 7104
rect 4672 7040 4688 7104
rect 4752 7040 4760 7104
rect 4440 6016 4760 7040
rect 4440 5952 4448 6016
rect 4512 5952 4528 6016
rect 4592 5952 4608 6016
rect 4672 5952 4688 6016
rect 4752 5952 4760 6016
rect 4440 4928 4760 5952
rect 4440 4864 4448 4928
rect 4512 4864 4528 4928
rect 4592 4864 4608 4928
rect 4672 4864 4688 4928
rect 4752 4864 4760 4928
rect 4440 3840 4760 4864
rect 4440 3776 4448 3840
rect 4512 3776 4528 3840
rect 4592 3776 4608 3840
rect 4672 3776 4688 3840
rect 4752 3776 4760 3840
rect 4440 2752 4760 3776
rect 4440 2688 4448 2752
rect 4512 2688 4528 2752
rect 4592 2688 4608 2752
rect 4672 2688 4688 2752
rect 4752 2688 4760 2752
rect 4440 2128 4760 2688
rect 6188 12000 6508 12560
rect 6188 11936 6196 12000
rect 6260 11936 6276 12000
rect 6340 11936 6356 12000
rect 6420 11936 6436 12000
rect 6500 11936 6508 12000
rect 6188 10912 6508 11936
rect 6188 10848 6196 10912
rect 6260 10848 6276 10912
rect 6340 10848 6356 10912
rect 6420 10848 6436 10912
rect 6500 10848 6508 10912
rect 6188 9824 6508 10848
rect 6188 9760 6196 9824
rect 6260 9760 6276 9824
rect 6340 9760 6356 9824
rect 6420 9760 6436 9824
rect 6500 9760 6508 9824
rect 6188 8736 6508 9760
rect 6188 8672 6196 8736
rect 6260 8672 6276 8736
rect 6340 8672 6356 8736
rect 6420 8672 6436 8736
rect 6500 8672 6508 8736
rect 6188 7648 6508 8672
rect 6188 7584 6196 7648
rect 6260 7584 6276 7648
rect 6340 7584 6356 7648
rect 6420 7584 6436 7648
rect 6500 7584 6508 7648
rect 6188 6560 6508 7584
rect 6188 6496 6196 6560
rect 6260 6496 6276 6560
rect 6340 6496 6356 6560
rect 6420 6496 6436 6560
rect 6500 6496 6508 6560
rect 6188 5472 6508 6496
rect 6188 5408 6196 5472
rect 6260 5408 6276 5472
rect 6340 5408 6356 5472
rect 6420 5408 6436 5472
rect 6500 5408 6508 5472
rect 6188 4384 6508 5408
rect 6188 4320 6196 4384
rect 6260 4320 6276 4384
rect 6340 4320 6356 4384
rect 6420 4320 6436 4384
rect 6500 4320 6508 4384
rect 6188 3296 6508 4320
rect 6188 3232 6196 3296
rect 6260 3232 6276 3296
rect 6340 3232 6356 3296
rect 6420 3232 6436 3296
rect 6500 3232 6508 3296
rect 6188 2208 6508 3232
rect 6188 2144 6196 2208
rect 6260 2144 6276 2208
rect 6340 2144 6356 2208
rect 6420 2144 6436 2208
rect 6500 2144 6508 2208
rect 6188 2128 6508 2144
rect 7936 12544 8256 12560
rect 7936 12480 7944 12544
rect 8008 12480 8024 12544
rect 8088 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8256 12544
rect 7936 11456 8256 12480
rect 7936 11392 7944 11456
rect 8008 11392 8024 11456
rect 8088 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8256 11456
rect 7936 10368 8256 11392
rect 7936 10304 7944 10368
rect 8008 10304 8024 10368
rect 8088 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8256 10368
rect 7936 9280 8256 10304
rect 7936 9216 7944 9280
rect 8008 9216 8024 9280
rect 8088 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8256 9280
rect 7936 8192 8256 9216
rect 7936 8128 7944 8192
rect 8008 8128 8024 8192
rect 8088 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8256 8192
rect 7936 7104 8256 8128
rect 7936 7040 7944 7104
rect 8008 7040 8024 7104
rect 8088 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8256 7104
rect 7936 6016 8256 7040
rect 7936 5952 7944 6016
rect 8008 5952 8024 6016
rect 8088 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8256 6016
rect 7936 4928 8256 5952
rect 7936 4864 7944 4928
rect 8008 4864 8024 4928
rect 8088 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8256 4928
rect 7936 3840 8256 4864
rect 7936 3776 7944 3840
rect 8008 3776 8024 3840
rect 8088 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8256 3840
rect 7936 2752 8256 3776
rect 7936 2688 7944 2752
rect 8008 2688 8024 2752
rect 8088 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8256 2752
rect 7936 2128 8256 2688
rect 9684 12000 10004 12560
rect 9684 11936 9692 12000
rect 9756 11936 9772 12000
rect 9836 11936 9852 12000
rect 9916 11936 9932 12000
rect 9996 11936 10004 12000
rect 9684 10912 10004 11936
rect 9684 10848 9692 10912
rect 9756 10848 9772 10912
rect 9836 10848 9852 10912
rect 9916 10848 9932 10912
rect 9996 10848 10004 10912
rect 9684 9824 10004 10848
rect 9684 9760 9692 9824
rect 9756 9760 9772 9824
rect 9836 9760 9852 9824
rect 9916 9760 9932 9824
rect 9996 9760 10004 9824
rect 9684 8736 10004 9760
rect 9684 8672 9692 8736
rect 9756 8672 9772 8736
rect 9836 8672 9852 8736
rect 9916 8672 9932 8736
rect 9996 8672 10004 8736
rect 9684 7648 10004 8672
rect 9684 7584 9692 7648
rect 9756 7584 9772 7648
rect 9836 7584 9852 7648
rect 9916 7584 9932 7648
rect 9996 7584 10004 7648
rect 9684 6560 10004 7584
rect 9684 6496 9692 6560
rect 9756 6496 9772 6560
rect 9836 6496 9852 6560
rect 9916 6496 9932 6560
rect 9996 6496 10004 6560
rect 9684 5472 10004 6496
rect 9684 5408 9692 5472
rect 9756 5408 9772 5472
rect 9836 5408 9852 5472
rect 9916 5408 9932 5472
rect 9996 5408 10004 5472
rect 9684 4384 10004 5408
rect 9684 4320 9692 4384
rect 9756 4320 9772 4384
rect 9836 4320 9852 4384
rect 9916 4320 9932 4384
rect 9996 4320 10004 4384
rect 9684 3296 10004 4320
rect 9684 3232 9692 3296
rect 9756 3232 9772 3296
rect 9836 3232 9852 3296
rect 9916 3232 9932 3296
rect 9996 3232 10004 3296
rect 9684 2208 10004 3232
rect 9684 2144 9692 2208
rect 9756 2144 9772 2208
rect 9836 2144 9852 2208
rect 9916 2144 9932 2208
rect 9996 2144 10004 2208
rect 9684 2128 10004 2144
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606969352
transform -1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_103
timestamp 1606969352
transform 1 0 10580 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _171_
timestamp 1606969352
transform 1 0 8464 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _183_
timestamp 1606969352
transform 1 0 10212 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606969352
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1606969352
transform 1 0 8924 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1606969352
transform 1 0 9752 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_98
timestamp 1606969352
transform 1 0 10120 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _102_
timestamp 1606969352
transform 1 0 6900 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606969352
transform 1 0 6808 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_72
timestamp 1606969352
transform 1 0 7728 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _157_
timestamp 1606969352
transform 1 0 5520 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_40
timestamp 1606969352
transform 1 0 4784 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_54
timestamp 1606969352
transform 1 0 6072 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _164_
timestamp 1606969352
transform 1 0 4324 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606969352
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606969352
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1606969352
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606969352
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606969352
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606969352
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606969352
transform -1 0 11592 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_106
timestamp 1606969352
transform 1 0 10856 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_110
timestamp 1606969352
transform 1 0 11224 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _179_
timestamp 1606969352
transform 1 0 9292 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 1606969352
transform 1 0 8556 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1606969352
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _103_
timestamp 1606969352
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _159_
timestamp 1606969352
transform 1 0 8096 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606969352
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_68
timestamp 1606969352
transform 1 0 7360 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _154_
timestamp 1606969352
transform 1 0 5520 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_17_40
timestamp 1606969352
transform 1 0 4784 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1606969352
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _162_
timestamp 1606969352
transform 1 0 4324 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _169_
timestamp 1606969352
transform 1 0 3128 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1606969352
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_27
timestamp 1606969352
transform 1 0 3588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606969352
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606969352
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1606969352
transform 1 0 2484 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606969352
transform -1 0 11592 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1606969352
transform 1 0 11224 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _161_
timestamp 1606969352
transform 1 0 9660 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606969352
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1606969352
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606969352
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_98
timestamp 1606969352
transform 1 0 10120 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_2  _158_
timestamp 1606969352
transform 1 0 7268 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_63
timestamp 1606969352
transform 1 0 6900 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_75
timestamp 1606969352
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_51
timestamp 1606969352
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _186_
timestamp 1606969352
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606969352
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1606969352
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _168_
timestamp 1606969352
transform 1 0 2760 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606969352
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606969352
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1606969352
transform 1 0 2484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606969352
transform -1 0 11592 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1606969352
transform 1 0 10764 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _156_
timestamp 1606969352
transform 1 0 9200 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_15_80
timestamp 1606969352
transform 1 0 8464 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1606969352
transform 1 0 9660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _086_
timestamp 1606969352
transform 1 0 6808 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _116_
timestamp 1606969352
transform 1 0 8004 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606969352
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_67
timestamp 1606969352
transform 1 0 7268 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _119_
timestamp 1606969352
transform 1 0 5520 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_15_40
timestamp 1606969352
transform 1 0 4784 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1606969352
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _137_
timestamp 1606969352
transform 1 0 4324 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _160_
timestamp 1606969352
transform 1 0 3128 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1606969352
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_27
timestamp 1606969352
transform 1 0 3588 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _165_
timestamp 1606969352
transform 1 0 1840 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606969352
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1606969352
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1606969352
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_13
timestamp 1606969352
transform 1 0 2300 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606969352
transform -1 0 11592 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606969352
transform -1 0 11592 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_110
timestamp 1606969352
transform 1 0 11224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_110
timestamp 1606969352
transform 1 0 11224 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _092_
timestamp 1606969352
transform 1 0 9660 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1606969352
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _146_
timestamp 1606969352
transform 1 0 9660 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606969352
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_85
timestamp 1606969352
transform 1 0 8924 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1606969352
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1606969352
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_98
timestamp 1606969352
transform 1 0 10120 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _089_
timestamp 1606969352
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _117_
timestamp 1606969352
transform 1 0 7268 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _144_
timestamp 1606969352
transform 1 0 8372 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606969352
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_71
timestamp 1606969352
transform 1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_73
timestamp 1606969352
transform 1 0 7820 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _091_
timestamp 1606969352
transform 1 0 5980 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _105_
timestamp 1606969352
transform 1 0 5428 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _120_
timestamp 1606969352
transform 1 0 4784 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1606969352
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_45
timestamp 1606969352
transform 1 0 5244 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_59
timestamp 1606969352
transform 1 0 6532 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _081_
timestamp 1606969352
transform 1 0 4232 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606969352
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_31
timestamp 1606969352
transform 1 0 3956 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1606969352
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1606969352
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1606969352
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_19
timestamp 1606969352
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _139_
timestamp 1606969352
transform 1 0 2300 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _155_
timestamp 1606969352
transform 1 0 2760 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1606969352
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_10
timestamp 1606969352
transform 1 0 2024 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _163_
timestamp 1606969352
transform 1 0 1564 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606969352
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606969352
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1606969352
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606969352
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606969352
transform -1 0 11592 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1606969352
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _088_
timestamp 1606969352
transform 1 0 9660 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606969352
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1606969352
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1606969352
transform 1 0 10120 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _153_
timestamp 1606969352
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_62
timestamp 1606969352
transform 1 0 6808 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_79
timestamp 1606969352
transform 1 0 8372 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _142_
timestamp 1606969352
transform 1 0 5704 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_42
timestamp 1606969352
transform 1 0 4968 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _141_
timestamp 1606969352
transform 1 0 4416 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606969352
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1606969352
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606969352
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _136_
timestamp 1606969352
transform 1 0 2760 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _140_
timestamp 1606969352
transform 1 0 1564 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606969352
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606969352
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_10
timestamp 1606969352
transform 1 0 2024 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606969352
transform -1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1606969352
transform 1 0 10580 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _143_
timestamp 1606969352
transform 1 0 10028 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _177_
timestamp 1606969352
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_89
timestamp 1606969352
transform 1 0 9292 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _172_
timestamp 1606969352
transform 1 0 6808 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606969352
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_72
timestamp 1606969352
transform 1 0 7728 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1606969352
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _173_
timestamp 1606969352
transform 1 0 4692 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_2  _181_
timestamp 1606969352
transform 1 0 3404 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_24
timestamp 1606969352
transform 1 0 3312 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_31
timestamp 1606969352
transform 1 0 3956 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _138_
timestamp 1606969352
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606969352
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_12
timestamp 1606969352
transform 1 0 2208 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606969352
transform -1 0 11592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_100
timestamp 1606969352
transform 1 0 10304 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_108
timestamp 1606969352
transform 1 0 11040 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _125_
timestamp 1606969352
transform 1 0 9660 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606969352
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1606969352
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _080_
timestamp 1606969352
transform 1 0 8096 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_68
timestamp 1606969352
transform 1 0 7360 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _129_
timestamp 1606969352
transform 1 0 5796 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_10_43
timestamp 1606969352
transform 1 0 5060 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _180_
timestamp 1606969352
transform 1 0 4140 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606969352
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1606969352
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1606969352
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _079_
timestamp 1606969352
transform 1 0 2760 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _118_
timestamp 1606969352
transform 1 0 1564 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606969352
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606969352
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_10
timestamp 1606969352
transform 1 0 2024 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606969352
transform -1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1606969352
transform 1 0 10764 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _132_
timestamp 1606969352
transform 1 0 8832 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1606969352
transform 1 0 9660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _149_
timestamp 1606969352
transform 1 0 6808 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606969352
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606969352
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_76
timestamp 1606969352
transform 1 0 8096 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_52
timestamp 1606969352
transform 1 0 5888 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _187_
timestamp 1606969352
transform 1 0 4140 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_24
timestamp 1606969352
transform 1 0 3312 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_32
timestamp 1606969352
transform 1 0 4048 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _167_
timestamp 1606969352
transform 1 0 2484 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606969352
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606969352
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606969352
transform -1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_103
timestamp 1606969352
transform 1 0 10580 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _127_
timestamp 1606969352
transform 1 0 9752 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606969352
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_83
timestamp 1606969352
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606969352
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1606969352
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _121_
timestamp 1606969352
transform 1 0 7912 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_66
timestamp 1606969352
transform 1 0 7176 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _099_
timestamp 1606969352
transform 1 0 5612 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1606969352
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _082_
timestamp 1606969352
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606969352
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1606969352
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _135_
timestamp 1606969352
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606969352
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1606969352
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_11
timestamp 1606969352
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606969352
transform -1 0 11592 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606969352
transform -1 0 11592 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_102
timestamp 1606969352
transform 1 0 10488 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_110
timestamp 1606969352
transform 1 0 11224 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1606969352
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _128_
timestamp 1606969352
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _130_
timestamp 1606969352
transform 1 0 8740 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606969352
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1606969352
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_97
timestamp 1606969352
transform 1 0 10028 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _083_
timestamp 1606969352
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _101_
timestamp 1606969352
transform 1 0 8096 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606969352
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_68
timestamp 1606969352
transform 1 0 7360 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_71
timestamp 1606969352
transform 1 0 7636 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _090_
timestamp 1606969352
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _106_
timestamp 1606969352
transform 1 0 4876 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1606969352
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1606969352
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _131_
timestamp 1606969352
transform 1 0 3312 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _188_
timestamp 1606969352
transform 1 0 4048 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606969352
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1606969352
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_33
timestamp 1606969352
transform 1 0 4140 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _104_
timestamp 1606969352
transform 1 0 2760 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _124_
timestamp 1606969352
transform 1 0 2024 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_10
timestamp 1606969352
transform 1 0 2024 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1606969352
transform 1 0 1932 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_16
timestamp 1606969352
transform 1 0 2576 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _134_
timestamp 1606969352
transform 1 0 1564 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606969352
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606969352
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606969352
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1606969352
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606969352
transform -1 0 11592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1606969352
transform 1 0 10580 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _126_
timestamp 1606969352
transform 1 0 9936 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_86
timestamp 1606969352
transform 1 0 9016 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1606969352
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _084_
timestamp 1606969352
transform 1 0 8372 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _098_
timestamp 1606969352
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606969352
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1606969352
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_71
timestamp 1606969352
transform 1 0 7636 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _085_
timestamp 1606969352
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_52
timestamp 1606969352
transform 1 0 5888 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _096_
timestamp 1606969352
transform 1 0 3680 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_20
timestamp 1606969352
transform 1 0 2944 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_35
timestamp 1606969352
transform 1 0 4324 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _133_
timestamp 1606969352
transform 1 0 2484 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606969352
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606969352
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606969352
transform -1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1606969352
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _115_
timestamp 1606969352
transform 1 0 9660 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1606969352
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1606969352
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1606969352
transform 1 0 10120 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_2  _175_
timestamp 1606969352
transform 1 0 7360 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_60
timestamp 1606969352
transform 1 0 6624 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_76
timestamp 1606969352
transform 1 0 8096 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _097_
timestamp 1606969352
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_43
timestamp 1606969352
transform 1 0 5060 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _087_
timestamp 1606969352
transform 1 0 4600 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1606969352
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1606969352
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 1606969352
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _151_
timestamp 1606969352
transform 1 0 2760 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _174_
timestamp 1606969352
transform 1 0 1564 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606969352
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1606969352
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_10
timestamp 1606969352
transform 1 0 2024 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606969352
transform -1 0 11592 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_110
timestamp 1606969352
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _147_
timestamp 1606969352
transform 1 0 9660 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_3_84
timestamp 1606969352
transform 1 0 8832 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_92
timestamp 1606969352
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606969352
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _114_
timestamp 1606969352
transform 1 0 8372 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _178_
timestamp 1606969352
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1606969352
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_71
timestamp 1606969352
transform 1 0 7636 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _108_
timestamp 1606969352
transform 1 0 5428 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1606969352
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _123_
timestamp 1606969352
transform 1 0 4232 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _170_
timestamp 1606969352
transform 1 0 3036 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_3_26
timestamp 1606969352
transform 1 0 3496 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 1606969352
transform 1 0 4692 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _184_
timestamp 1606969352
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606969352
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_7
timestamp 1606969352
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1606969352
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606969352
transform -1 0 11592 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_110
timestamp 1606969352
transform 1 0 11224 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _112_
timestamp 1606969352
transform 1 0 9660 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1606969352
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_82
timestamp 1606969352
transform 1 0 8648 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606969352
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1606969352
transform 1 0 10120 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _110_
timestamp 1606969352
transform 1 0 8188 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1606969352
transform 1 0 6808 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp 1606969352
transform 1 0 7912 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _107_
timestamp 1606969352
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _122_
timestamp 1606969352
transform 1 0 5060 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_2_48
timestamp 1606969352
transform 1 0 5520 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp 1606969352
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1606969352
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1606969352
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_35
timestamp 1606969352
transform 1 0 4324 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _182_
timestamp 1606969352
transform 1 0 2300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606969352
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1606969352
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1606969352
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_17
timestamp 1606969352
transform 1 0 2668 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606969352
transform -1 0 11592 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606969352
transform -1 0 11592 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1606969352
transform 1 0 10580 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _093_
timestamp 1606969352
transform 1 0 9752 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _111_
timestamp 1606969352
transform 1 0 10120 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1606969352
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1606969352
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_99
timestamp 1606969352
transform 1 0 10212 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_90
timestamp 1606969352
transform 1 0 9384 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _095_
timestamp 1606969352
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _100_
timestamp 1606969352
transform 1 0 8096 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_2  _113_
timestamp 1606969352
transform 1 0 6808 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _150_
timestamp 1606969352
transform 1 0 6900 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1606969352
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1606969352
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68
timestamp 1606969352
transform 1 0 7360 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_67
timestamp 1606969352
transform 1 0 7268 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1606969352
transform 1 0 8004 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _148_
timestamp 1606969352
transform 1 0 5520 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _152_
timestamp 1606969352
transform 1 0 5612 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp 1606969352
transform 1 0 4876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1606969352
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_40
timestamp 1606969352
transform 1 0 4784 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1606969352
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606969352
transform 1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _166_
timestamp 1606969352
transform 1 0 4324 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _176_
timestamp 1606969352
transform 1 0 4416 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1606969352
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23
timestamp 1606969352
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1606969352
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1606969352
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _185_
timestamp 1606969352
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606969352
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606969352
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1606969352
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1606969352
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606969352
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1606969352
transform 1 0 2484 0 1 2720
box -38 -48 774 592
<< labels >>
rlabel metal2 s 3422 14113 3478 14913 4 cbitin
port 1 nsew
rlabel metal2 s 3422 0 3478 800 4 cbitout
port 2 nsew
rlabel metal2 s 2042 14113 2098 14913 4 confclk
port 3 nsew
rlabel metal2 s 2042 0 2098 800 4 confclko
port 4 nsew
rlabel metal2 s 9126 0 9182 800 4 dempty
port 5 nsew
rlabel metal2 s 11978 0 12034 800 4 din[0]
port 6 nsew
rlabel metal2 s 10598 0 10654 800 4 din[1]
port 7 nsew
rlabel metal2 s 6274 0 6330 800 4 dout[0]
port 8 nsew
rlabel metal2 s 4894 0 4950 800 4 dout[1]
port 9 nsew
rlabel metal3 s 0 6128 800 6248 4 hempty
port 10 nsew
rlabel metal3 s 11969 8712 12769 8832 4 hempty2
port 11 nsew
rlabel metal3 s 0 8712 800 8832 4 lempty
port 12 nsew
rlabel metal3 s 0 13608 800 13728 4 lin[0]
port 13 nsew
rlabel metal3 s 0 11160 800 11280 4 lin[1]
port 14 nsew
rlabel metal3 s 0 3680 800 3800 4 lout[0]
port 15 nsew
rlabel metal3 s 0 1232 800 1352 4 lout[1]
port 16 nsew
rlabel metal3 s 11969 6128 12769 6248 4 rempty
port 17 nsew
rlabel metal2 s 662 14113 718 14913 4 reset
port 18 nsew
rlabel metal2 s 662 0 718 800 4 reseto
port 19 nsew
rlabel metal3 s 11969 3680 12769 3800 4 rin[0]
port 20 nsew
rlabel metal3 s 11969 1232 12769 1352 4 rin[1]
port 21 nsew
rlabel metal3 s 11969 13608 12769 13728 4 rout[0]
port 22 nsew
rlabel metal3 s 11969 11160 12769 11280 4 rout[1]
port 23 nsew
rlabel metal2 s 7746 14113 7802 14913 4 uempty
port 24 nsew
rlabel metal2 s 6274 14113 6330 14913 4 uin[0]
port 25 nsew
rlabel metal2 s 4894 14113 4950 14913 4 uin[1]
port 26 nsew
rlabel metal2 s 11978 14113 12034 14913 4 uout[0]
port 27 nsew
rlabel metal2 s 10598 14113 10654 14913 4 uout[1]
port 28 nsew
rlabel metal2 s 9126 14113 9182 14913 4 vempty
port 29 nsew
rlabel metal2 s 7746 0 7802 800 4 vempty2
port 30 nsew
rlabel metal4 s 2692 2128 3012 12560 4 VPWR
port 31 nsew
rlabel metal4 s 4440 2128 4760 12560 4 VGND
port 32 nsew
<< properties >>
string FIXED_BBOX 0 0 12769 14913
string GDS_FILE /project/openlane/morphle_ycell/runs/morphle_ycell/results/magic/ycell.gds
string GDS_END 496734
string GDS_START 176590
<< end >>
