// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module user_proj_example(wb_clk_i, wb_rst_i, wbs_ack_o, wbs_cyc_i, wbs_stb_i, wbs_we_i, vccd1, vssd1, vccd2, vssd2, vdda1, vssa1, vdda2, vssa2, io_in, io_oeb, io_out, la_data_in, la_data_out, la_oen, wbs_adr_i, wbs_dat_i, wbs_dat_o, wbs_sel_i);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire \clknet_0_counter.clk ;
  wire \clknet_1_0_0_counter.clk ;
  wire \clknet_1_1_0_counter.clk ;
  wire \clknet_2_0_0_counter.clk ;
  wire \clknet_2_1_0_counter.clk ;
  wire \clknet_2_2_0_counter.clk ;
  wire \clknet_2_3_0_counter.clk ;
  wire \clknet_3_0_0_counter.clk ;
  wire \clknet_3_1_0_counter.clk ;
  wire \clknet_3_2_0_counter.clk ;
  wire \clknet_3_3_0_counter.clk ;
  wire \clknet_3_4_0_counter.clk ;
  wire \clknet_3_5_0_counter.clk ;
  wire \clknet_3_6_0_counter.clk ;
  wire \clknet_3_7_0_counter.clk ;
  wire \counter.clk ;
  input [37:0] io_in;
  output [37:0] io_oeb;
  output [37:0] io_out;
  input [127:0] la_data_in;
  output [127:0] la_data_out;
  input [127:0] la_oen;
  input vccd1;
  input vccd2;
  input vdda1;
  input vdda2;
  input vssa1;
  input vssa2;
  input vssd1;
  input vssd2;
  input wb_clk_i;
  input wb_rst_i;
  output wbs_ack_o;
  input [31:0] wbs_adr_i;
  input wbs_cyc_i;
  input [31:0] wbs_dat_i;
  output [31:0] wbs_dat_o;
  input [3:0] wbs_sel_i;
  input wbs_stb_i;
  input wbs_we_i;
  sky130_fd_sc_hd__diode_2 ANTENNA_0 (
    .DIODE(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_1 (
    .DIODE(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_2 (
    .DIODE(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_3 (
    .DIODE(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_101 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1021 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1024 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1036 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1048 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1055 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1067 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1079 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1098 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1148 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_116 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1179 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1210 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1222 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1234 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1241 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_125 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1253 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1259 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_1263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1272 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_156 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_167 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_204 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_209 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_218 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_223 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_240 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_268 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_294 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_311 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_331 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_339 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_350 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_363 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_371 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_382 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_394 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_413 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_425 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_433 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_442 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_457 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_470 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_482 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_494 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_518 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_526 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_549 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_557 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_580 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_588 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_599 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_619 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_63 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_630 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_641 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_649 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_652 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_674 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_692 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_711 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_723 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_734 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_742 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_748 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_759 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_771 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_807 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_819 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_831 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_838 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_85 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_850 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_862 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_869 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_881 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_893 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_900 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_912 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_924 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_931 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_943 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_955 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_962 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_974 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_986 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_993 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_997 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_100_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_100_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_101_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_101_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_101_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_102_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_102_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_103_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_103_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_103_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_104_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_104_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_105_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_105_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_105_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_106_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_106_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_107_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_107_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_107_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_108_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_108_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_109_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_109_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_109_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_145 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_189 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_237 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_272 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_284 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_301 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_360 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_387 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_404 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_424 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_457 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_478 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_505 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_516 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_529 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_541 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_545 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_555 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_572 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_584 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_592 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_612 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_620 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_630 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_638 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_645 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_110_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_110_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_111_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_111_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_111_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_112_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_112_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_113_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_113_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_113_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_114_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_114_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_115_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_115_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_115_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_116_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_116_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_117_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_117_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_117_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_118_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_118_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_119_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_119_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_119_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_152 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_163 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_175 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_211 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_241 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_325 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_352 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_360 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_375 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_401 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_419 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_447 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_458 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_480 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_503 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_539 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_547 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_560 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_571 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_579 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_589 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_600 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_614 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_625 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_636 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_651 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_663 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_697 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_709 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_721 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_729 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_120_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_120_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_121_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_121_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_121_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_122_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_122_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_123_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_123_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_123_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_124_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_124_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_125_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_125_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_125_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_126_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_126_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_127_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_127_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_127_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_128_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_128_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_129_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_129_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_129_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_162 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_177 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_189 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_231 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_280 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_307 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_356 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_383 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_387 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_435 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_450 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_465 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_485 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_506 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_518 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_529 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_541 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_551 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_563 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_575 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_579 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_584 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_595 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_606 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_130_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_130_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_131_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_131_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_131_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_132_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_132_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_133_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_133_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_133_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_134_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_134_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_135_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_135_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_135_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_136_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_136_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_137_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_137_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_137_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_138_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_138_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_139_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_139_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_139_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_175 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_189 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_204 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_216 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_253 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_327 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_352 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_363 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_386 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_413 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_421 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_437 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_445 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_466 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_478 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_486 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_493 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_519 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_534 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_546 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_554 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_565 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_576 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_587 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_602 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_621 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_633 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_645 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_657 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_669 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_140_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_140_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_141_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_141_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_141_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_142_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_142_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_143_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_143_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_143_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_144_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_144_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_145_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_145_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_145_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_146_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_146_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_147_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_147_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_147_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_148_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_148_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_149_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_149_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_149_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_174 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_180 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_188 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_194 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_234 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_260 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_272 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_283 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_310 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_356 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_383 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_394 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_406 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_423 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_450 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_472 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_506 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_518 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_524 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_536 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_548 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_559 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_570 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_578 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_609 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_613 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_625 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_637 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_150_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_150_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_151_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_151_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_151_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_152_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_152_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_153_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_153_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_153_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_154_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_154_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_155_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_155_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_155_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_156_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_156_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_157_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_157_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_157_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_158_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_158_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_159_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_159_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_159_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_188 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_192 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_235 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_283 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_325 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_347 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_377 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_404 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_419 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_463 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_478 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_486 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_493 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_517 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_529 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_540 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_548 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_572 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_584 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_596 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_160_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_160_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_161_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_161_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_161_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_162_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_162_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_163_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_163_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_163_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_164_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_164_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_165_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_165_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_165_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_166_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_166_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_167_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_167_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_167_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_168_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_168_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_169_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_169_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_169_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_219 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_231 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_246 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_266 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_274 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_284 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_295 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_307 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_311 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_325 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_341 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_365 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_387 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_420 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_442 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_454 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_466 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_474 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_491 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_506 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_518 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_523 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_534 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_546 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_558 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_570 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_578 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_170_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_170_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_171_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_171_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_171_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_172_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_172_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_173_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_173_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_174_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_174_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_175_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_175_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_176_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_176_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_177_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_177_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_177_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_178_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_178_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_179_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_179_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_179_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_213 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_224 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_256 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_291 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_303 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_319 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_334 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_352 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_364 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_376 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_388 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_399 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_416 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_438 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_453 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_480 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_508 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_519 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_531 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_543 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_180_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_180_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_181_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_181_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_181_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_182_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_182_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_183_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_183_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_183_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_184_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_184_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_185_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_185_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_185_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_186_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_186_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_187_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_187_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_187_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_188_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_188_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_189_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_189_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_189_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_231 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_255 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_285 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_303 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_320 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_332 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_346 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_366 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_374 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_389 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_417 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_432 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_444 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_456 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_465 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_503 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_515 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_190_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_190_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_191_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_191_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_191_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_192_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_192_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_193_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_193_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_193_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_194_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_194_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_195_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_195_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_195_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_196_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_196_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_197_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_197_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_197_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_198_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_198_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_199_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_199_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_199_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_248 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_260 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_287 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_314 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_323 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_331 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_340 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_348 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_377 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_392 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_407 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_419 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_432 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_443 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_455 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_463 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_475 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_487 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_492 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_504 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_516 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_528 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_540 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_548 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1002 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1024 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1036 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1041 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1052 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1063 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1085 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1097 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1102 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1124 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1146 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1158 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1163 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1174 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1185 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1207 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1219 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1224 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1235 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1246 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1268 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_131 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_158 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_175 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_204 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_216 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_235 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_292 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_304 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_355 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_363 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_376 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_393 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_405 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_418 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_426 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_444 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_461 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_473 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_485 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_493 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_510 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_522 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_541 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_559 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_576 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_609 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_620 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_637 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_670 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_681 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_698 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_731 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_736 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_747 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_758 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_780 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_792 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_797 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_808 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_819 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_83 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_841 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_853 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_858 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_869 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_880 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_902 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_914 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_919 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_930 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_941 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_963 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_975 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_980 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_99 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_991 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_200_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_200_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_201_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_201_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_201_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_202_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_202_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_203_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_203_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_203_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_204_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_204_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_205_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_205_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_205_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_206_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_206_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_207_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_207_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_207_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_208_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_208_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_1028 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_103 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1036 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1054 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1059 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1071 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_1083 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_1089 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1097 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_209_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1118 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1146 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_115 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1158 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_1171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1179 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1183 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1195 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1207 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_121 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1219 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1224 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_209_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_1248 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_1267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_1275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_189 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_201 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_213 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_219 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_231 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_283 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_295 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_303 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_316 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_340 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_344 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_365 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_383 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_407 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_417 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_425 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_451 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_463 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_47 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_475 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_487 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_493 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_505 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_209_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_53 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_548 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_554 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_566 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_578 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_588 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_600 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_619 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_624 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_636 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_648 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_658 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_670 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_692 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_209_70 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_704 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_716 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_724 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_761 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_77 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_773 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_785 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_798 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_810 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_822 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_859 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_864 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_876 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_209_888 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_89 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_892 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_897 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_909 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_209_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_924 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_930 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_942 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_954 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_209_97 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_209_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_996 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_244 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_255 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_286 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_303 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_344 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_356 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_368 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_378 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_389 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_414 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_421 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_432 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_444 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_456 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_210_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_210_1126 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_210_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1149 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1161 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1173 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_210_1185 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_210_1189 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_210_1267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_210_1275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_210_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1005 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1017 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1024 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1036 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1048 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1055 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_106 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1067 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1079 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1098 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1148 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1179 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_118 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1210 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1222 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1234 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1241 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_125 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_1253 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_1265 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_211_1272 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_211_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_137 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_149 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_156 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_168 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_180 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_187 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_199 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_211 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_218 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_230 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_242 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_249 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_261 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_211_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_280 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_292 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_304 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_311 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_323 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_335 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_366 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_397 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_404 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_416 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_435 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_447 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_466 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_478 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_490 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_497 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_509 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_521 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_528 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_540 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_552 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_559 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_571 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_583 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_590 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_602 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_614 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_621 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_63 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_633 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_645 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_652 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_664 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_676 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_683 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_695 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_707 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_714 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_726 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_738 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_75 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_807 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_819 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_831 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_838 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_850 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_862 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_869 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_87 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_881 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_893 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_900 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_912 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_924 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_931 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_94 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_943 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_955 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_962 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_974 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_986 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_993 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_262 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_274 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_286 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_296 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_304 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_310 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_333 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_345 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_356 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_364 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_371 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_383 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_406 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_417 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_425 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_431 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_443 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_455 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_467 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_479 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_487 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_283 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_295 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_310 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_325 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_333 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_340 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_351 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_366 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_381 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_393 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_414 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_426 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_438 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_450 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_277 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_313 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_321 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_326 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_338 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_347 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_370 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_382 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_394 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_414 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_426 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_309 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_313 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_317 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_346 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_369 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_381 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_393 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_314 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_319 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_331 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_338 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_365 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_321 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_333 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_28_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_28_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_29_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_29_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_29_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1005 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1037 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1041 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1053 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_1065 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1073 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1085 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1089 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1101 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1109 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1125 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1136 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1148 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1152 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1164 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1176 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1188 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1224 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_1248 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_125 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1256 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_133 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_145 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_173 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_200 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_212 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_234 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_261 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_295 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_322 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_333 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_357 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_381 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_393 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_466 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_511 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_554 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_571 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_579 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_589 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_600 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_627 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_639 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_646 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_671 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_688 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_700 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_712 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_729 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_740 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_76 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_767 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_778 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_789 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_801 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_805 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_809 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_821 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_84 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_841 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_853 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_857 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_869 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_881 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_889 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_901 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_905 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_917 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_925 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_929 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_941 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_945 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_953 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_965 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_969 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_981 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_993 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_30_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_30_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_31_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_31_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_31_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_32_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_32_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_33_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_33_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_33_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_34_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_34_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_35_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_35_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_35_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_36_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_36_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_37_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_37_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_37_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_38_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_38_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_39_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_39_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_39_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_106 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_118 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_169 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_181 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_230 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_242 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_272 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_294 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_302 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_325 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_352 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_364 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_384 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_419 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_432 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_456 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_480 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_497 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_515 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_523 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_541 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_559 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_571 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_589 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_601 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_609 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_619 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_637 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_661 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_669 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_688 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_705 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_722 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_730 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_736 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_747 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_759 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_771 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_783 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_79 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_791 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_40_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_40_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_41_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_41_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_41_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_42_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_42_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_43_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_43_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_43_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_44_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_44_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_45_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_45_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_45_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_46_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_46_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_47_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_47_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_47_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_48_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_48_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_49_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_49_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_49_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_125 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_145 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_173 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_181 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_198 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_210 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_234 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_261 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_298 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_341 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_411 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_426 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_450 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_475 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_487 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_511 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_524 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_548 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_572 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_597 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_609 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_613 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_630 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_638 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_645 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_653 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_670 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_694 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_712 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_84 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_50_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_50_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_51_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_51_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_51_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_52_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_52_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_53_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_53_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_53_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_54_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_54_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_55_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_55_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_55_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_56_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_56_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_57_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_57_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_57_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_58_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_58_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_59_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_59_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_59_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_127 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_137 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_161 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_169 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_175 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_188 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_212 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_254 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_289 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_310 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_327 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_365 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_409 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_421 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_435 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_480 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_506 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_534 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_546 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_559 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_567 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_627 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_638 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_646 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_663 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_680 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_697 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_719 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_731 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_82 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_88 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_99 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_60_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_60_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_61_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_61_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_61_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_62_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_62_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_63_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_63_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_63_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_64_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_64_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_65_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_65_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_65_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_66_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_66_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_67_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_67_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_67_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_68_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_68_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_69_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_69_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_69_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_121 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_145 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_158 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_182 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_219 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_304 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_365 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_389 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_416 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_438 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_450 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_466 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_474 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_487 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_504 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_516 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_530 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_557 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_569 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_577 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_610 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_627 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_639 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_651 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_668 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_685 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_697 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_701 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_706 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_718 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_730 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_742 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_754 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_762 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_97 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_70_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_70_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_71_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_71_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_71_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_72_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_72_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_73_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_73_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_73_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_74_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_74_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_75_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_75_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_75_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_76_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_76_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_77_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_77_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_77_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_78_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_78_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_79_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_79_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_79_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_149 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_168 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_180 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_254 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_279 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_287 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_310 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_334 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_376 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_418 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_426 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_432 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_461 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_478 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_486 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_500 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_512 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_516 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_526 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_541 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_560 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_575 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_587 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_602 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_614 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_643 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_663 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_681 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_698 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_710 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_722 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_730 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_736 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_748 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_760 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_772 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_784 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_792 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_80_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_80_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_81_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_81_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_81_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_82_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_82_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_83_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_83_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_83_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_84_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_84_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_85_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_85_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_85_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_86_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_86_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_87_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_87_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_87_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_88_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_88_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_89_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_89_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_89_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_128 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_143 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_151 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_163 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_187 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_204 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_212 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_224 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_259 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_282 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_299 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_307 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_350 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_377 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_389 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_431 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_448 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_456 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_478 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_505 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_517 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_528 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_549 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_566 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_578 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_602 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_661 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_673 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_694 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_734 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_746 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_758 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_762 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_90_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_90_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_91_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_91_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_91_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_92_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_92_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_93_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_93_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_93_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_94_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_94_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_95_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_95_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_95_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_96_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_96_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_97_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_97_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_97_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1008 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1020 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1032 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1044 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1056 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1069 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1081 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1093 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_1264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_98_1276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_98_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_434 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_471 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_495 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_532 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_581 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_593 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_605 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_629 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_642 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_654 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_666 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_678 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_690 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_739 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_751 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_764 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_776 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_788 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_800 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_812 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_825 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_837 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_849 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_861 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_873 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_886 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_898 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_910 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_922 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_934 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_947 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_959 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_971 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_983 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_995 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_99_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_440 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_452 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_464 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_476 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_99_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_537 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_586 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_99_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_598 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_611 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_623 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_635 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_659 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_672 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_684 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_696 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_708 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_720 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1001 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1013 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1025 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1038 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1050 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1062 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1074 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1086 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1099 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_131 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_146 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_158 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_175 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_188 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_212 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_249 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_314 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_331 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_393 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_421 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_447 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_474 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_485 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_514 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_541 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_569 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_596 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_620 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_647 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_658 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_670 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_691 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_703 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_715 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_727 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_731 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_733 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_745 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_757 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_769 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_781 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_794 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_806 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_818 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_830 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_842 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_855 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_867 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_879 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_891 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_903 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_916 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_928 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_940 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_952 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_964 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_977 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_989 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_100 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_101 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_102 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_103 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_104 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_106 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_107 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_108 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_109 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_112 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_115 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_116 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_118 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_119 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_120 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_121 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_122 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_123 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_124 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_125 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_126 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_127 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_128 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_129 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_131 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_132 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_133 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_134 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_135 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_136 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_137 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_138 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_139 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_140 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_141 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_143 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_144 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_145 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_146 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_148 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_149 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_150 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_151 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_152 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_153 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_155 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_156 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_157 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_158 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_160 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_161 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_162 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_163 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_164 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_165 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_167 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_168 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_169 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_170 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_173 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_174 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_175 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_176 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_177 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_178 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_179 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_180 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_181 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_182 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_183 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_185 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_186 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_187 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_188 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_189 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_191 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_192 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_193 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_194 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_195 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_197 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_198 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_199 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_200 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_201 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_203 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_204 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_205 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_207 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_208 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_209 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_210 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_211 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_212 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_213 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_214 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_216 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_217 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_218 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_219 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_220 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_222 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_223 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_224 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_225 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_226 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_228 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_229 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_230 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_231 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_232 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_234 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_235 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_236 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_237 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_238 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_239 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_240 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_241 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_242 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_243 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_244 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_246 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_247 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_248 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_249 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_250 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_251 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_253 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_254 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_255 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_256 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_257 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_258 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_259 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_260 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_261 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_262 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_263 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_265 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_266 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_267 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_268 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_270 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_271 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_272 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_274 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_276 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_277 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_278 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_279 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_280 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_281 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_282 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_283 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_284 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_285 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_286 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_287 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_289 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_290 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_291 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_292 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_293 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_294 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_295 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_296 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_297 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_298 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_299 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_301 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_302 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_303 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_304 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_305 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_307 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_308 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_309 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_310 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_311 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_312 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_313 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_314 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_315 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_316 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_317 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_319 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_320 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_321 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_322 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_323 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_324 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_325 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_326 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_327 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_328 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_329 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_33 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_331 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_332 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_333 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_334 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_335 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_336 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_337 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_338 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_339 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_34 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_340 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_341 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_342 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_343 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_344 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_345 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_346 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_347 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_348 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_35 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_350 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_351 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_352 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_353 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_355 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_356 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_357 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_358 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_359 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_36 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_360 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_362 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_363 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_364 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_365 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_366 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_368 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_369 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_37 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_370 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_371 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_372 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_373 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_374 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_375 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_376 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_377 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_378 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_38 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_380 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_381 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_382 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_383 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_384 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_386 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_387 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_388 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_389 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_390 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_392 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_393 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_394 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_395 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_396 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_397 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_399 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_40 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_400 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_401 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4014 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4015 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4016 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4017 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4018 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4019 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4020 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4021 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4022 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4023 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4024 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4025 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4026 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4027 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4028 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4029 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_403 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4030 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4031 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4032 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4033 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4034 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4035 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4036 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4037 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4038 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4039 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_404 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4040 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4041 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4042 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4043 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4044 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4045 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4046 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4047 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4048 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4049 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_405 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4050 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4051 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4052 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4053 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4054 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4055 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4056 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4057 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4058 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4059 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_406 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4060 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4061 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4062 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4063 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4064 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4065 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4066 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4067 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4068 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4069 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_407 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4070 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4071 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4072 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4073 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4074 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4075 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4076 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4077 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4078 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4079 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_408 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4080 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4081 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4082 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4083 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4084 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4085 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4086 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4087 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4088 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4089 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_409 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4090 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4091 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4092 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4093 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4094 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4095 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4096 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4097 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4098 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4099 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_41 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_410 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4100 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4101 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4102 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4103 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4104 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4105 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4106 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4107 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4108 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4109 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_411 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4110 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4111 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4112 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4113 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4114 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4115 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4116 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4117 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4118 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4119 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_412 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4120 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4121 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4122 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4123 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4124 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4125 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4126 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4127 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4128 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4129 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_413 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4130 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4131 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4132 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4133 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4134 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4135 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4136 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4137 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4138 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4139 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_414 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4140 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4141 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4142 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4143 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4144 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4145 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4146 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4147 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4148 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4149 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_415 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4150 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4151 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4152 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4153 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4154 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4155 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4156 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4157 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4158 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4159 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_416 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4160 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4161 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4162 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4163 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4164 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4165 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4166 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4167 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4168 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4169 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_417 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4170 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4171 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4172 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4173 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4174 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4175 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4176 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4177 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4178 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4179 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_418 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4180 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4181 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4182 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4183 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4184 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4185 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4186 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4187 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4188 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4189 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_419 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4190 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4191 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4192 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4193 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4194 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4195 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4196 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4197 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4198 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4199 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_42 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_420 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4200 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4201 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4202 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4203 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4204 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4205 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4206 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4207 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4208 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4209 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_421 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4210 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4211 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4212 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4213 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4214 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4215 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4216 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4217 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4218 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4219 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_422 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4220 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4221 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4222 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4223 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4224 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4225 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4226 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4227 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4228 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4229 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_423 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4230 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4231 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4232 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4233 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4234 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4235 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4236 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4237 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4238 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4239 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4240 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4241 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4242 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4243 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4244 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4245 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4246 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4247 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4248 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4249 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4250 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4251 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4252 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4253 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4254 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4255 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4256 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4257 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4258 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4259 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4260 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4261 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4262 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4263 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4264 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4265 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4266 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4267 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4268 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4269 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4270 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4271 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4272 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4273 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4274 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4275 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4276 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4277 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4278 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4279 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4280 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4281 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4282 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4283 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4284 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4285 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4286 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4287 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4288 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4289 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4290 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4291 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4292 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4293 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4294 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4295 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4296 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4297 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4298 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4299 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_43 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4300 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4301 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4302 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4303 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4304 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4305 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4306 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4307 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4308 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4309 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4310 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4311 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4312 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4313 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4314 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4315 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4316 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4317 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4318 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4319 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4320 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4321 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4322 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4323 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4324 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4325 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4326 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4327 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4328 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4329 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4330 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4331 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4332 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4333 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4334 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4335 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4336 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4337 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4338 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4339 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4340 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4341 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4342 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4343 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4344 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4345 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4346 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4347 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4348 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4349 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4350 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4351 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4352 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4353 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4354 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4355 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4356 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4357 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4358 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4359 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4360 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4361 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4362 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4363 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4364 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4365 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4366 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4367 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4368 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4369 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4370 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4371 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4372 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4373 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4374 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4375 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4376 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4377 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4378 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4379 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4380 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4381 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4382 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4383 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4384 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4385 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4386 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4387 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4388 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4389 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4390 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4391 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4392 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4393 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4394 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4395 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4396 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4397 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4398 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4399 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4400 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4401 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4402 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4403 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4404 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4405 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4406 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4407 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4408 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4409 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4410 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4411 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4412 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4413 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4414 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4415 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4416 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4417 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4418 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4419 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4420 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4421 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4422 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4423 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4424 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4425 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4426 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4427 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4428 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4429 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4430 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4431 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4432 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4433 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4434 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4435 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4436 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4437 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4438 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4439 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4440 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4441 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4442 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4443 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4444 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4445 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4446 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4447 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4448 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4449 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4450 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4451 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4452 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4453 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4454 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4455 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4456 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4457 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4458 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4459 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4460 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4461 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4462 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4463 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4464 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4465 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4466 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4467 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4468 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4469 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4470 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4471 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4472 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4473 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4474 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4475 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4476 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4477 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4478 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4479 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4480 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4481 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4482 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4483 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4484 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4485 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4486 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4487 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4488 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4489 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4490 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4491 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4492 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4493 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4494 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4495 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4496 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4497 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4498 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4499 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_45 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4500 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4501 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4502 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4503 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4504 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4505 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4506 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4507 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4508 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4509 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4510 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4511 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4512 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4513 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4514 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4515 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4516 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4517 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4518 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4519 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4520 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4521 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4522 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4523 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4524 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4525 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4526 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4527 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4528 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4529 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4530 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4531 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4532 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4533 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4534 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4535 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4536 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4537 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4538 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4539 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4540 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4541 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4542 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4543 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4544 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4545 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4546 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4547 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4548 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4549 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4550 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4551 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4552 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4553 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4554 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4555 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4556 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4557 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4558 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4559 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4560 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4561 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4562 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4563 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4564 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4565 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4566 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4567 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4568 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4569 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4570 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4571 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4572 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4573 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4574 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4575 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4576 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4577 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4578 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4579 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4580 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4581 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4582 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4583 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4584 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4585 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4586 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4587 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4588 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4589 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4590 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4591 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4592 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4593 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4594 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4595 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4596 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4597 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4598 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4599 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_46 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4600 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4601 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4602 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4603 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4604 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4605 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4606 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4607 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4608 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4609 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4610 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4611 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4612 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4613 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4614 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4615 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4616 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4617 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4618 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4619 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4620 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4621 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4622 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4623 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4624 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4625 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4626 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4627 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4628 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4629 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4630 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4631 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4632 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4633 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4634 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4635 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4636 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4637 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4638 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4639 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4640 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4641 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4642 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4643 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4644 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4645 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4646 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4647 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4648 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4649 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4650 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4651 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4652 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4653 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4654 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4655 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4656 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4657 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4658 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4659 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4660 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4661 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4662 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4663 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4664 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4665 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4666 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4667 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4668 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4669 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4670 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4671 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4672 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4673 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4674 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4675 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4676 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4677 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4678 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4679 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4680 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4681 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4682 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4683 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4684 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4685 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4686 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4687 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4688 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4689 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4690 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4691 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4692 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4693 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4694 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4695 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4696 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4697 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4698 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4699 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_47 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4700 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4701 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4702 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4703 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4704 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4705 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4706 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4707 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4708 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4709 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4710 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4711 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4712 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4713 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4714 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4715 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4716 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4717 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4718 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4719 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4720 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4721 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4722 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4723 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4724 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4725 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4726 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4727 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4728 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4729 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4730 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4731 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4732 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4733 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4734 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4735 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4736 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4737 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4738 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4739 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4740 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4741 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4742 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4743 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4744 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4745 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4746 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4747 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4748 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4749 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4750 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4751 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4752 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4753 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4754 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4755 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4756 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4757 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4758 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4759 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4760 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4761 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4762 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4763 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4764 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4765 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4766 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4767 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4768 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4769 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4770 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4771 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4772 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4773 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4774 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4775 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4776 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4777 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4778 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4779 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4780 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4781 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4782 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4783 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4784 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4785 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4786 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4787 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4788 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4789 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4790 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4791 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4792 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4793 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4794 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4795 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4796 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4797 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4798 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4799 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_48 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4800 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4801 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4802 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4803 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4804 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4805 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4806 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4807 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4808 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4809 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4810 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_49 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_50 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_52 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_53 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_54 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_55 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_57 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_58 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_60 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_61 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_63 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_64 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_65 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_66 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_67 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_69 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_70 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_71 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_72 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_73 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_75 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_76 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_77 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_78 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_79 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_81 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_82 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_83 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_84 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_85 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_87 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_88 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_89 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_90 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_92 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_94 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_95 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_96 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_97 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_99 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__inv_2 _0402_ (
    .A(la_oen[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0097_)
  );
  sky130_fd_sc_hd__o22a_4 _0403_ (
    .A1(la_data_in[65]),
    .A2(la_oen[65]),
    .B1(wb_rst_i),
    .B2(_0097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0098_)
  );
  sky130_fd_sc_hd__buf_2 _0404_ (
    .A(_0098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0099_)
  );
  sky130_fd_sc_hd__buf_4 _0405_ (
    .A(_0099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[36])
  );
  sky130_fd_sc_hd__inv_2 _0406_ (
    .A(_0099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0100_)
  );
  sky130_fd_sc_hd__buf_2 _0407_ (
    .A(_0100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0101_)
  );
  sky130_fd_sc_hd__and2_4 _0408_ (
    .A(wbs_stb_i),
    .B(wbs_cyc_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0102_)
  );
  sky130_fd_sc_hd__buf_2 _0409_ (
    .A(_0102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0103_)
  );
  sky130_fd_sc_hd__buf_2 _0410_ (
    .A(_0103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0104_)
  );
  sky130_fd_sc_hd__buf_2 _0411_ (
    .A(_0104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0105_)
  );
  sky130_fd_sc_hd__inv_2 _0412_ (
    .A(_0105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0106_)
  );
  sky130_fd_sc_hd__inv_2 _0413_ (
    .A(wbs_we_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0107_)
  );
  sky130_fd_sc_hd__inv_2 _0414_ (
    .A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0108_)
  );
  sky130_fd_sc_hd__or4_4 _0415_ (
    .A(wbs_ack_o),
    .B(_0106_),
    .C(_0107_),
    .D(_0108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0109_)
  );
  sky130_fd_sc_hd__buf_2 _0416_ (
    .A(_0109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0110_)
  );
  sky130_fd_sc_hd__or2_4 _0417_ (
    .A(wbs_dat_i[30]),
    .B(_0110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0111_)
  );
  sky130_fd_sc_hd__inv_2 _0418_ (
    .A(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0112_)
  );
  sky130_fd_sc_hd__inv_2 _0419_ (
    .A(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0113_)
  );
  sky130_fd_sc_hd__inv_2 _0420_ (
    .A(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0114_)
  );
  sky130_fd_sc_hd__inv_2 _0421_ (
    .A(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0115_)
  );
  sky130_fd_sc_hd__inv_2 _0422_ (
    .A(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0116_)
  );
  sky130_fd_sc_hd__inv_2 _0423_ (
    .A(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0117_)
  );
  sky130_fd_sc_hd__inv_2 _0424_ (
    .A(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0118_)
  );
  sky130_fd_sc_hd__or2_4 _0425_ (
    .A(_0117_),
    .B(_0118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0119_)
  );
  sky130_fd_sc_hd__inv_2 _0426_ (
    .A(io_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0120_)
  );
  sky130_fd_sc_hd__inv_2 _0427_ (
    .A(io_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0121_)
  );
  sky130_fd_sc_hd__inv_2 _0428_ (
    .A(io_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0122_)
  );
  sky130_fd_sc_hd__inv_2 _0429_ (
    .A(io_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0123_)
  );
  sky130_fd_sc_hd__or4_4 _0430_ (
    .A(_0120_),
    .B(_0121_),
    .C(_0122_),
    .D(_0123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0124_)
  );
  sky130_fd_sc_hd__inv_2 _0431_ (
    .A(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0125_)
  );
  sky130_fd_sc_hd__inv_2 _0432_ (
    .A(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0126_)
  );
  sky130_fd_sc_hd__inv_2 _0433_ (
    .A(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0127_)
  );
  sky130_fd_sc_hd__inv_2 _0434_ (
    .A(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0128_)
  );
  sky130_fd_sc_hd__or4_4 _0435_ (
    .A(_0125_),
    .B(_0126_),
    .C(_0127_),
    .D(_0128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0129_)
  );
  sky130_fd_sc_hd__inv_2 _0436_ (
    .A(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0130_)
  );
  sky130_fd_sc_hd__inv_2 _0437_ (
    .A(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0131_)
  );
  sky130_fd_sc_hd__inv_2 _0438_ (
    .A(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0132_)
  );
  sky130_fd_sc_hd__inv_2 _0439_ (
    .A(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0133_)
  );
  sky130_fd_sc_hd__or2_4 _0440_ (
    .A(_0132_),
    .B(_0133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0134_)
  );
  sky130_fd_sc_hd__inv_2 _0441_ (
    .A(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0135_)
  );
  sky130_fd_sc_hd__inv_2 _0442_ (
    .A(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0136_)
  );
  sky130_fd_sc_hd__inv_2 _0443_ (
    .A(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0137_)
  );
  sky130_fd_sc_hd__inv_2 _0444_ (
    .A(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0138_)
  );
  sky130_fd_sc_hd__or4_4 _0445_ (
    .A(_0135_),
    .B(_0136_),
    .C(_0137_),
    .D(_0138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0139_)
  );
  sky130_fd_sc_hd__or4_4 _0446_ (
    .A(_0130_),
    .B(_0131_),
    .C(_0134_),
    .D(_0139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0140_)
  );
  sky130_fd_sc_hd__inv_2 _0447_ (
    .A(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0141_)
  );
  sky130_fd_sc_hd__inv_2 _0448_ (
    .A(io_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0142_)
  );
  sky130_fd_sc_hd__inv_2 _0449_ (
    .A(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0143_)
  );
  sky130_fd_sc_hd__or2_4 _0450_ (
    .A(_0142_),
    .B(_0143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0144_)
  );
  sky130_fd_sc_hd__inv_2 _0451_ (
    .A(io_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0145_)
  );
  sky130_fd_sc_hd__inv_2 _0452_ (
    .A(io_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0146_)
  );
  sky130_fd_sc_hd__inv_2 _0453_ (
    .A(io_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0147_)
  );
  sky130_fd_sc_hd__inv_2 _0454_ (
    .A(io_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0148_)
  );
  sky130_fd_sc_hd__inv_2 _0455_ (
    .A(io_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0149_)
  );
  sky130_fd_sc_hd__or4_4 _0456_ (
    .A(_0146_),
    .B(_0147_),
    .C(_0148_),
    .D(_0149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0150_)
  );
  sky130_fd_sc_hd__or4_4 _0457_ (
    .A(_0141_),
    .B(_0144_),
    .C(_0145_),
    .D(_0150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0151_)
  );
  sky130_fd_sc_hd__or2_4 _0458_ (
    .A(_0140_),
    .B(_0151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0152_)
  );
  sky130_fd_sc_hd__nor2_4 _0459_ (
    .A(la_oen[32]),
    .B(_0104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0153_)
  );
  sky130_fd_sc_hd__nor2_4 _0460_ (
    .A(la_oen[34]),
    .B(_0104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0154_)
  );
  sky130_fd_sc_hd__buf_2 _0461_ (
    .A(_0103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0155_)
  );
  sky130_fd_sc_hd__nor2_4 _0462_ (
    .A(la_oen[35]),
    .B(_0155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0156_)
  );
  sky130_fd_sc_hd__buf_2 _0463_ (
    .A(_0103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0157_)
  );
  sky130_fd_sc_hd__nor2_4 _0464_ (
    .A(la_oen[33]),
    .B(_0157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0158_)
  );
  sky130_fd_sc_hd__or4_4 _0465_ (
    .A(_0153_),
    .B(_0154_),
    .C(_0156_),
    .D(_0158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0159_)
  );
  sky130_fd_sc_hd__nor2_4 _0466_ (
    .A(la_oen[36]),
    .B(_0104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0160_)
  );
  sky130_fd_sc_hd__nor2_4 _0467_ (
    .A(la_oen[38]),
    .B(_0155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0161_)
  );
  sky130_fd_sc_hd__buf_2 _0468_ (
    .A(_0103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0162_)
  );
  sky130_fd_sc_hd__nor2_4 _0469_ (
    .A(la_oen[39]),
    .B(_0162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0163_)
  );
  sky130_fd_sc_hd__nor2_4 _0470_ (
    .A(la_oen[37]),
    .B(_0157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0164_)
  );
  sky130_fd_sc_hd__or4_4 _0471_ (
    .A(_0160_),
    .B(_0161_),
    .C(_0163_),
    .D(_0164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0165_)
  );
  sky130_fd_sc_hd__nor2_4 _0472_ (
    .A(la_oen[40]),
    .B(_0162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0166_)
  );
  sky130_fd_sc_hd__nor2_4 _0473_ (
    .A(la_oen[42]),
    .B(_0162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0167_)
  );
  sky130_fd_sc_hd__buf_2 _0474_ (
    .A(_0103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0168_)
  );
  sky130_fd_sc_hd__nor2_4 _0475_ (
    .A(la_oen[43]),
    .B(_0168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0169_)
  );
  sky130_fd_sc_hd__buf_2 _0476_ (
    .A(_0104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0170_)
  );
  sky130_fd_sc_hd__nor2_4 _0477_ (
    .A(la_oen[41]),
    .B(_0170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0171_)
  );
  sky130_fd_sc_hd__or4_4 _0478_ (
    .A(_0166_),
    .B(_0167_),
    .C(_0169_),
    .D(_0171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0172_)
  );
  sky130_fd_sc_hd__nor2_4 _0479_ (
    .A(la_oen[44]),
    .B(_0157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0173_)
  );
  sky130_fd_sc_hd__nor2_4 _0480_ (
    .A(la_oen[46]),
    .B(_0157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0174_)
  );
  sky130_fd_sc_hd__nor2_4 _0481_ (
    .A(la_oen[47]),
    .B(_0170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0175_)
  );
  sky130_fd_sc_hd__nor2_4 _0482_ (
    .A(la_oen[45]),
    .B(_0105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0176_)
  );
  sky130_fd_sc_hd__or4_4 _0483_ (
    .A(_0173_),
    .B(_0174_),
    .C(_0175_),
    .D(_0176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0177_)
  );
  sky130_fd_sc_hd__or4_4 _0484_ (
    .A(_0159_),
    .B(_0165_),
    .C(_0172_),
    .D(_0177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0178_)
  );
  sky130_fd_sc_hd__nor2_4 _0485_ (
    .A(la_oen[48]),
    .B(_0155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0179_)
  );
  sky130_fd_sc_hd__nor2_4 _0486_ (
    .A(la_oen[50]),
    .B(_0155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0180_)
  );
  sky130_fd_sc_hd__nor2_4 _0487_ (
    .A(la_oen[51]),
    .B(_0162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0181_)
  );
  sky130_fd_sc_hd__nor2_4 _0488_ (
    .A(la_oen[49]),
    .B(_0170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0182_)
  );
  sky130_fd_sc_hd__or4_4 _0489_ (
    .A(_0179_),
    .B(_0180_),
    .C(_0181_),
    .D(_0182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0183_)
  );
  sky130_fd_sc_hd__nor2_4 _0490_ (
    .A(la_oen[52]),
    .B(_0155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0184_)
  );
  sky130_fd_sc_hd__nor2_4 _0491_ (
    .A(la_oen[54]),
    .B(_0162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0185_)
  );
  sky130_fd_sc_hd__nor2_4 _0492_ (
    .A(la_oen[55]),
    .B(_0168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0186_)
  );
  sky130_fd_sc_hd__nor2_4 _0493_ (
    .A(la_oen[53]),
    .B(_0170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0187_)
  );
  sky130_fd_sc_hd__or4_4 _0494_ (
    .A(_0184_),
    .B(_0185_),
    .C(_0186_),
    .D(_0187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0188_)
  );
  sky130_fd_sc_hd__nor2_4 _0495_ (
    .A(la_oen[56]),
    .B(_0168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0189_)
  );
  sky130_fd_sc_hd__nor2_4 _0496_ (
    .A(la_oen[58]),
    .B(_0168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0190_)
  );
  sky130_fd_sc_hd__nor2_4 _0497_ (
    .A(la_oen[59]),
    .B(_0168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0191_)
  );
  sky130_fd_sc_hd__nor2_4 _0498_ (
    .A(la_oen[57]),
    .B(_0105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0192_)
  );
  sky130_fd_sc_hd__or4_4 _0499_ (
    .A(_0189_),
    .B(_0190_),
    .C(_0191_),
    .D(_0192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0193_)
  );
  sky130_fd_sc_hd__nor2_4 _0500_ (
    .A(la_oen[60]),
    .B(_0157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0194_)
  );
  sky130_fd_sc_hd__nor2_4 _0501_ (
    .A(la_oen[62]),
    .B(_0170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0195_)
  );
  sky130_fd_sc_hd__nor2_4 _0502_ (
    .A(la_oen[63]),
    .B(_0105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0196_)
  );
  sky130_fd_sc_hd__nor2_4 _0503_ (
    .A(la_oen[61]),
    .B(_0105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0197_)
  );
  sky130_fd_sc_hd__or4_4 _0504_ (
    .A(_0194_),
    .B(_0195_),
    .C(_0196_),
    .D(_0197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0198_)
  );
  sky130_fd_sc_hd__or4_4 _0505_ (
    .A(_0183_),
    .B(_0188_),
    .C(_0193_),
    .D(_0198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0199_)
  );
  sky130_fd_sc_hd__or2_4 _0506_ (
    .A(_0178_),
    .B(_0199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0200_)
  );
  sky130_fd_sc_hd__or4_4 _0507_ (
    .A(_0124_),
    .B(_0129_),
    .C(_0152_),
    .D(_0200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0201_)
  );
  sky130_fd_sc_hd__or4_4 _0508_ (
    .A(_0115_),
    .B(_0116_),
    .C(_0119_),
    .D(_0201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0202_)
  );
  sky130_fd_sc_hd__or3_4 _0509_ (
    .A(_0113_),
    .B(_0114_),
    .C(_0202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0203_)
  );
  sky130_fd_sc_hd__nand2_4 _0510_ (
    .A(_0112_),
    .B(_0203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0204_)
  );
  sky130_fd_sc_hd__or2_4 _0511_ (
    .A(_0112_),
    .B(_0203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0205_)
  );
  sky130_fd_sc_hd__buf_2 _0512_ (
    .A(_0109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0206_)
  );
  sky130_fd_sc_hd__inv_2 _0513_ (
    .A(_0206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0207_)
  );
  sky130_fd_sc_hd__a21o_4 _0514_ (
    .A1(_0204_),
    .A2(_0205_),
    .B1(_0207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0208_)
  );
  sky130_fd_sc_hd__and3_4 _0515_ (
    .A(_0101_),
    .B(_0111_),
    .C(_0208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0095_)
  );
  sky130_fd_sc_hd__buf_2 _0516_ (
    .A(_0206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0209_)
  );
  sky130_fd_sc_hd__nor2_4 _0517_ (
    .A(_0114_),
    .B(_0202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0210_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0518_ (
    .A1_N(io_out[29]),
    .A2_N(_0210_),
    .B1(io_out[29]),
    .B2(_0210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0211_)
  );
  sky130_fd_sc_hd__nor2_4 _0519_ (
    .A(wbs_dat_i[29]),
    .B(_0110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0212_)
  );
  sky130_fd_sc_hd__a211o_4 _0520_ (
    .A1(_0209_),
    .A2(_0211_),
    .B1(io_oeb[36]),
    .C1(_0212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0213_)
  );
  sky130_fd_sc_hd__inv_2 _0521_ (
    .A(_0213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0094_)
  );
  sky130_fd_sc_hd__or2_4 _0522_ (
    .A(wbs_dat_i[28]),
    .B(_0110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0214_)
  );
  sky130_fd_sc_hd__and2_4 _0523_ (
    .A(_0114_),
    .B(_0202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0215_)
  );
  sky130_fd_sc_hd__o21ai_4 _0524_ (
    .A1(_0210_),
    .A2(_0215_),
    .B1(_0209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0216_)
  );
  sky130_fd_sc_hd__and3_4 _0525_ (
    .A(_0101_),
    .B(_0214_),
    .C(_0216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0093_)
  );
  sky130_fd_sc_hd__or3_4 _0526_ (
    .A(_0115_),
    .B(_0116_),
    .C(_0201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0217_)
  );
  sky130_fd_sc_hd__inv_2 _0527_ (
    .A(_0217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0218_)
  );
  sky130_fd_sc_hd__or2_4 _0528_ (
    .A(_0118_),
    .B(_0217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0219_)
  );
  sky130_fd_sc_hd__a32o_4 _0529_ (
    .A1(io_out[26]),
    .A2(_0218_),
    .A3(io_out[27]),
    .B1(_0117_),
    .B2(_0219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0220_)
  );
  sky130_fd_sc_hd__nor2_4 _0530_ (
    .A(wbs_dat_i[27]),
    .B(_0110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0221_)
  );
  sky130_fd_sc_hd__a211o_4 _0531_ (
    .A1(_0209_),
    .A2(_0220_),
    .B1(io_oeb[36]),
    .C1(_0221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0222_)
  );
  sky130_fd_sc_hd__inv_2 _0532_ (
    .A(_0222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0092_)
  );
  sky130_fd_sc_hd__buf_2 _0533_ (
    .A(_0100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0223_)
  );
  sky130_fd_sc_hd__or2_4 _0534_ (
    .A(io_out[26]),
    .B(_0218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0224_)
  );
  sky130_fd_sc_hd__a32o_4 _0535_ (
    .A1(_0206_),
    .A2(_0219_),
    .A3(_0224_),
    .B1(wbs_dat_i[26]),
    .B2(_0207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0225_)
  );
  sky130_fd_sc_hd__and2_4 _0536_ (
    .A(_0223_),
    .B(_0225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0091_)
  );
  sky130_fd_sc_hd__nor2_4 _0537_ (
    .A(_0116_),
    .B(_0201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0226_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0538_ (
    .A1_N(io_out[25]),
    .A2_N(_0226_),
    .B1(io_out[25]),
    .B2(_0226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0227_)
  );
  sky130_fd_sc_hd__nor2_4 _0539_ (
    .A(wbs_dat_i[25]),
    .B(_0110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0228_)
  );
  sky130_fd_sc_hd__a211o_4 _0540_ (
    .A1(_0209_),
    .A2(_0227_),
    .B1(io_oeb[36]),
    .C1(_0228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0229_)
  );
  sky130_fd_sc_hd__inv_2 _0541_ (
    .A(_0229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0090_)
  );
  sky130_fd_sc_hd__or2_4 _0542_ (
    .A(wbs_dat_i[24]),
    .B(_0206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0230_)
  );
  sky130_fd_sc_hd__and2_4 _0543_ (
    .A(_0116_),
    .B(_0201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0231_)
  );
  sky130_fd_sc_hd__o21ai_4 _0544_ (
    .A1(_0226_),
    .A2(_0231_),
    .B1(_0209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0232_)
  );
  sky130_fd_sc_hd__and3_4 _0545_ (
    .A(_0101_),
    .B(_0230_),
    .C(_0232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0089_)
  );
  sky130_fd_sc_hd__inv_2 _0546_ (
    .A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0233_)
  );
  sky130_fd_sc_hd__or4_4 _0547_ (
    .A(wbs_ack_o),
    .B(_0106_),
    .C(_0107_),
    .D(_0233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0234_)
  );
  sky130_fd_sc_hd__buf_2 _0548_ (
    .A(_0234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0235_)
  );
  sky130_fd_sc_hd__or2_4 _0549_ (
    .A(wbs_dat_i[23]),
    .B(_0235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0236_)
  );
  sky130_fd_sc_hd__or2_4 _0550_ (
    .A(_0200_),
    .B(_0152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0237_)
  );
  sky130_fd_sc_hd__or2_4 _0551_ (
    .A(_0124_),
    .B(_0237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0238_)
  );
  sky130_fd_sc_hd__or3_4 _0552_ (
    .A(_0125_),
    .B(_0126_),
    .C(_0238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0239_)
  );
  sky130_fd_sc_hd__or2_4 _0553_ (
    .A(_0128_),
    .B(_0239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0240_)
  );
  sky130_fd_sc_hd__buf_2 _0554_ (
    .A(_0234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0241_)
  );
  sky130_fd_sc_hd__inv_2 _0555_ (
    .A(_0241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0242_)
  );
  sky130_fd_sc_hd__nor2_4 _0556_ (
    .A(io_out[23]),
    .B(_0240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0243_)
  );
  sky130_fd_sc_hd__a211o_4 _0557_ (
    .A1(io_out[23]),
    .A2(_0240_),
    .B1(_0242_),
    .C1(_0243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0244_)
  );
  sky130_fd_sc_hd__and3_4 _0558_ (
    .A(_0101_),
    .B(_0236_),
    .C(_0244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0088_)
  );
  sky130_fd_sc_hd__or2_4 _0559_ (
    .A(wbs_dat_i[22]),
    .B(_0235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0245_)
  );
  sky130_fd_sc_hd__nand2_4 _0560_ (
    .A(_0128_),
    .B(_0239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0246_)
  );
  sky130_fd_sc_hd__a21o_4 _0561_ (
    .A1(_0240_),
    .A2(_0246_),
    .B1(_0242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0247_)
  );
  sky130_fd_sc_hd__and3_4 _0562_ (
    .A(_0101_),
    .B(_0245_),
    .C(_0247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0087_)
  );
  sky130_fd_sc_hd__buf_2 _0563_ (
    .A(_0241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0248_)
  );
  sky130_fd_sc_hd__nor2_4 _0564_ (
    .A(_0126_),
    .B(_0238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0249_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0565_ (
    .A1_N(io_out[21]),
    .A2_N(_0249_),
    .B1(io_out[21]),
    .B2(_0249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0250_)
  );
  sky130_fd_sc_hd__nor2_4 _0566_ (
    .A(wbs_dat_i[21]),
    .B(_0235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0251_)
  );
  sky130_fd_sc_hd__a211o_4 _0567_ (
    .A1(_0248_),
    .A2(_0250_),
    .B1(io_oeb[36]),
    .C1(_0251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0252_)
  );
  sky130_fd_sc_hd__inv_2 _0568_ (
    .A(_0252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0086_)
  );
  sky130_fd_sc_hd__buf_2 _0569_ (
    .A(_0100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0253_)
  );
  sky130_fd_sc_hd__or2_4 _0570_ (
    .A(wbs_dat_i[20]),
    .B(_0241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0254_)
  );
  sky130_fd_sc_hd__and2_4 _0571_ (
    .A(_0126_),
    .B(_0238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0255_)
  );
  sky130_fd_sc_hd__o21ai_4 _0572_ (
    .A1(_0249_),
    .A2(_0255_),
    .B1(_0248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0256_)
  );
  sky130_fd_sc_hd__and3_4 _0573_ (
    .A(_0253_),
    .B(_0254_),
    .C(_0256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0085_)
  );
  sky130_fd_sc_hd__buf_2 _0574_ (
    .A(_0200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0257_)
  );
  sky130_fd_sc_hd__or4_4 _0575_ (
    .A(_0120_),
    .B(_0121_),
    .C(_0257_),
    .D(_0152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0258_)
  );
  sky130_fd_sc_hd__inv_2 _0576_ (
    .A(_0258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0259_)
  );
  sky130_fd_sc_hd__or2_4 _0577_ (
    .A(_0123_),
    .B(_0258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0260_)
  );
  sky130_fd_sc_hd__a32o_4 _0578_ (
    .A1(io_out[18]),
    .A2(_0259_),
    .A3(io_out[19]),
    .B1(_0122_),
    .B2(_0260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0261_)
  );
  sky130_fd_sc_hd__buf_2 _0579_ (
    .A(_0099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0262_)
  );
  sky130_fd_sc_hd__nor2_4 _0580_ (
    .A(wbs_dat_i[19]),
    .B(_0235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0263_)
  );
  sky130_fd_sc_hd__a211o_4 _0581_ (
    .A1(_0248_),
    .A2(_0261_),
    .B1(_0262_),
    .C1(_0263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0264_)
  );
  sky130_fd_sc_hd__inv_2 _0582_ (
    .A(_0264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0084_)
  );
  sky130_fd_sc_hd__or2_4 _0583_ (
    .A(io_out[18]),
    .B(_0259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0265_)
  );
  sky130_fd_sc_hd__a32o_4 _0584_ (
    .A1(_0241_),
    .A2(_0260_),
    .A3(_0265_),
    .B1(wbs_dat_i[18]),
    .B2(_0242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0266_)
  );
  sky130_fd_sc_hd__and2_4 _0585_ (
    .A(_0223_),
    .B(_0266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0083_)
  );
  sky130_fd_sc_hd__nor2_4 _0586_ (
    .A(_0121_),
    .B(_0237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0267_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0587_ (
    .A1_N(io_out[17]),
    .A2_N(_0267_),
    .B1(io_out[17]),
    .B2(_0267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0268_)
  );
  sky130_fd_sc_hd__nor2_4 _0588_ (
    .A(wbs_dat_i[17]),
    .B(_0235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0269_)
  );
  sky130_fd_sc_hd__a211o_4 _0589_ (
    .A1(_0248_),
    .A2(_0268_),
    .B1(_0262_),
    .C1(_0269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0270_)
  );
  sky130_fd_sc_hd__inv_2 _0590_ (
    .A(_0270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0082_)
  );
  sky130_fd_sc_hd__or2_4 _0591_ (
    .A(wbs_dat_i[16]),
    .B(_0241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0271_)
  );
  sky130_fd_sc_hd__and2_4 _0592_ (
    .A(_0121_),
    .B(_0237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0272_)
  );
  sky130_fd_sc_hd__o21ai_4 _0593_ (
    .A1(_0267_),
    .A2(_0272_),
    .B1(_0248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0273_)
  );
  sky130_fd_sc_hd__and3_4 _0594_ (
    .A(_0253_),
    .B(_0271_),
    .C(_0273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0081_)
  );
  sky130_fd_sc_hd__inv_2 _0595_ (
    .A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0274_)
  );
  sky130_fd_sc_hd__or4_4 _0596_ (
    .A(wbs_ack_o),
    .B(_0106_),
    .C(_0107_),
    .D(_0274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0275_)
  );
  sky130_fd_sc_hd__buf_2 _0597_ (
    .A(_0275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0276_)
  );
  sky130_fd_sc_hd__or2_4 _0598_ (
    .A(wbs_dat_i[15]),
    .B(_0276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0277_)
  );
  sky130_fd_sc_hd__buf_2 _0599_ (
    .A(_0275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0278_)
  );
  sky130_fd_sc_hd__inv_2 _0600_ (
    .A(_0278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0279_)
  );
  sky130_fd_sc_hd__or2_4 _0601_ (
    .A(_0200_),
    .B(_0140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0280_)
  );
  sky130_fd_sc_hd__or2_4 _0602_ (
    .A(_0150_),
    .B(_0280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0281_)
  );
  sky130_fd_sc_hd__or4_4 _0603_ (
    .A(_0142_),
    .B(_0143_),
    .C(_0141_),
    .D(_0281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0282_)
  );
  sky130_fd_sc_hd__inv_2 _0604_ (
    .A(_0282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0283_)
  );
  sky130_fd_sc_hd__o22a_4 _0605_ (
    .A1(io_out[15]),
    .A2(_0283_),
    .B1(_0151_),
    .B2(_0280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0284_)
  );
  sky130_fd_sc_hd__or2_4 _0606_ (
    .A(_0279_),
    .B(_0284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0285_)
  );
  sky130_fd_sc_hd__and3_4 _0607_ (
    .A(_0253_),
    .B(_0277_),
    .C(_0285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0080_)
  );
  sky130_fd_sc_hd__buf_2 _0608_ (
    .A(_0278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0286_)
  );
  sky130_fd_sc_hd__or2_4 _0609_ (
    .A(_0141_),
    .B(_0281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0287_)
  );
  sky130_fd_sc_hd__or2_4 _0610_ (
    .A(_0143_),
    .B(_0287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0288_)
  );
  sky130_fd_sc_hd__a21o_4 _0611_ (
    .A1(_0142_),
    .A2(_0288_),
    .B1(_0283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0289_)
  );
  sky130_fd_sc_hd__nor2_4 _0612_ (
    .A(wbs_dat_i[14]),
    .B(_0276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0290_)
  );
  sky130_fd_sc_hd__a211o_4 _0613_ (
    .A1(_0286_),
    .A2(_0289_),
    .B1(_0262_),
    .C1(_0290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0291_)
  );
  sky130_fd_sc_hd__inv_2 _0614_ (
    .A(_0291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0079_)
  );
  sky130_fd_sc_hd__inv_2 _0615_ (
    .A(_0287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0292_)
  );
  sky130_fd_sc_hd__or2_4 _0616_ (
    .A(io_out[13]),
    .B(_0292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0293_)
  );
  sky130_fd_sc_hd__a32o_4 _0617_ (
    .A1(_0278_),
    .A2(_0288_),
    .A3(_0293_),
    .B1(wbs_dat_i[13]),
    .B2(_0279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0294_)
  );
  sky130_fd_sc_hd__and2_4 _0618_ (
    .A(_0223_),
    .B(_0294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0078_)
  );
  sky130_fd_sc_hd__or2_4 _0619_ (
    .A(wbs_dat_i[12]),
    .B(_0276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0295_)
  );
  sky130_fd_sc_hd__and2_4 _0620_ (
    .A(_0141_),
    .B(_0281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0296_)
  );
  sky130_fd_sc_hd__o21ai_4 _0621_ (
    .A1(_0292_),
    .A2(_0296_),
    .B1(_0286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0297_)
  );
  sky130_fd_sc_hd__and3_4 _0622_ (
    .A(_0253_),
    .B(_0295_),
    .C(_0297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0077_)
  );
  sky130_fd_sc_hd__or4_4 _0623_ (
    .A(_0146_),
    .B(_0147_),
    .C(_0257_),
    .D(_0140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0298_)
  );
  sky130_fd_sc_hd__inv_2 _0624_ (
    .A(_0298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0299_)
  );
  sky130_fd_sc_hd__or2_4 _0625_ (
    .A(_0149_),
    .B(_0298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0300_)
  );
  sky130_fd_sc_hd__a32o_4 _0626_ (
    .A1(io_out[10]),
    .A2(_0299_),
    .A3(io_out[11]),
    .B1(_0148_),
    .B2(_0300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0301_)
  );
  sky130_fd_sc_hd__nor2_4 _0627_ (
    .A(wbs_dat_i[11]),
    .B(_0276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0302_)
  );
  sky130_fd_sc_hd__a211o_4 _0628_ (
    .A1(_0286_),
    .A2(_0301_),
    .B1(_0262_),
    .C1(_0302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0303_)
  );
  sky130_fd_sc_hd__inv_2 _0629_ (
    .A(_0303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0076_)
  );
  sky130_fd_sc_hd__or2_4 _0630_ (
    .A(io_out[10]),
    .B(_0299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0304_)
  );
  sky130_fd_sc_hd__a32o_4 _0631_ (
    .A1(_0278_),
    .A2(_0300_),
    .A3(_0304_),
    .B1(wbs_dat_i[10]),
    .B2(_0279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0305_)
  );
  sky130_fd_sc_hd__and2_4 _0632_ (
    .A(_0223_),
    .B(_0305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0075_)
  );
  sky130_fd_sc_hd__nor2_4 _0633_ (
    .A(_0147_),
    .B(_0280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0306_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0634_ (
    .A1_N(io_out[9]),
    .A2_N(_0306_),
    .B1(io_out[9]),
    .B2(_0306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0307_)
  );
  sky130_fd_sc_hd__nor2_4 _0635_ (
    .A(wbs_dat_i[9]),
    .B(_0276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0308_)
  );
  sky130_fd_sc_hd__a211o_4 _0636_ (
    .A1(_0286_),
    .A2(_0307_),
    .B1(_0262_),
    .C1(_0308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0309_)
  );
  sky130_fd_sc_hd__inv_2 _0637_ (
    .A(_0309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0074_)
  );
  sky130_fd_sc_hd__or2_4 _0638_ (
    .A(wbs_dat_i[8]),
    .B(_0278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0310_)
  );
  sky130_fd_sc_hd__and2_4 _0639_ (
    .A(_0147_),
    .B(_0280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0311_)
  );
  sky130_fd_sc_hd__o21ai_4 _0640_ (
    .A1(_0306_),
    .A2(_0311_),
    .B1(_0286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0312_)
  );
  sky130_fd_sc_hd__and3_4 _0641_ (
    .A(_0253_),
    .B(_0310_),
    .C(_0312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0073_)
  );
  sky130_fd_sc_hd__buf_2 _0642_ (
    .A(_0100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0313_)
  );
  sky130_fd_sc_hd__inv_2 _0643_ (
    .A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0314_)
  );
  sky130_fd_sc_hd__or4_4 _0644_ (
    .A(wbs_ack_o),
    .B(_0106_),
    .C(_0107_),
    .D(_0314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0315_)
  );
  sky130_fd_sc_hd__buf_2 _0645_ (
    .A(_0315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0316_)
  );
  sky130_fd_sc_hd__or2_4 _0646_ (
    .A(wbs_dat_i[7]),
    .B(_0316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0317_)
  );
  sky130_fd_sc_hd__or2_4 _0647_ (
    .A(_0257_),
    .B(_0139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0318_)
  );
  sky130_fd_sc_hd__or2_4 _0648_ (
    .A(_0131_),
    .B(_0318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0319_)
  );
  sky130_fd_sc_hd__or2_4 _0649_ (
    .A(_0130_),
    .B(_0319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0320_)
  );
  sky130_fd_sc_hd__or2_4 _0650_ (
    .A(_0133_),
    .B(_0320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0321_)
  );
  sky130_fd_sc_hd__inv_2 _0651_ (
    .A(_0315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0322_)
  );
  sky130_fd_sc_hd__nor2_4 _0652_ (
    .A(io_out[7]),
    .B(_0321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0323_)
  );
  sky130_fd_sc_hd__a211o_4 _0653_ (
    .A1(io_out[7]),
    .A2(_0321_),
    .B1(_0322_),
    .C1(_0323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0324_)
  );
  sky130_fd_sc_hd__and3_4 _0654_ (
    .A(_0313_),
    .B(_0317_),
    .C(_0324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0072_)
  );
  sky130_fd_sc_hd__or2_4 _0655_ (
    .A(wbs_dat_i[6]),
    .B(_0316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0325_)
  );
  sky130_fd_sc_hd__nand2_4 _0656_ (
    .A(_0133_),
    .B(_0320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0326_)
  );
  sky130_fd_sc_hd__a21o_4 _0657_ (
    .A1(_0321_),
    .A2(_0326_),
    .B1(_0322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0327_)
  );
  sky130_fd_sc_hd__and3_4 _0658_ (
    .A(_0313_),
    .B(_0325_),
    .C(_0327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0071_)
  );
  sky130_fd_sc_hd__or2_4 _0659_ (
    .A(wbs_dat_i[5]),
    .B(_0316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0328_)
  );
  sky130_fd_sc_hd__nand2_4 _0660_ (
    .A(_0130_),
    .B(_0319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0329_)
  );
  sky130_fd_sc_hd__a21o_4 _0661_ (
    .A1(_0320_),
    .A2(_0329_),
    .B1(_0322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0330_)
  );
  sky130_fd_sc_hd__and3_4 _0662_ (
    .A(_0313_),
    .B(_0328_),
    .C(_0330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0070_)
  );
  sky130_fd_sc_hd__or2_4 _0663_ (
    .A(wbs_dat_i[4]),
    .B(_0316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0331_)
  );
  sky130_fd_sc_hd__nand2_4 _0664_ (
    .A(_0131_),
    .B(_0318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0332_)
  );
  sky130_fd_sc_hd__a21o_4 _0665_ (
    .A1(_0319_),
    .A2(_0332_),
    .B1(_0322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0333_)
  );
  sky130_fd_sc_hd__and3_4 _0666_ (
    .A(_0313_),
    .B(_0331_),
    .C(_0333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0069_)
  );
  sky130_fd_sc_hd__or2_4 _0667_ (
    .A(_0138_),
    .B(_0257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0334_)
  );
  sky130_fd_sc_hd__or2_4 _0668_ (
    .A(_0137_),
    .B(_0334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0335_)
  );
  sky130_fd_sc_hd__inv_2 _0669_ (
    .A(_0335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0336_)
  );
  sky130_fd_sc_hd__a21o_4 _0670_ (
    .A1(io_out[2]),
    .A2(_0336_),
    .B1(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0337_)
  );
  sky130_fd_sc_hd__a32o_4 _0671_ (
    .A1(_0318_),
    .A2(_0315_),
    .A3(_0337_),
    .B1(wbs_dat_i[3]),
    .B2(_0322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0338_)
  );
  sky130_fd_sc_hd__and2_4 _0672_ (
    .A(_0223_),
    .B(_0338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0068_)
  );
  sky130_fd_sc_hd__buf_2 _0673_ (
    .A(_0315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0339_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0674_ (
    .A1_N(_0136_),
    .A2_N(_0335_),
    .B1(_0136_),
    .B2(_0335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0340_)
  );
  sky130_fd_sc_hd__nor2_4 _0675_ (
    .A(wbs_dat_i[2]),
    .B(_0339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0341_)
  );
  sky130_fd_sc_hd__a211o_4 _0676_ (
    .A1(_0339_),
    .A2(_0340_),
    .B1(_0099_),
    .C1(_0341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0342_)
  );
  sky130_fd_sc_hd__inv_2 _0677_ (
    .A(_0342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0067_)
  );
  sky130_fd_sc_hd__or2_4 _0678_ (
    .A(wbs_dat_i[1]),
    .B(_0316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0343_)
  );
  sky130_fd_sc_hd__and2_4 _0679_ (
    .A(_0137_),
    .B(_0334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0344_)
  );
  sky130_fd_sc_hd__o21ai_4 _0680_ (
    .A1(_0336_),
    .A2(_0344_),
    .B1(_0339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0345_)
  );
  sky130_fd_sc_hd__and3_4 _0681_ (
    .A(_0313_),
    .B(_0343_),
    .C(_0345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0066_)
  );
  sky130_fd_sc_hd__a21bo_4 _0682_ (
    .A1(_0138_),
    .A2(_0257_),
    .B1_N(_0334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0346_)
  );
  sky130_fd_sc_hd__nor2_4 _0683_ (
    .A(wbs_dat_i[0]),
    .B(_0339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0347_)
  );
  sky130_fd_sc_hd__a211o_4 _0684_ (
    .A1(_0339_),
    .A2(_0346_),
    .B1(_0099_),
    .C1(_0347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0348_)
  );
  sky130_fd_sc_hd__inv_2 _0685_ (
    .A(_0348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0065_)
  );
  sky130_fd_sc_hd__or3_4 _0686_ (
    .A(wbs_ack_o),
    .B(_0106_),
    .C(_0098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0349_)
  );
  sky130_fd_sc_hd__inv_2 _0687_ (
    .A(_0349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0350_)
  );
  sky130_fd_sc_hd__buf_2 _0688_ (
    .A(_0350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0064_)
  );
  sky130_fd_sc_hd__inv_2 _0689_ (
    .A(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0351_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0690_ (
    .A1_N(_0351_),
    .A2_N(_0196_),
    .B1(la_data_in[63]),
    .B2(_0196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0063_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0691_ (
    .A1_N(_0112_),
    .A2_N(_0195_),
    .B1(la_data_in[62]),
    .B2(_0195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0062_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0692_ (
    .A1_N(_0113_),
    .A2_N(_0197_),
    .B1(la_data_in[61]),
    .B2(_0197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0061_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0693_ (
    .A1_N(_0114_),
    .A2_N(_0194_),
    .B1(la_data_in[60]),
    .B2(_0194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0060_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0694_ (
    .A1_N(_0117_),
    .A2_N(_0191_),
    .B1(la_data_in[59]),
    .B2(_0191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0059_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0695_ (
    .A1_N(_0118_),
    .A2_N(_0190_),
    .B1(la_data_in[58]),
    .B2(_0190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0058_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0696_ (
    .A1_N(_0115_),
    .A2_N(_0192_),
    .B1(la_data_in[57]),
    .B2(_0192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0057_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0697_ (
    .A1_N(_0116_),
    .A2_N(_0189_),
    .B1(la_data_in[56]),
    .B2(_0189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0056_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0698_ (
    .A1_N(_0127_),
    .A2_N(_0186_),
    .B1(la_data_in[55]),
    .B2(_0186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0055_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0699_ (
    .A1_N(_0128_),
    .A2_N(_0185_),
    .B1(la_data_in[54]),
    .B2(_0185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0054_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0700_ (
    .A1_N(_0125_),
    .A2_N(_0187_),
    .B1(la_data_in[53]),
    .B2(_0187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0053_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0701_ (
    .A1_N(_0126_),
    .A2_N(_0184_),
    .B1(la_data_in[52]),
    .B2(_0184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0052_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0702_ (
    .A1_N(_0122_),
    .A2_N(_0181_),
    .B1(la_data_in[51]),
    .B2(_0181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0051_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0703_ (
    .A1_N(_0123_),
    .A2_N(_0180_),
    .B1(la_data_in[50]),
    .B2(_0180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0050_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0704_ (
    .A1_N(_0120_),
    .A2_N(_0182_),
    .B1(la_data_in[49]),
    .B2(_0182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0049_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0705_ (
    .A1_N(_0121_),
    .A2_N(_0179_),
    .B1(la_data_in[48]),
    .B2(_0179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0048_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0706_ (
    .A1_N(_0145_),
    .A2_N(_0175_),
    .B1(la_data_in[47]),
    .B2(_0175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0047_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0707_ (
    .A1_N(_0142_),
    .A2_N(_0174_),
    .B1(la_data_in[46]),
    .B2(_0174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0046_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0708_ (
    .A1_N(_0143_),
    .A2_N(_0176_),
    .B1(la_data_in[45]),
    .B2(_0176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0045_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0709_ (
    .A1_N(_0141_),
    .A2_N(_0173_),
    .B1(la_data_in[44]),
    .B2(_0173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0044_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0710_ (
    .A1_N(_0148_),
    .A2_N(_0169_),
    .B1(la_data_in[43]),
    .B2(_0169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0043_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0711_ (
    .A1_N(_0149_),
    .A2_N(_0167_),
    .B1(la_data_in[42]),
    .B2(_0167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0042_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0712_ (
    .A1_N(_0146_),
    .A2_N(_0171_),
    .B1(la_data_in[41]),
    .B2(_0171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0041_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0713_ (
    .A1_N(_0147_),
    .A2_N(_0166_),
    .B1(la_data_in[40]),
    .B2(_0166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0040_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0714_ (
    .A1_N(_0132_),
    .A2_N(_0163_),
    .B1(la_data_in[39]),
    .B2(_0163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0039_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0715_ (
    .A1_N(_0133_),
    .A2_N(_0161_),
    .B1(la_data_in[38]),
    .B2(_0161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0038_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0716_ (
    .A1_N(_0130_),
    .A2_N(_0164_),
    .B1(la_data_in[37]),
    .B2(_0164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0037_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0717_ (
    .A1_N(_0131_),
    .A2_N(_0160_),
    .B1(la_data_in[36]),
    .B2(_0160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0036_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0718_ (
    .A1_N(_0135_),
    .A2_N(_0156_),
    .B1(la_data_in[35]),
    .B2(_0156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0035_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0719_ (
    .A1_N(_0136_),
    .A2_N(_0154_),
    .B1(la_data_in[34]),
    .B2(_0154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0034_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0720_ (
    .A1_N(_0137_),
    .A2_N(_0158_),
    .B1(la_data_in[33]),
    .B2(_0158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0033_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0721_ (
    .A1_N(_0138_),
    .A2_N(_0153_),
    .B1(la_data_in[32]),
    .B2(_0153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0032_)
  );
  sky130_fd_sc_hd__inv_2 _0722_ (
    .A(wbs_dat_o[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0352_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0723_ (
    .A1_N(_0352_),
    .A2_N(_0064_),
    .B1(io_out[31]),
    .B2(_0064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0031_)
  );
  sky130_fd_sc_hd__inv_2 _0724_ (
    .A(wbs_dat_o[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0353_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0725_ (
    .A1_N(_0353_),
    .A2_N(_0064_),
    .B1(io_out[30]),
    .B2(_0064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0030_)
  );
  sky130_fd_sc_hd__inv_2 _0726_ (
    .A(wbs_dat_o[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0354_)
  );
  sky130_fd_sc_hd__buf_2 _0727_ (
    .A(_0350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0355_)
  );
  sky130_fd_sc_hd__buf_2 _0728_ (
    .A(_0355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0356_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0729_ (
    .A1_N(_0354_),
    .A2_N(_0356_),
    .B1(io_out[29]),
    .B2(_0356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0029_)
  );
  sky130_fd_sc_hd__inv_2 _0730_ (
    .A(wbs_dat_o[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0357_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0731_ (
    .A1_N(_0357_),
    .A2_N(_0356_),
    .B1(io_out[28]),
    .B2(_0356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0028_)
  );
  sky130_fd_sc_hd__inv_2 _0732_ (
    .A(wbs_dat_o[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0358_)
  );
  sky130_fd_sc_hd__buf_2 _0733_ (
    .A(_0350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0359_)
  );
  sky130_fd_sc_hd__buf_2 _0734_ (
    .A(_0359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0360_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0735_ (
    .A1_N(_0358_),
    .A2_N(_0356_),
    .B1(io_out[27]),
    .B2(_0360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0027_)
  );
  sky130_fd_sc_hd__inv_2 _0736_ (
    .A(wbs_dat_o[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0361_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0737_ (
    .A1_N(_0361_),
    .A2_N(_0360_),
    .B1(io_out[26]),
    .B2(_0360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0026_)
  );
  sky130_fd_sc_hd__inv_2 _0738_ (
    .A(wbs_dat_o[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0362_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0739_ (
    .A1_N(_0362_),
    .A2_N(_0360_),
    .B1(io_out[25]),
    .B2(_0360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0025_)
  );
  sky130_fd_sc_hd__inv_2 _0740_ (
    .A(wbs_dat_o[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0363_)
  );
  sky130_fd_sc_hd__buf_2 _0741_ (
    .A(_0355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0364_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0742_ (
    .A1_N(_0363_),
    .A2_N(_0364_),
    .B1(io_out[24]),
    .B2(_0364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0024_)
  );
  sky130_fd_sc_hd__inv_2 _0743_ (
    .A(wbs_dat_o[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0365_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0744_ (
    .A1_N(_0365_),
    .A2_N(_0364_),
    .B1(io_out[23]),
    .B2(_0364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0023_)
  );
  sky130_fd_sc_hd__inv_2 _0745_ (
    .A(wbs_dat_o[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0366_)
  );
  sky130_fd_sc_hd__buf_2 _0746_ (
    .A(_0359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0367_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0747_ (
    .A1_N(_0366_),
    .A2_N(_0364_),
    .B1(io_out[22]),
    .B2(_0367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0022_)
  );
  sky130_fd_sc_hd__inv_2 _0748_ (
    .A(wbs_dat_o[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0368_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0749_ (
    .A1_N(_0368_),
    .A2_N(_0367_),
    .B1(io_out[21]),
    .B2(_0367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0021_)
  );
  sky130_fd_sc_hd__inv_2 _0750_ (
    .A(wbs_dat_o[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0369_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0751_ (
    .A1_N(_0369_),
    .A2_N(_0367_),
    .B1(io_out[20]),
    .B2(_0367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0020_)
  );
  sky130_fd_sc_hd__inv_2 _0752_ (
    .A(wbs_dat_o[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0370_)
  );
  sky130_fd_sc_hd__buf_2 _0753_ (
    .A(_0355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0371_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0754_ (
    .A1_N(_0370_),
    .A2_N(_0371_),
    .B1(io_out[19]),
    .B2(_0371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0019_)
  );
  sky130_fd_sc_hd__inv_2 _0755_ (
    .A(wbs_dat_o[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0372_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0756_ (
    .A1_N(_0372_),
    .A2_N(_0371_),
    .B1(io_out[18]),
    .B2(_0371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0018_)
  );
  sky130_fd_sc_hd__inv_2 _0757_ (
    .A(wbs_dat_o[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0373_)
  );
  sky130_fd_sc_hd__buf_2 _0758_ (
    .A(_0359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0374_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0759_ (
    .A1_N(_0373_),
    .A2_N(_0371_),
    .B1(io_out[17]),
    .B2(_0374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0017_)
  );
  sky130_fd_sc_hd__inv_2 _0760_ (
    .A(wbs_dat_o[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0375_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0761_ (
    .A1_N(_0375_),
    .A2_N(_0374_),
    .B1(io_out[16]),
    .B2(_0374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0016_)
  );
  sky130_fd_sc_hd__inv_2 _0762_ (
    .A(wbs_dat_o[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0376_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0763_ (
    .A1_N(_0376_),
    .A2_N(_0374_),
    .B1(io_out[15]),
    .B2(_0374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0015_)
  );
  sky130_fd_sc_hd__inv_2 _0764_ (
    .A(wbs_dat_o[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0377_)
  );
  sky130_fd_sc_hd__buf_2 _0765_ (
    .A(_0355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0378_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0766_ (
    .A1_N(_0377_),
    .A2_N(_0378_),
    .B1(io_out[14]),
    .B2(_0378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0014_)
  );
  sky130_fd_sc_hd__inv_2 _0767_ (
    .A(wbs_dat_o[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0379_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0768_ (
    .A1_N(_0379_),
    .A2_N(_0378_),
    .B1(io_out[13]),
    .B2(_0378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0013_)
  );
  sky130_fd_sc_hd__inv_2 _0769_ (
    .A(wbs_dat_o[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0380_)
  );
  sky130_fd_sc_hd__buf_2 _0770_ (
    .A(_0359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0381_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0771_ (
    .A1_N(_0380_),
    .A2_N(_0378_),
    .B1(io_out[12]),
    .B2(_0381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0012_)
  );
  sky130_fd_sc_hd__inv_2 _0772_ (
    .A(wbs_dat_o[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0382_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0773_ (
    .A1_N(_0382_),
    .A2_N(_0381_),
    .B1(io_out[11]),
    .B2(_0381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0011_)
  );
  sky130_fd_sc_hd__inv_2 _0774_ (
    .A(wbs_dat_o[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0383_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0775_ (
    .A1_N(_0383_),
    .A2_N(_0381_),
    .B1(io_out[10]),
    .B2(_0381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0010_)
  );
  sky130_fd_sc_hd__inv_2 _0776_ (
    .A(wbs_dat_o[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0384_)
  );
  sky130_fd_sc_hd__buf_2 _0777_ (
    .A(_0355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0385_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0778_ (
    .A1_N(_0384_),
    .A2_N(_0385_),
    .B1(io_out[9]),
    .B2(_0385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0009_)
  );
  sky130_fd_sc_hd__inv_2 _0779_ (
    .A(wbs_dat_o[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0386_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0780_ (
    .A1_N(_0386_),
    .A2_N(_0385_),
    .B1(io_out[8]),
    .B2(_0385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0008_)
  );
  sky130_fd_sc_hd__inv_2 _0781_ (
    .A(wbs_dat_o[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0387_)
  );
  sky130_fd_sc_hd__buf_2 _0782_ (
    .A(_0350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0388_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0783_ (
    .A1_N(_0387_),
    .A2_N(_0385_),
    .B1(io_out[7]),
    .B2(_0388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0007_)
  );
  sky130_fd_sc_hd__inv_2 _0784_ (
    .A(wbs_dat_o[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0389_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0785_ (
    .A1_N(_0389_),
    .A2_N(_0388_),
    .B1(io_out[6]),
    .B2(_0388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0006_)
  );
  sky130_fd_sc_hd__inv_2 _0786_ (
    .A(wbs_dat_o[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0390_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0787_ (
    .A1_N(_0390_),
    .A2_N(_0388_),
    .B1(io_out[5]),
    .B2(_0388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0005_)
  );
  sky130_fd_sc_hd__inv_2 _0788_ (
    .A(wbs_dat_o[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0391_)
  );
  sky130_fd_sc_hd__buf_2 _0789_ (
    .A(_0359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0392_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0790_ (
    .A1_N(_0391_),
    .A2_N(_0392_),
    .B1(io_out[4]),
    .B2(_0392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0004_)
  );
  sky130_fd_sc_hd__inv_2 _0791_ (
    .A(wbs_dat_o[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0393_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0792_ (
    .A1_N(_0393_),
    .A2_N(_0392_),
    .B1(io_out[3]),
    .B2(_0392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0003_)
  );
  sky130_fd_sc_hd__inv_2 _0793_ (
    .A(wbs_dat_o[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0394_)
  );
  sky130_fd_sc_hd__buf_2 _0794_ (
    .A(_0350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0395_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0795_ (
    .A1_N(_0394_),
    .A2_N(_0392_),
    .B1(io_out[2]),
    .B2(_0395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0002_)
  );
  sky130_fd_sc_hd__inv_2 _0796_ (
    .A(wbs_dat_o[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0396_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0797_ (
    .A1_N(_0396_),
    .A2_N(_0395_),
    .B1(io_out[1]),
    .B2(_0395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0001_)
  );
  sky130_fd_sc_hd__inv_2 _0798_ (
    .A(wbs_dat_o[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0397_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _0799_ (
    .A1_N(_0397_),
    .A2_N(_0395_),
    .B1(io_out[0]),
    .B2(_0395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0000_)
  );
  sky130_fd_sc_hd__inv_2 _0800_ (
    .A(la_oen[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0398_)
  );
  sky130_fd_sc_hd__o22a_4 _0801_ (
    .A1(la_data_in[64]),
    .A2(la_oen[64]),
    .B1(wb_clk_i),
    .B2(_0398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\counter.clk )
  );
  sky130_fd_sc_hd__or2_4 _0802_ (
    .A(wbs_dat_i[31]),
    .B(_0206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0399_)
  );
  sky130_fd_sc_hd__nor2_4 _0803_ (
    .A(io_out[31]),
    .B(_0205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_0400_)
  );
  sky130_fd_sc_hd__a211o_4 _0804_ (
    .A1(io_out[31]),
    .A2(_0205_),
    .B1(_0207_),
    .C1(_0400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0401_)
  );
  sky130_fd_sc_hd__and3_4 _0805_ (
    .A(_0100_),
    .B(_0399_),
    .C(_0401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_0096_)
  );
  sky130_fd_sc_hd__conb_1 _0806_ (
    .LO(io_oeb[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0807_ (
    .LO(io_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0808_ (
    .LO(io_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0809_ (
    .LO(io_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0810_ (
    .LO(io_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0811_ (
    .LO(io_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0812_ (
    .LO(io_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0813_ (
    .LO(la_data_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0814_ (
    .LO(la_data_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0815_ (
    .LO(la_data_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0816_ (
    .LO(la_data_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0817_ (
    .LO(la_data_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0818_ (
    .LO(la_data_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0819_ (
    .LO(la_data_out[38]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0820_ (
    .LO(la_data_out[39]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0821_ (
    .LO(la_data_out[40]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0822_ (
    .LO(la_data_out[41]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0823_ (
    .LO(la_data_out[42]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0824_ (
    .LO(la_data_out[43]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0825_ (
    .LO(la_data_out[44]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0826_ (
    .LO(la_data_out[45]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0827_ (
    .LO(la_data_out[46]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0828_ (
    .LO(la_data_out[47]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0829_ (
    .LO(la_data_out[48]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0830_ (
    .LO(la_data_out[49]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0831_ (
    .LO(la_data_out[50]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0832_ (
    .LO(la_data_out[51]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0833_ (
    .LO(la_data_out[52]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0834_ (
    .LO(la_data_out[53]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0835_ (
    .LO(la_data_out[54]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0836_ (
    .LO(la_data_out[55]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0837_ (
    .LO(la_data_out[56]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0838_ (
    .LO(la_data_out[57]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0839_ (
    .LO(la_data_out[58]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0840_ (
    .LO(la_data_out[59]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0841_ (
    .LO(la_data_out[60]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0842_ (
    .LO(la_data_out[61]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0843_ (
    .LO(la_data_out[62]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0844_ (
    .LO(la_data_out[63]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0845_ (
    .LO(la_data_out[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0846_ (
    .LO(la_data_out[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0847_ (
    .LO(la_data_out[66]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0848_ (
    .LO(la_data_out[67]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0849_ (
    .LO(la_data_out[68]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0850_ (
    .LO(la_data_out[69]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0851_ (
    .LO(la_data_out[70]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0852_ (
    .LO(la_data_out[71]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0853_ (
    .LO(la_data_out[72]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0854_ (
    .LO(la_data_out[73]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0855_ (
    .LO(la_data_out[74]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0856_ (
    .LO(la_data_out[75]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0857_ (
    .LO(la_data_out[76]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0858_ (
    .LO(la_data_out[77]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0859_ (
    .LO(la_data_out[78]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0860_ (
    .LO(la_data_out[79]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0861_ (
    .LO(la_data_out[80]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0862_ (
    .LO(la_data_out[81]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0863_ (
    .LO(la_data_out[82]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0864_ (
    .LO(la_data_out[83]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0865_ (
    .LO(la_data_out[84]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0866_ (
    .LO(la_data_out[85]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0867_ (
    .LO(la_data_out[86]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0868_ (
    .LO(la_data_out[87]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0869_ (
    .LO(la_data_out[88]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0870_ (
    .LO(la_data_out[89]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0871_ (
    .LO(la_data_out[90]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0872_ (
    .LO(la_data_out[91]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0873_ (
    .LO(la_data_out[92]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0874_ (
    .LO(la_data_out[93]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0875_ (
    .LO(la_data_out[94]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0876_ (
    .LO(la_data_out[95]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0877_ (
    .LO(la_data_out[96]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0878_ (
    .LO(la_data_out[97]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0879_ (
    .LO(la_data_out[98]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0880_ (
    .LO(la_data_out[99]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0881_ (
    .LO(la_data_out[100]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0882_ (
    .LO(la_data_out[101]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0883_ (
    .LO(la_data_out[102]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0884_ (
    .LO(la_data_out[103]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0885_ (
    .LO(la_data_out[104]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0886_ (
    .LO(la_data_out[105]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0887_ (
    .LO(la_data_out[106]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0888_ (
    .LO(la_data_out[107]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0889_ (
    .LO(la_data_out[108]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0890_ (
    .LO(la_data_out[109]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0891_ (
    .LO(la_data_out[110]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0892_ (
    .LO(la_data_out[111]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0893_ (
    .LO(la_data_out[112]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0894_ (
    .LO(la_data_out[113]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0895_ (
    .LO(la_data_out[114]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0896_ (
    .LO(la_data_out[115]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0897_ (
    .LO(la_data_out[116]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0898_ (
    .LO(la_data_out[117]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0899_ (
    .LO(la_data_out[118]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0900_ (
    .LO(la_data_out[119]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0901_ (
    .LO(la_data_out[120]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0902_ (
    .LO(la_data_out[121]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0903_ (
    .LO(la_data_out[122]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0904_ (
    .LO(la_data_out[123]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0905_ (
    .LO(la_data_out[124]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0906_ (
    .LO(la_data_out[125]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0907_ (
    .LO(la_data_out[126]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 _0908_ (
    .LO(la_data_out[127]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__buf_2 _0909_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[0])
  );
  sky130_fd_sc_hd__buf_2 _0910_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[1])
  );
  sky130_fd_sc_hd__buf_2 _0911_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[2])
  );
  sky130_fd_sc_hd__buf_2 _0912_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[3])
  );
  sky130_fd_sc_hd__buf_2 _0913_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[4])
  );
  sky130_fd_sc_hd__buf_2 _0914_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[5])
  );
  sky130_fd_sc_hd__buf_2 _0915_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[6])
  );
  sky130_fd_sc_hd__buf_2 _0916_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[7])
  );
  sky130_fd_sc_hd__buf_2 _0917_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[8])
  );
  sky130_fd_sc_hd__buf_2 _0918_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[9])
  );
  sky130_fd_sc_hd__buf_2 _0919_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[10])
  );
  sky130_fd_sc_hd__buf_2 _0920_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[11])
  );
  sky130_fd_sc_hd__buf_2 _0921_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[12])
  );
  sky130_fd_sc_hd__buf_2 _0922_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[13])
  );
  sky130_fd_sc_hd__buf_2 _0923_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[14])
  );
  sky130_fd_sc_hd__buf_2 _0924_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[15])
  );
  sky130_fd_sc_hd__buf_2 _0925_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[16])
  );
  sky130_fd_sc_hd__buf_2 _0926_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[17])
  );
  sky130_fd_sc_hd__buf_2 _0927_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[18])
  );
  sky130_fd_sc_hd__buf_2 _0928_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[19])
  );
  sky130_fd_sc_hd__buf_2 _0929_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[20])
  );
  sky130_fd_sc_hd__buf_2 _0930_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[21])
  );
  sky130_fd_sc_hd__buf_2 _0931_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[22])
  );
  sky130_fd_sc_hd__buf_2 _0932_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[23])
  );
  sky130_fd_sc_hd__buf_2 _0933_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[24])
  );
  sky130_fd_sc_hd__buf_2 _0934_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[25])
  );
  sky130_fd_sc_hd__buf_2 _0935_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[26])
  );
  sky130_fd_sc_hd__buf_2 _0936_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[27])
  );
  sky130_fd_sc_hd__buf_2 _0937_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[28])
  );
  sky130_fd_sc_hd__buf_2 _0938_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[29])
  );
  sky130_fd_sc_hd__buf_2 _0939_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[30])
  );
  sky130_fd_sc_hd__buf_2 _0940_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[31])
  );
  sky130_fd_sc_hd__buf_2 _0941_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[32])
  );
  sky130_fd_sc_hd__buf_2 _0942_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[33])
  );
  sky130_fd_sc_hd__buf_2 _0943_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[34])
  );
  sky130_fd_sc_hd__buf_2 _0944_ (
    .A(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[35])
  );
  sky130_fd_sc_hd__buf_2 _0945_ (
    .A(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[0])
  );
  sky130_fd_sc_hd__buf_2 _0946_ (
    .A(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[1])
  );
  sky130_fd_sc_hd__buf_2 _0947_ (
    .A(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[2])
  );
  sky130_fd_sc_hd__buf_2 _0948_ (
    .A(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[3])
  );
  sky130_fd_sc_hd__buf_2 _0949_ (
    .A(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[4])
  );
  sky130_fd_sc_hd__buf_2 _0950_ (
    .A(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[5])
  );
  sky130_fd_sc_hd__buf_2 _0951_ (
    .A(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[6])
  );
  sky130_fd_sc_hd__buf_2 _0952_ (
    .A(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[7])
  );
  sky130_fd_sc_hd__buf_2 _0953_ (
    .A(io_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[8])
  );
  sky130_fd_sc_hd__buf_2 _0954_ (
    .A(io_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[9])
  );
  sky130_fd_sc_hd__buf_2 _0955_ (
    .A(io_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[10])
  );
  sky130_fd_sc_hd__buf_2 _0956_ (
    .A(io_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[11])
  );
  sky130_fd_sc_hd__buf_2 _0957_ (
    .A(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[12])
  );
  sky130_fd_sc_hd__buf_2 _0958_ (
    .A(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[13])
  );
  sky130_fd_sc_hd__buf_2 _0959_ (
    .A(io_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[14])
  );
  sky130_fd_sc_hd__buf_2 _0960_ (
    .A(io_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[15])
  );
  sky130_fd_sc_hd__buf_2 _0961_ (
    .A(io_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[16])
  );
  sky130_fd_sc_hd__buf_2 _0962_ (
    .A(io_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[17])
  );
  sky130_fd_sc_hd__buf_2 _0963_ (
    .A(io_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[18])
  );
  sky130_fd_sc_hd__buf_2 _0964_ (
    .A(io_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[19])
  );
  sky130_fd_sc_hd__buf_2 _0965_ (
    .A(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[20])
  );
  sky130_fd_sc_hd__buf_2 _0966_ (
    .A(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[21])
  );
  sky130_fd_sc_hd__buf_2 _0967_ (
    .A(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[22])
  );
  sky130_fd_sc_hd__buf_2 _0968_ (
    .A(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[23])
  );
  sky130_fd_sc_hd__buf_2 _0969_ (
    .A(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[24])
  );
  sky130_fd_sc_hd__buf_2 _0970_ (
    .A(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[25])
  );
  sky130_fd_sc_hd__buf_2 _0971_ (
    .A(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[26])
  );
  sky130_fd_sc_hd__buf_2 _0972_ (
    .A(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[27])
  );
  sky130_fd_sc_hd__buf_2 _0973_ (
    .A(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[28])
  );
  sky130_fd_sc_hd__buf_2 _0974_ (
    .A(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[29])
  );
  sky130_fd_sc_hd__buf_2 _0975_ (
    .A(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[30])
  );
  sky130_fd_sc_hd__buf_2 _0976_ (
    .A(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[31])
  );
  sky130_fd_sc_hd__dfxtp_4 _0977_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0000_),
    .Q(wbs_dat_o[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0978_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0001_),
    .Q(wbs_dat_o[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0979_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0002_),
    .Q(wbs_dat_o[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0980_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0003_),
    .Q(wbs_dat_o[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0981_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0004_),
    .Q(wbs_dat_o[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0982_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0005_),
    .Q(wbs_dat_o[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0983_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0006_),
    .Q(wbs_dat_o[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0984_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0007_),
    .Q(wbs_dat_o[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0985_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0008_),
    .Q(wbs_dat_o[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0986_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0009_),
    .Q(wbs_dat_o[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0987_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0010_),
    .Q(wbs_dat_o[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0988_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0011_),
    .Q(wbs_dat_o[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0989_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0012_),
    .Q(wbs_dat_o[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0990_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0013_),
    .Q(wbs_dat_o[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0991_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0014_),
    .Q(wbs_dat_o[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0992_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0015_),
    .Q(wbs_dat_o[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0993_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0016_),
    .Q(wbs_dat_o[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0994_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0017_),
    .Q(wbs_dat_o[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0995_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0018_),
    .Q(wbs_dat_o[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0996_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0019_),
    .Q(wbs_dat_o[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0997_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0020_),
    .Q(wbs_dat_o[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0998_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0021_),
    .Q(wbs_dat_o[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _0999_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0022_),
    .Q(wbs_dat_o[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1000_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0023_),
    .Q(wbs_dat_o[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1001_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0024_),
    .Q(wbs_dat_o[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1002_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0025_),
    .Q(wbs_dat_o[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1003_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0026_),
    .Q(wbs_dat_o[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1004_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0027_),
    .Q(wbs_dat_o[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1005_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0028_),
    .Q(wbs_dat_o[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1006_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0029_),
    .Q(wbs_dat_o[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1007_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0030_),
    .Q(wbs_dat_o[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1008_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0031_),
    .Q(wbs_dat_o[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1009_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0032_),
    .Q(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1010_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0033_),
    .Q(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1011_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0034_),
    .Q(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1012_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0035_),
    .Q(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1013_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0036_),
    .Q(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1014_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0037_),
    .Q(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1015_ (
    .CLK(\clknet_3_1_0_counter.clk ),
    .D(_0038_),
    .Q(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1016_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0039_),
    .Q(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1017_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0040_),
    .Q(io_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1018_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0041_),
    .Q(io_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1019_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0042_),
    .Q(io_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1020_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0043_),
    .Q(io_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1021_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0044_),
    .Q(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1022_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0045_),
    .Q(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1023_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0046_),
    .Q(io_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1024_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0047_),
    .Q(io_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1025_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0048_),
    .Q(io_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1026_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0049_),
    .Q(io_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1027_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0050_),
    .Q(io_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1028_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0051_),
    .Q(io_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1029_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0052_),
    .Q(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1030_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0053_),
    .Q(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1031_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0054_),
    .Q(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1032_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0055_),
    .Q(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1033_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0056_),
    .Q(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1034_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0057_),
    .Q(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1035_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0058_),
    .Q(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1036_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0059_),
    .Q(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1037_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0060_),
    .Q(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1038_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0061_),
    .Q(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1039_ (
    .CLK(\clknet_3_5_0_counter.clk ),
    .D(_0062_),
    .Q(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1040_ (
    .CLK(\clknet_3_4_0_counter.clk ),
    .D(_0063_),
    .Q(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1041_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0064_),
    .Q(wbs_ack_o),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1042_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0065_),
    .Q(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1043_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0066_),
    .Q(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1044_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0067_),
    .Q(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1045_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0068_),
    .Q(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1046_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0069_),
    .Q(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1047_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0070_),
    .Q(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1048_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0071_),
    .Q(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1049_ (
    .CLK(\clknet_3_0_0_counter.clk ),
    .D(_0072_),
    .Q(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1050_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0073_),
    .Q(io_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1051_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0074_),
    .Q(io_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1052_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0075_),
    .Q(io_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1053_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0076_),
    .Q(io_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1054_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0077_),
    .Q(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1055_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0078_),
    .Q(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1056_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0079_),
    .Q(io_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1057_ (
    .CLK(\clknet_3_2_0_counter.clk ),
    .D(_0080_),
    .Q(io_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1058_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0081_),
    .Q(io_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1059_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0082_),
    .Q(io_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1060_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0083_),
    .Q(io_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1061_ (
    .CLK(\clknet_3_3_0_counter.clk ),
    .D(_0084_),
    .Q(io_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1062_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0085_),
    .Q(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1063_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0086_),
    .Q(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1064_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0087_),
    .Q(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1065_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0088_),
    .Q(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1066_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0089_),
    .Q(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1067_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0090_),
    .Q(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1068_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0091_),
    .Q(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1069_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0092_),
    .Q(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1070_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0093_),
    .Q(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1071_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0094_),
    .Q(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1072_ (
    .CLK(\clknet_3_7_0_counter.clk ),
    .D(_0095_),
    .Q(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _1073_ (
    .CLK(\clknet_3_6_0_counter.clk ),
    .D(_0096_),
    .Q(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_counter.clk  (
    .A(\counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_1_0_0_counter.clk  (
    .A(\clknet_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_1_1_0_counter.clk  (
    .A(\clknet_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_0_0_counter.clk  (
    .A(\clknet_1_0_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_2_0_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_1_0_counter.clk  (
    .A(\clknet_1_0_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_2_1_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_2_0_counter.clk  (
    .A(\clknet_1_1_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_2_2_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_3_0_counter.clk  (
    .A(\clknet_1_1_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_2_3_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_0_0_counter.clk  (
    .A(\clknet_2_0_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_0_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_1_0_counter.clk  (
    .A(\clknet_2_0_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_1_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_2_0_counter.clk  (
    .A(\clknet_2_1_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_2_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_3_0_counter.clk  (
    .A(\clknet_2_1_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_3_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_4_0_counter.clk  (
    .A(\clknet_2_2_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_4_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_5_0_counter.clk  (
    .A(\clknet_2_2_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_5_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_6_0_counter.clk  (
    .A(\clknet_2_3_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_6_0_counter.clk )
  );
  sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_7_0_counter.clk  (
    .A(\clknet_2_3_0_counter.clk ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_3_7_0_counter.clk )
  );
endmodule
