*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* NGSPICE file created from storage.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sram_1rw1r_32_256_8_sky130 abstract view
.subckt sram_1rw1r_32_256_8_sky130 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5]
+ din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24]
+ din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0] addr0[1]
+ addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1] addr1[2]
+ addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 web0 clk0 clk1 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5]
+ dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22]
+ dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30]
+ dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7]
+ dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16]
+ dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24]
+ dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] vdd gnd
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

.subckt storage mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3] mgmt_addr[4] mgmt_addr[5]
+ mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0] mgmt_addr_ro[1] mgmt_addr_ro[2] mgmt_addr_ro[3]
+ mgmt_addr_ro[4] mgmt_addr_ro[5] mgmt_addr_ro[6] mgmt_addr_ro[7] mgmt_clk mgmt_ena[0]
+ mgmt_ena[1] mgmt_ena_ro mgmt_rdata[0] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12]
+ mgmt_rdata[13] mgmt_rdata[14] mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18]
+ mgmt_rdata[19] mgmt_rdata[1] mgmt_rdata[20] mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23]
+ mgmt_rdata[24] mgmt_rdata[25] mgmt_rdata[26] mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29]
+ mgmt_rdata[2] mgmt_rdata[30] mgmt_rdata[31] mgmt_rdata[32] mgmt_rdata[33] mgmt_rdata[34]
+ mgmt_rdata[35] mgmt_rdata[36] mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39] mgmt_rdata[3]
+ mgmt_rdata[40] mgmt_rdata[41] mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45]
+ mgmt_rdata[46] mgmt_rdata[47] mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[4] mgmt_rdata[50]
+ mgmt_rdata[51] mgmt_rdata[52] mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56]
+ mgmt_rdata[57] mgmt_rdata[58] mgmt_rdata[59] mgmt_rdata[5] mgmt_rdata[60] mgmt_rdata[61]
+ mgmt_rdata[62] mgmt_rdata[63] mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8] mgmt_rdata[9]
+ mgmt_rdata_ro[0] mgmt_rdata_ro[10] mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13]
+ mgmt_rdata_ro[14] mgmt_rdata_ro[15] mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18]
+ mgmt_rdata_ro[19] mgmt_rdata_ro[1] mgmt_rdata_ro[20] mgmt_rdata_ro[21] mgmt_rdata_ro[22]
+ mgmt_rdata_ro[23] mgmt_rdata_ro[24] mgmt_rdata_ro[25] mgmt_rdata_ro[26] mgmt_rdata_ro[27]
+ mgmt_rdata_ro[28] mgmt_rdata_ro[29] mgmt_rdata_ro[2] mgmt_rdata_ro[30] mgmt_rdata_ro[31]
+ mgmt_rdata_ro[3] mgmt_rdata_ro[4] mgmt_rdata_ro[5] mgmt_rdata_ro[6] mgmt_rdata_ro[7]
+ mgmt_rdata_ro[8] mgmt_rdata_ro[9] mgmt_wdata[0] mgmt_wdata[10] mgmt_wdata[11] mgmt_wdata[12]
+ mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17] mgmt_wdata[18]
+ mgmt_wdata[19] mgmt_wdata[1] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[2] mgmt_wdata[30] mgmt_wdata[31] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wen[0] mgmt_wen[1]
+ mgmt_wen_mask[0] mgmt_wen_mask[1] mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_wen_mask[4]
+ mgmt_wen_mask[5] mgmt_wen_mask[6] mgmt_wen_mask[7] VPWR VGND
XFILLER_338_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_329_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[23] mgmt_wdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_296_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_293_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_295_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_288_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_292_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_283_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[22] mgmt_wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_332_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_296_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_314_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_302_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_332_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_283_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_325_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[21] mgmt_wdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_265_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_331_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_287_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_318_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[20] mgmt_wdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_265_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_326_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_268_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[7] mgmt_addr_ro[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSRAM_0 mgmt_wdata[0] mgmt_wdata[1] mgmt_wdata[2] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wdata[10] mgmt_wdata[11]
+ mgmt_wdata[12] mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17]
+ mgmt_wdata[18] mgmt_wdata[19] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[30] mgmt_wdata[31] mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3]
+ mgmt_addr[4] mgmt_addr[5] mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0] mgmt_addr_ro[1]
+ mgmt_addr_ro[2] mgmt_addr_ro[3] mgmt_addr_ro[4] mgmt_addr_ro[5] mgmt_addr_ro[6]
+ mgmt_addr_ro[7] mgmt_ena[0] mgmt_ena_ro mgmt_wen[0] mgmt_clk mgmt_clk mgmt_wen_mask[0]
+ mgmt_wen_mask[1] mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_rdata[0] mgmt_rdata[1] mgmt_rdata[2]
+ mgmt_rdata[3] mgmt_rdata[4] mgmt_rdata[5] mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8]
+ mgmt_rdata[9] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12] mgmt_rdata[13] mgmt_rdata[14]
+ mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18] mgmt_rdata[19] mgmt_rdata[20]
+ mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23] mgmt_rdata[24] mgmt_rdata[25] mgmt_rdata[26]
+ mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29] mgmt_rdata[30] mgmt_rdata[31] mgmt_rdata_ro[0]
+ mgmt_rdata_ro[1] mgmt_rdata_ro[2] mgmt_rdata_ro[3] mgmt_rdata_ro[4] mgmt_rdata_ro[5]
+ mgmt_rdata_ro[6] mgmt_rdata_ro[7] mgmt_rdata_ro[8] mgmt_rdata_ro[9] mgmt_rdata_ro[10]
+ mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13] mgmt_rdata_ro[14] mgmt_rdata_ro[15]
+ mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18] mgmt_rdata_ro[19] mgmt_rdata_ro[20]
+ mgmt_rdata_ro[21] mgmt_rdata_ro[22] mgmt_rdata_ro[23] mgmt_rdata_ro[24] mgmt_rdata_ro[25]
+ mgmt_rdata_ro[26] mgmt_rdata_ro[27] mgmt_rdata_ro[28] mgmt_rdata_ro[29] mgmt_rdata_ro[30]
+ mgmt_rdata_ro[31] VPWR VGND sram_1rw1r_32_256_8_sky130
XFILLER_156_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_300_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_310_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_289_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_302_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_clk0 mgmt_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_323_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[6] mgmt_addr_ro[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSRAM_1 mgmt_wdata[0] mgmt_wdata[1] mgmt_wdata[2] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wdata[10] mgmt_wdata[11]
+ mgmt_wdata[12] mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17]
+ mgmt_wdata[18] mgmt_wdata[19] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[30] mgmt_wdata[31] mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3]
+ mgmt_addr[4] mgmt_addr[5] mgmt_addr[6] mgmt_addr[7] SRAM_1/addr1[0] SRAM_1/addr1[1]
+ SRAM_1/addr1[2] SRAM_1/addr1[3] SRAM_1/addr1[4] SRAM_1/addr1[5] SRAM_1/addr1[6]
+ SRAM_1/addr1[7] mgmt_ena[1] SRAM_1/csb1 mgmt_wen[1] mgmt_clk SRAM_1/clk1 mgmt_wen_mask[4]
+ mgmt_wen_mask[5] mgmt_wen_mask[6] mgmt_wen_mask[7] mgmt_rdata[32] mgmt_rdata[33]
+ mgmt_rdata[34] mgmt_rdata[35] mgmt_rdata[36] mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39]
+ mgmt_rdata[40] mgmt_rdata[41] mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45]
+ mgmt_rdata[46] mgmt_rdata[47] mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[50] mgmt_rdata[51]
+ mgmt_rdata[52] mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56] mgmt_rdata[57]
+ mgmt_rdata[58] mgmt_rdata[59] mgmt_rdata[60] mgmt_rdata[61] mgmt_rdata[62] mgmt_rdata[63]
+ SRAM_1/dout1[0] SRAM_1/dout1[1] SRAM_1/dout1[2] SRAM_1/dout1[3] SRAM_1/dout1[4]
+ SRAM_1/dout1[5] SRAM_1/dout1[6] SRAM_1/dout1[7] SRAM_1/dout1[8] SRAM_1/dout1[9]
+ SRAM_1/dout1[10] SRAM_1/dout1[11] SRAM_1/dout1[12] SRAM_1/dout1[13] SRAM_1/dout1[14]
+ SRAM_1/dout1[15] SRAM_1/dout1[16] SRAM_1/dout1[17] SRAM_1/dout1[18] SRAM_1/dout1[19]
+ SRAM_1/dout1[20] SRAM_1/dout1[21] SRAM_1/dout1[22] SRAM_1/dout1[23] SRAM_1/dout1[24]
+ SRAM_1/dout1[25] SRAM_1/dout1[26] SRAM_1/dout1[27] SRAM_1/dout1[28] SRAM_1/dout1[29]
+ SRAM_1/dout1[30] SRAM_1/dout1[31] VPWR VGND sram_1rw1r_32_256_8_sky130
XFILLER_305_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_301_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_302_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_327_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_295_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[29] mgmt_wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_313_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_259_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_clk1 mgmt_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_310_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[5] mgmt_addr_ro[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[28] mgmt_wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_277_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_313_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_308_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_308_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_319_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_316_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_321_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_266_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_addr1[4] mgmt_addr_ro[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_313_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_304_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_289_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_327_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[27] mgmt_wdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_324_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_324_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_296_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_326_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_335_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_wmask0[3] mgmt_wen_mask[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_308_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[3] mgmt_addr_ro[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_289_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_327_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_SRAM_0_din0[26] mgmt_wdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_339_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_337_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_289_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_271_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_319_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_334_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_325_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_wmask0[2] mgmt_wen_mask[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_316_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_307_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[2] mgmt_addr_ro[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_321_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_289_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_csb0 mgmt_ena[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_SRAM_0_din0[25] mgmt_wdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_338_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_291_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_264_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_334_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_270_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_wmask0[1] mgmt_wen_mask[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_316_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[1] mgmt_addr_ro[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_314_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_310_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_264_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[24] mgmt_wdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_264_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_329_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_261_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_wmask0[0] mgmt_wen_mask[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_307_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[0] mgmt_addr_ro[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[23] mgmt_wdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_280_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_280_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_274_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_337_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_319_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_287_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_306_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_278_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_0_din0[22] mgmt_wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_294_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_285_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_314_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_319_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_340_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_286_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_322_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_297_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_0_din0[21] mgmt_wdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_294_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_291_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_273_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_255_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_292_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_din0[9] mgmt_wdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_305_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[19] mgmt_wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[20] mgmt_wdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_277_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_259_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_334_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_335_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[8] mgmt_wdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_300_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_297_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_din0[18] mgmt_wdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_294_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_276_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_267_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_334_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_340_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_300_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_313_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_304_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_SRAM_1_din0[7] mgmt_wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[17] mgmt_wdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_310_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_285_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_267_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[3] mgmt_wen_mask[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_258_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_333_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_300_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_252_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_330_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_addr0[7] mgmt_addr[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_340_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_303_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_SRAM_1_din0[6] mgmt_wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_289_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[16] mgmt_wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_267_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[2] mgmt_wen_mask[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_314_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_330_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_309_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_addr0[6] mgmt_addr[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_276_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_312_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[5] mgmt_wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_306_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_297_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_din0[15] mgmt_wdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_317_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[1] mgmt_wen_mask[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_314_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_314_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_325_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_307_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_addr0[5] mgmt_addr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_292_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[31] mgmt_wdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[4] mgmt_wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_322_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_276_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_297_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[14] mgmt_wdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_317_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[0] mgmt_wen_mask[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_264_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_addr0[4] mgmt_addr[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_306_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_336_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_din0[30] mgmt_wdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_din0[3] mgmt_wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[13] mgmt_wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_328_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_csb0 mgmt_ena[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_301_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_281_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_249_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_299_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_251_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_addr0[3] mgmt_addr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_306_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_336_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_din0[2] mgmt_wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[12] mgmt_wdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_300_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_csb1 mgmt_ena_ro VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_337_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_254_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_249_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_265_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_addr0[2] mgmt_addr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_din0[1] mgmt_wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[11] mgmt_wdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_282_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_270_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_258_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_327_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_255_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_addr0[1] mgmt_addr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_276_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_din0[0] mgmt_wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_317_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[10] mgmt_wdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_din0[9] mgmt_wdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_267_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_293_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_268_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_290_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_257_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_263_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_318_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_309_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_330_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_addr0[0] mgmt_addr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_312_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_297_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_287_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_web0 mgmt_wen[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_312_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_din0[8] mgmt_wdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_284_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_290_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_309_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_292_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[19] mgmt_wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_298_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[7] mgmt_wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_285_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_339_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_295_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_306_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[18] mgmt_wdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[6] mgmt_wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_287_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_315_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_334_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_257_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_330_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_321_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[17] mgmt_wdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_312_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[5] mgmt_wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_308_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_293_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_266_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_addr0[7] mgmt_addr[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_0_din0[16] mgmt_wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_320_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_338_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_297_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[4] mgmt_wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_320_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_304_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[6] mgmt_addr[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[15] mgmt_wdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_320_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_311_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_302_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_296_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_287_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[3] mgmt_wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_307_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_clk0 mgmt_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_304_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_263_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_SRAM_0_addr0[5] mgmt_addr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_333_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_254_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[31] mgmt_wdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_306_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[14] mgmt_wdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_282_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_311_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_312_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[2] mgmt_wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_287_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_307_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_323_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_290_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_din0[29] mgmt_wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_335_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_320_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_256_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[4] mgmt_addr[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_0_din0[30] mgmt_wdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_317_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_323_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[13] mgmt_wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_305_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_336_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[1] mgmt_wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_287_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_288_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_323_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_286_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_269_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_318_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_318_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[28] mgmt_wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_0_addr0[3] mgmt_addr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_296_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_0_din0[12] mgmt_wdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_305_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_326_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[0] mgmt_wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_334_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_336_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_din0[27] mgmt_wdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_addr0[2] mgmt_addr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_309_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[11] mgmt_wdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_305_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_329_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_272_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[26] mgmt_wdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_260_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_335_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_SRAM_0_addr0[1] mgmt_addr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_326_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_254_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[10] mgmt_wdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_266_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_302_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_334_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_258_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_283_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_SRAM_1_din0[25] mgmt_wdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_280_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[0] mgmt_addr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_262_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_308_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_266_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_320_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_282_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_web0 mgmt_wen[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_302_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_339_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_274_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_274_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_290_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_277_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[24] mgmt_wdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_280_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_269_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_262_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_282_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_277_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_293_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_290_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_290_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_275_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

