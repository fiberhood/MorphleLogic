// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module mgmt_protect(caravel_clk, caravel_clk2, caravel_rstn, mprj_cyc_o_core, mprj_cyc_o_user, mprj_stb_o_core, mprj_stb_o_user, mprj_we_o_core, mprj_we_o_user, user1_vcc_powergood, user1_vdd_powergood, user2_vcc_powergood, user2_vdd_powergood, user_clock, user_clock2, user_reset, user_resetn, vccd, vssd, vccd1, vssd1, vccd2, vssd2, vdda1, vssa1, vdda2, vssa2, la_data_in_core, la_data_in_mprj, la_data_out_core, la_data_out_mprj, la_oen_core, la_oen_mprj, mprj_adr_o_core, mprj_adr_o_user, mprj_dat_o_core, mprj_dat_o_user, mprj_sel_o_core, mprj_sel_o_user);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  input caravel_clk;
  input caravel_clk2;
  input caravel_rstn;
  output [127:0] la_data_in_core;
  output [127:0] la_data_in_mprj;
  wire \la_data_in_mprj_bar[0] ;
  wire \la_data_in_mprj_bar[100] ;
  wire \la_data_in_mprj_bar[101] ;
  wire \la_data_in_mprj_bar[102] ;
  wire \la_data_in_mprj_bar[103] ;
  wire \la_data_in_mprj_bar[104] ;
  wire \la_data_in_mprj_bar[105] ;
  wire \la_data_in_mprj_bar[106] ;
  wire \la_data_in_mprj_bar[107] ;
  wire \la_data_in_mprj_bar[108] ;
  wire \la_data_in_mprj_bar[109] ;
  wire \la_data_in_mprj_bar[10] ;
  wire \la_data_in_mprj_bar[110] ;
  wire \la_data_in_mprj_bar[111] ;
  wire \la_data_in_mprj_bar[112] ;
  wire \la_data_in_mprj_bar[113] ;
  wire \la_data_in_mprj_bar[114] ;
  wire \la_data_in_mprj_bar[115] ;
  wire \la_data_in_mprj_bar[116] ;
  wire \la_data_in_mprj_bar[117] ;
  wire \la_data_in_mprj_bar[118] ;
  wire \la_data_in_mprj_bar[119] ;
  wire \la_data_in_mprj_bar[11] ;
  wire \la_data_in_mprj_bar[120] ;
  wire \la_data_in_mprj_bar[121] ;
  wire \la_data_in_mprj_bar[122] ;
  wire \la_data_in_mprj_bar[123] ;
  wire \la_data_in_mprj_bar[124] ;
  wire \la_data_in_mprj_bar[125] ;
  wire \la_data_in_mprj_bar[126] ;
  wire \la_data_in_mprj_bar[127] ;
  wire \la_data_in_mprj_bar[12] ;
  wire \la_data_in_mprj_bar[13] ;
  wire \la_data_in_mprj_bar[14] ;
  wire \la_data_in_mprj_bar[15] ;
  wire \la_data_in_mprj_bar[16] ;
  wire \la_data_in_mprj_bar[17] ;
  wire \la_data_in_mprj_bar[18] ;
  wire \la_data_in_mprj_bar[19] ;
  wire \la_data_in_mprj_bar[1] ;
  wire \la_data_in_mprj_bar[20] ;
  wire \la_data_in_mprj_bar[21] ;
  wire \la_data_in_mprj_bar[22] ;
  wire \la_data_in_mprj_bar[23] ;
  wire \la_data_in_mprj_bar[24] ;
  wire \la_data_in_mprj_bar[25] ;
  wire \la_data_in_mprj_bar[26] ;
  wire \la_data_in_mprj_bar[27] ;
  wire \la_data_in_mprj_bar[28] ;
  wire \la_data_in_mprj_bar[29] ;
  wire \la_data_in_mprj_bar[2] ;
  wire \la_data_in_mprj_bar[30] ;
  wire \la_data_in_mprj_bar[31] ;
  wire \la_data_in_mprj_bar[32] ;
  wire \la_data_in_mprj_bar[33] ;
  wire \la_data_in_mprj_bar[34] ;
  wire \la_data_in_mprj_bar[35] ;
  wire \la_data_in_mprj_bar[36] ;
  wire \la_data_in_mprj_bar[37] ;
  wire \la_data_in_mprj_bar[38] ;
  wire \la_data_in_mprj_bar[39] ;
  wire \la_data_in_mprj_bar[3] ;
  wire \la_data_in_mprj_bar[40] ;
  wire \la_data_in_mprj_bar[41] ;
  wire \la_data_in_mprj_bar[42] ;
  wire \la_data_in_mprj_bar[43] ;
  wire \la_data_in_mprj_bar[44] ;
  wire \la_data_in_mprj_bar[45] ;
  wire \la_data_in_mprj_bar[46] ;
  wire \la_data_in_mprj_bar[47] ;
  wire \la_data_in_mprj_bar[48] ;
  wire \la_data_in_mprj_bar[49] ;
  wire \la_data_in_mprj_bar[4] ;
  wire \la_data_in_mprj_bar[50] ;
  wire \la_data_in_mprj_bar[51] ;
  wire \la_data_in_mprj_bar[52] ;
  wire \la_data_in_mprj_bar[53] ;
  wire \la_data_in_mprj_bar[54] ;
  wire \la_data_in_mprj_bar[55] ;
  wire \la_data_in_mprj_bar[56] ;
  wire \la_data_in_mprj_bar[57] ;
  wire \la_data_in_mprj_bar[58] ;
  wire \la_data_in_mprj_bar[59] ;
  wire \la_data_in_mprj_bar[5] ;
  wire \la_data_in_mprj_bar[60] ;
  wire \la_data_in_mprj_bar[61] ;
  wire \la_data_in_mprj_bar[62] ;
  wire \la_data_in_mprj_bar[63] ;
  wire \la_data_in_mprj_bar[64] ;
  wire \la_data_in_mprj_bar[65] ;
  wire \la_data_in_mprj_bar[66] ;
  wire \la_data_in_mprj_bar[67] ;
  wire \la_data_in_mprj_bar[68] ;
  wire \la_data_in_mprj_bar[69] ;
  wire \la_data_in_mprj_bar[6] ;
  wire \la_data_in_mprj_bar[70] ;
  wire \la_data_in_mprj_bar[71] ;
  wire \la_data_in_mprj_bar[72] ;
  wire \la_data_in_mprj_bar[73] ;
  wire \la_data_in_mprj_bar[74] ;
  wire \la_data_in_mprj_bar[75] ;
  wire \la_data_in_mprj_bar[76] ;
  wire \la_data_in_mprj_bar[77] ;
  wire \la_data_in_mprj_bar[78] ;
  wire \la_data_in_mprj_bar[79] ;
  wire \la_data_in_mprj_bar[7] ;
  wire \la_data_in_mprj_bar[80] ;
  wire \la_data_in_mprj_bar[81] ;
  wire \la_data_in_mprj_bar[82] ;
  wire \la_data_in_mprj_bar[83] ;
  wire \la_data_in_mprj_bar[84] ;
  wire \la_data_in_mprj_bar[85] ;
  wire \la_data_in_mprj_bar[86] ;
  wire \la_data_in_mprj_bar[87] ;
  wire \la_data_in_mprj_bar[88] ;
  wire \la_data_in_mprj_bar[89] ;
  wire \la_data_in_mprj_bar[8] ;
  wire \la_data_in_mprj_bar[90] ;
  wire \la_data_in_mprj_bar[91] ;
  wire \la_data_in_mprj_bar[92] ;
  wire \la_data_in_mprj_bar[93] ;
  wire \la_data_in_mprj_bar[94] ;
  wire \la_data_in_mprj_bar[95] ;
  wire \la_data_in_mprj_bar[96] ;
  wire \la_data_in_mprj_bar[97] ;
  wire \la_data_in_mprj_bar[98] ;
  wire \la_data_in_mprj_bar[99] ;
  wire \la_data_in_mprj_bar[9] ;
  input [127:0] la_data_out_core;
  input [127:0] la_data_out_mprj;
  output [127:0] la_oen_core;
  input [127:0] la_oen_mprj;
  wire mprj2_logic1;
  wire mprj2_vdd_logic1;
  input [31:0] mprj_adr_o_core;
  output [31:0] mprj_adr_o_user;
  input mprj_cyc_o_core;
  output mprj_cyc_o_user;
  input [31:0] mprj_dat_o_core;
  output [31:0] mprj_dat_o_user;
  wire \mprj_logic1[0] ;
  wire \mprj_logic1[100] ;
  wire \mprj_logic1[101] ;
  wire \mprj_logic1[102] ;
  wire \mprj_logic1[103] ;
  wire \mprj_logic1[104] ;
  wire \mprj_logic1[105] ;
  wire \mprj_logic1[106] ;
  wire \mprj_logic1[107] ;
  wire \mprj_logic1[108] ;
  wire \mprj_logic1[109] ;
  wire \mprj_logic1[10] ;
  wire \mprj_logic1[110] ;
  wire \mprj_logic1[111] ;
  wire \mprj_logic1[112] ;
  wire \mprj_logic1[113] ;
  wire \mprj_logic1[114] ;
  wire \mprj_logic1[115] ;
  wire \mprj_logic1[116] ;
  wire \mprj_logic1[117] ;
  wire \mprj_logic1[118] ;
  wire \mprj_logic1[119] ;
  wire \mprj_logic1[11] ;
  wire \mprj_logic1[120] ;
  wire \mprj_logic1[121] ;
  wire \mprj_logic1[122] ;
  wire \mprj_logic1[123] ;
  wire \mprj_logic1[124] ;
  wire \mprj_logic1[125] ;
  wire \mprj_logic1[126] ;
  wire \mprj_logic1[127] ;
  wire \mprj_logic1[128] ;
  wire \mprj_logic1[129] ;
  wire \mprj_logic1[12] ;
  wire \mprj_logic1[130] ;
  wire \mprj_logic1[131] ;
  wire \mprj_logic1[132] ;
  wire \mprj_logic1[133] ;
  wire \mprj_logic1[134] ;
  wire \mprj_logic1[135] ;
  wire \mprj_logic1[136] ;
  wire \mprj_logic1[137] ;
  wire \mprj_logic1[138] ;
  wire \mprj_logic1[139] ;
  wire \mprj_logic1[13] ;
  wire \mprj_logic1[140] ;
  wire \mprj_logic1[141] ;
  wire \mprj_logic1[142] ;
  wire \mprj_logic1[143] ;
  wire \mprj_logic1[144] ;
  wire \mprj_logic1[145] ;
  wire \mprj_logic1[146] ;
  wire \mprj_logic1[147] ;
  wire \mprj_logic1[148] ;
  wire \mprj_logic1[149] ;
  wire \mprj_logic1[14] ;
  wire \mprj_logic1[150] ;
  wire \mprj_logic1[151] ;
  wire \mprj_logic1[152] ;
  wire \mprj_logic1[153] ;
  wire \mprj_logic1[154] ;
  wire \mprj_logic1[155] ;
  wire \mprj_logic1[156] ;
  wire \mprj_logic1[157] ;
  wire \mprj_logic1[158] ;
  wire \mprj_logic1[159] ;
  wire \mprj_logic1[15] ;
  wire \mprj_logic1[160] ;
  wire \mprj_logic1[161] ;
  wire \mprj_logic1[162] ;
  wire \mprj_logic1[163] ;
  wire \mprj_logic1[164] ;
  wire \mprj_logic1[165] ;
  wire \mprj_logic1[166] ;
  wire \mprj_logic1[167] ;
  wire \mprj_logic1[168] ;
  wire \mprj_logic1[169] ;
  wire \mprj_logic1[16] ;
  wire \mprj_logic1[170] ;
  wire \mprj_logic1[171] ;
  wire \mprj_logic1[172] ;
  wire \mprj_logic1[173] ;
  wire \mprj_logic1[174] ;
  wire \mprj_logic1[175] ;
  wire \mprj_logic1[176] ;
  wire \mprj_logic1[177] ;
  wire \mprj_logic1[178] ;
  wire \mprj_logic1[179] ;
  wire \mprj_logic1[17] ;
  wire \mprj_logic1[180] ;
  wire \mprj_logic1[181] ;
  wire \mprj_logic1[182] ;
  wire \mprj_logic1[183] ;
  wire \mprj_logic1[184] ;
  wire \mprj_logic1[185] ;
  wire \mprj_logic1[186] ;
  wire \mprj_logic1[187] ;
  wire \mprj_logic1[188] ;
  wire \mprj_logic1[189] ;
  wire \mprj_logic1[18] ;
  wire \mprj_logic1[190] ;
  wire \mprj_logic1[191] ;
  wire \mprj_logic1[192] ;
  wire \mprj_logic1[193] ;
  wire \mprj_logic1[194] ;
  wire \mprj_logic1[195] ;
  wire \mprj_logic1[196] ;
  wire \mprj_logic1[197] ;
  wire \mprj_logic1[198] ;
  wire \mprj_logic1[199] ;
  wire \mprj_logic1[19] ;
  wire \mprj_logic1[1] ;
  wire \mprj_logic1[200] ;
  wire \mprj_logic1[201] ;
  wire \mprj_logic1[202] ;
  wire \mprj_logic1[203] ;
  wire \mprj_logic1[204] ;
  wire \mprj_logic1[205] ;
  wire \mprj_logic1[206] ;
  wire \mprj_logic1[207] ;
  wire \mprj_logic1[208] ;
  wire \mprj_logic1[209] ;
  wire \mprj_logic1[20] ;
  wire \mprj_logic1[210] ;
  wire \mprj_logic1[211] ;
  wire \mprj_logic1[212] ;
  wire \mprj_logic1[213] ;
  wire \mprj_logic1[214] ;
  wire \mprj_logic1[215] ;
  wire \mprj_logic1[216] ;
  wire \mprj_logic1[217] ;
  wire \mprj_logic1[218] ;
  wire \mprj_logic1[219] ;
  wire \mprj_logic1[21] ;
  wire \mprj_logic1[220] ;
  wire \mprj_logic1[221] ;
  wire \mprj_logic1[222] ;
  wire \mprj_logic1[223] ;
  wire \mprj_logic1[224] ;
  wire \mprj_logic1[225] ;
  wire \mprj_logic1[226] ;
  wire \mprj_logic1[227] ;
  wire \mprj_logic1[228] ;
  wire \mprj_logic1[229] ;
  wire \mprj_logic1[22] ;
  wire \mprj_logic1[230] ;
  wire \mprj_logic1[231] ;
  wire \mprj_logic1[232] ;
  wire \mprj_logic1[233] ;
  wire \mprj_logic1[234] ;
  wire \mprj_logic1[235] ;
  wire \mprj_logic1[236] ;
  wire \mprj_logic1[237] ;
  wire \mprj_logic1[238] ;
  wire \mprj_logic1[239] ;
  wire \mprj_logic1[23] ;
  wire \mprj_logic1[240] ;
  wire \mprj_logic1[241] ;
  wire \mprj_logic1[242] ;
  wire \mprj_logic1[243] ;
  wire \mprj_logic1[244] ;
  wire \mprj_logic1[245] ;
  wire \mprj_logic1[246] ;
  wire \mprj_logic1[247] ;
  wire \mprj_logic1[248] ;
  wire \mprj_logic1[249] ;
  wire \mprj_logic1[24] ;
  wire \mprj_logic1[250] ;
  wire \mprj_logic1[251] ;
  wire \mprj_logic1[252] ;
  wire \mprj_logic1[253] ;
  wire \mprj_logic1[254] ;
  wire \mprj_logic1[255] ;
  wire \mprj_logic1[256] ;
  wire \mprj_logic1[257] ;
  wire \mprj_logic1[258] ;
  wire \mprj_logic1[259] ;
  wire \mprj_logic1[25] ;
  wire \mprj_logic1[260] ;
  wire \mprj_logic1[261] ;
  wire \mprj_logic1[262] ;
  wire \mprj_logic1[263] ;
  wire \mprj_logic1[264] ;
  wire \mprj_logic1[265] ;
  wire \mprj_logic1[266] ;
  wire \mprj_logic1[267] ;
  wire \mprj_logic1[268] ;
  wire \mprj_logic1[269] ;
  wire \mprj_logic1[26] ;
  wire \mprj_logic1[270] ;
  wire \mprj_logic1[271] ;
  wire \mprj_logic1[272] ;
  wire \mprj_logic1[273] ;
  wire \mprj_logic1[274] ;
  wire \mprj_logic1[275] ;
  wire \mprj_logic1[276] ;
  wire \mprj_logic1[277] ;
  wire \mprj_logic1[278] ;
  wire \mprj_logic1[279] ;
  wire \mprj_logic1[27] ;
  wire \mprj_logic1[280] ;
  wire \mprj_logic1[281] ;
  wire \mprj_logic1[282] ;
  wire \mprj_logic1[283] ;
  wire \mprj_logic1[284] ;
  wire \mprj_logic1[285] ;
  wire \mprj_logic1[286] ;
  wire \mprj_logic1[287] ;
  wire \mprj_logic1[288] ;
  wire \mprj_logic1[289] ;
  wire \mprj_logic1[28] ;
  wire \mprj_logic1[290] ;
  wire \mprj_logic1[291] ;
  wire \mprj_logic1[292] ;
  wire \mprj_logic1[293] ;
  wire \mprj_logic1[294] ;
  wire \mprj_logic1[295] ;
  wire \mprj_logic1[296] ;
  wire \mprj_logic1[297] ;
  wire \mprj_logic1[298] ;
  wire \mprj_logic1[299] ;
  wire \mprj_logic1[29] ;
  wire \mprj_logic1[2] ;
  wire \mprj_logic1[300] ;
  wire \mprj_logic1[301] ;
  wire \mprj_logic1[302] ;
  wire \mprj_logic1[303] ;
  wire \mprj_logic1[304] ;
  wire \mprj_logic1[305] ;
  wire \mprj_logic1[306] ;
  wire \mprj_logic1[307] ;
  wire \mprj_logic1[308] ;
  wire \mprj_logic1[309] ;
  wire \mprj_logic1[30] ;
  wire \mprj_logic1[310] ;
  wire \mprj_logic1[311] ;
  wire \mprj_logic1[312] ;
  wire \mprj_logic1[313] ;
  wire \mprj_logic1[314] ;
  wire \mprj_logic1[315] ;
  wire \mprj_logic1[316] ;
  wire \mprj_logic1[317] ;
  wire \mprj_logic1[318] ;
  wire \mprj_logic1[319] ;
  wire \mprj_logic1[31] ;
  wire \mprj_logic1[320] ;
  wire \mprj_logic1[321] ;
  wire \mprj_logic1[322] ;
  wire \mprj_logic1[323] ;
  wire \mprj_logic1[324] ;
  wire \mprj_logic1[325] ;
  wire \mprj_logic1[326] ;
  wire \mprj_logic1[327] ;
  wire \mprj_logic1[328] ;
  wire \mprj_logic1[329] ;
  wire \mprj_logic1[32] ;
  wire \mprj_logic1[330] ;
  wire \mprj_logic1[331] ;
  wire \mprj_logic1[332] ;
  wire \mprj_logic1[333] ;
  wire \mprj_logic1[334] ;
  wire \mprj_logic1[335] ;
  wire \mprj_logic1[336] ;
  wire \mprj_logic1[337] ;
  wire \mprj_logic1[338] ;
  wire \mprj_logic1[339] ;
  wire \mprj_logic1[33] ;
  wire \mprj_logic1[340] ;
  wire \mprj_logic1[341] ;
  wire \mprj_logic1[342] ;
  wire \mprj_logic1[343] ;
  wire \mprj_logic1[344] ;
  wire \mprj_logic1[345] ;
  wire \mprj_logic1[346] ;
  wire \mprj_logic1[347] ;
  wire \mprj_logic1[348] ;
  wire \mprj_logic1[349] ;
  wire \mprj_logic1[34] ;
  wire \mprj_logic1[350] ;
  wire \mprj_logic1[351] ;
  wire \mprj_logic1[352] ;
  wire \mprj_logic1[353] ;
  wire \mprj_logic1[354] ;
  wire \mprj_logic1[355] ;
  wire \mprj_logic1[356] ;
  wire \mprj_logic1[357] ;
  wire \mprj_logic1[358] ;
  wire \mprj_logic1[359] ;
  wire \mprj_logic1[35] ;
  wire \mprj_logic1[360] ;
  wire \mprj_logic1[361] ;
  wire \mprj_logic1[362] ;
  wire \mprj_logic1[363] ;
  wire \mprj_logic1[364] ;
  wire \mprj_logic1[365] ;
  wire \mprj_logic1[366] ;
  wire \mprj_logic1[367] ;
  wire \mprj_logic1[368] ;
  wire \mprj_logic1[369] ;
  wire \mprj_logic1[36] ;
  wire \mprj_logic1[370] ;
  wire \mprj_logic1[371] ;
  wire \mprj_logic1[372] ;
  wire \mprj_logic1[373] ;
  wire \mprj_logic1[374] ;
  wire \mprj_logic1[375] ;
  wire \mprj_logic1[376] ;
  wire \mprj_logic1[377] ;
  wire \mprj_logic1[378] ;
  wire \mprj_logic1[379] ;
  wire \mprj_logic1[37] ;
  wire \mprj_logic1[380] ;
  wire \mprj_logic1[381] ;
  wire \mprj_logic1[382] ;
  wire \mprj_logic1[383] ;
  wire \mprj_logic1[384] ;
  wire \mprj_logic1[385] ;
  wire \mprj_logic1[386] ;
  wire \mprj_logic1[387] ;
  wire \mprj_logic1[388] ;
  wire \mprj_logic1[389] ;
  wire \mprj_logic1[38] ;
  wire \mprj_logic1[390] ;
  wire \mprj_logic1[391] ;
  wire \mprj_logic1[392] ;
  wire \mprj_logic1[393] ;
  wire \mprj_logic1[394] ;
  wire \mprj_logic1[395] ;
  wire \mprj_logic1[396] ;
  wire \mprj_logic1[397] ;
  wire \mprj_logic1[398] ;
  wire \mprj_logic1[399] ;
  wire \mprj_logic1[39] ;
  wire \mprj_logic1[3] ;
  wire \mprj_logic1[400] ;
  wire \mprj_logic1[401] ;
  wire \mprj_logic1[402] ;
  wire \mprj_logic1[403] ;
  wire \mprj_logic1[404] ;
  wire \mprj_logic1[405] ;
  wire \mprj_logic1[406] ;
  wire \mprj_logic1[407] ;
  wire \mprj_logic1[408] ;
  wire \mprj_logic1[409] ;
  wire \mprj_logic1[40] ;
  wire \mprj_logic1[410] ;
  wire \mprj_logic1[411] ;
  wire \mprj_logic1[412] ;
  wire \mprj_logic1[413] ;
  wire \mprj_logic1[414] ;
  wire \mprj_logic1[415] ;
  wire \mprj_logic1[416] ;
  wire \mprj_logic1[417] ;
  wire \mprj_logic1[418] ;
  wire \mprj_logic1[419] ;
  wire \mprj_logic1[41] ;
  wire \mprj_logic1[420] ;
  wire \mprj_logic1[421] ;
  wire \mprj_logic1[422] ;
  wire \mprj_logic1[423] ;
  wire \mprj_logic1[424] ;
  wire \mprj_logic1[425] ;
  wire \mprj_logic1[426] ;
  wire \mprj_logic1[427] ;
  wire \mprj_logic1[428] ;
  wire \mprj_logic1[429] ;
  wire \mprj_logic1[42] ;
  wire \mprj_logic1[430] ;
  wire \mprj_logic1[431] ;
  wire \mprj_logic1[432] ;
  wire \mprj_logic1[433] ;
  wire \mprj_logic1[434] ;
  wire \mprj_logic1[435] ;
  wire \mprj_logic1[436] ;
  wire \mprj_logic1[437] ;
  wire \mprj_logic1[438] ;
  wire \mprj_logic1[439] ;
  wire \mprj_logic1[43] ;
  wire \mprj_logic1[440] ;
  wire \mprj_logic1[441] ;
  wire \mprj_logic1[442] ;
  wire \mprj_logic1[443] ;
  wire \mprj_logic1[444] ;
  wire \mprj_logic1[445] ;
  wire \mprj_logic1[446] ;
  wire \mprj_logic1[447] ;
  wire \mprj_logic1[448] ;
  wire \mprj_logic1[449] ;
  wire \mprj_logic1[44] ;
  wire \mprj_logic1[450] ;
  wire \mprj_logic1[451] ;
  wire \mprj_logic1[452] ;
  wire \mprj_logic1[453] ;
  wire \mprj_logic1[454] ;
  wire \mprj_logic1[455] ;
  wire \mprj_logic1[456] ;
  wire \mprj_logic1[457] ;
  wire \mprj_logic1[458] ;
  wire \mprj_logic1[45] ;
  wire \mprj_logic1[46] ;
  wire \mprj_logic1[47] ;
  wire \mprj_logic1[48] ;
  wire \mprj_logic1[49] ;
  wire \mprj_logic1[4] ;
  wire \mprj_logic1[50] ;
  wire \mprj_logic1[51] ;
  wire \mprj_logic1[52] ;
  wire \mprj_logic1[53] ;
  wire \mprj_logic1[54] ;
  wire \mprj_logic1[55] ;
  wire \mprj_logic1[56] ;
  wire \mprj_logic1[57] ;
  wire \mprj_logic1[58] ;
  wire \mprj_logic1[59] ;
  wire \mprj_logic1[5] ;
  wire \mprj_logic1[60] ;
  wire \mprj_logic1[61] ;
  wire \mprj_logic1[62] ;
  wire \mprj_logic1[63] ;
  wire \mprj_logic1[64] ;
  wire \mprj_logic1[65] ;
  wire \mprj_logic1[66] ;
  wire \mprj_logic1[67] ;
  wire \mprj_logic1[68] ;
  wire \mprj_logic1[69] ;
  wire \mprj_logic1[6] ;
  wire \mprj_logic1[70] ;
  wire \mprj_logic1[71] ;
  wire \mprj_logic1[72] ;
  wire \mprj_logic1[73] ;
  wire \mprj_logic1[74] ;
  wire \mprj_logic1[75] ;
  wire \mprj_logic1[76] ;
  wire \mprj_logic1[77] ;
  wire \mprj_logic1[78] ;
  wire \mprj_logic1[79] ;
  wire \mprj_logic1[7] ;
  wire \mprj_logic1[80] ;
  wire \mprj_logic1[81] ;
  wire \mprj_logic1[82] ;
  wire \mprj_logic1[83] ;
  wire \mprj_logic1[84] ;
  wire \mprj_logic1[85] ;
  wire \mprj_logic1[86] ;
  wire \mprj_logic1[87] ;
  wire \mprj_logic1[88] ;
  wire \mprj_logic1[89] ;
  wire \mprj_logic1[8] ;
  wire \mprj_logic1[90] ;
  wire \mprj_logic1[91] ;
  wire \mprj_logic1[92] ;
  wire \mprj_logic1[93] ;
  wire \mprj_logic1[94] ;
  wire \mprj_logic1[95] ;
  wire \mprj_logic1[96] ;
  wire \mprj_logic1[97] ;
  wire \mprj_logic1[98] ;
  wire \mprj_logic1[99] ;
  wire \mprj_logic1[9] ;
  input [3:0] mprj_sel_o_core;
  output [3:0] mprj_sel_o_user;
  input mprj_stb_o_core;
  output mprj_stb_o_user;
  wire mprj_vdd_logic1;
  input mprj_we_o_core;
  output mprj_we_o_user;
  output user1_vcc_powergood;
  output user1_vdd_powergood;
  output user2_vcc_powergood;
  output user2_vdd_powergood;
  output user_clock;
  output user_clock2;
  output user_reset;
  output user_resetn;
  input vccd;
  input vccd1;
  input vccd2;
  input vdda1;
  input vdda2;
  input vssa1;
  input vssa2;
  input vssd;
  input vssd1;
  input vssd2;
  sky130_fd_sc_hd__diode_2 ANTENNA__330__A (
    .DIODE(la_oen_mprj[62]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__331__A (
    .DIODE(la_oen_mprj[63]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__332__A (
    .DIODE(la_oen_mprj[64]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__333__A (
    .DIODE(la_oen_mprj[65]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__334__A (
    .DIODE(la_oen_mprj[66]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__335__A (
    .DIODE(la_oen_mprj[67]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__336__A (
    .DIODE(la_oen_mprj[68]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__337__A (
    .DIODE(la_oen_mprj[69]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__338__A (
    .DIODE(la_oen_mprj[70]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__339__A (
    .DIODE(la_oen_mprj[71]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__340__A (
    .DIODE(la_oen_mprj[72]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__341__A (
    .DIODE(la_oen_mprj[73]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__342__A (
    .DIODE(la_oen_mprj[74]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__343__A (
    .DIODE(la_oen_mprj[75]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__344__A (
    .DIODE(la_oen_mprj[76]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__345__A (
    .DIODE(la_oen_mprj[77]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__346__A (
    .DIODE(la_oen_mprj[78]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__347__A (
    .DIODE(la_oen_mprj[79]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__348__A (
    .DIODE(la_oen_mprj[80]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__349__A (
    .DIODE(la_oen_mprj[81]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__350__A (
    .DIODE(la_oen_mprj[82]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__351__A (
    .DIODE(la_oen_mprj[83]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__352__A (
    .DIODE(la_oen_mprj[84]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__353__A (
    .DIODE(la_oen_mprj[85]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__354__A (
    .DIODE(la_oen_mprj[86]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__355__A (
    .DIODE(la_oen_mprj[87]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__356__A (
    .DIODE(la_oen_mprj[88]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__357__A (
    .DIODE(la_oen_mprj[89]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__358__A (
    .DIODE(la_oen_mprj[90]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__359__A (
    .DIODE(la_oen_mprj[91]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__360__A (
    .DIODE(la_oen_mprj[92]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__361__A (
    .DIODE(la_oen_mprj[93]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__362__A (
    .DIODE(la_oen_mprj[94]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__363__A (
    .DIODE(la_oen_mprj[95]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__364__A (
    .DIODE(la_oen_mprj[96]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__365__A (
    .DIODE(la_oen_mprj[97]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__366__A (
    .DIODE(la_oen_mprj[98]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__367__A (
    .DIODE(la_oen_mprj[99]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__368__A (
    .DIODE(la_oen_mprj[100]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__369__A (
    .DIODE(la_oen_mprj[101]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__370__A (
    .DIODE(la_oen_mprj[102]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__371__A (
    .DIODE(la_oen_mprj[103]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__372__A (
    .DIODE(la_oen_mprj[104]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__373__A (
    .DIODE(la_oen_mprj[105]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__374__A (
    .DIODE(la_oen_mprj[106]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__375__A (
    .DIODE(la_oen_mprj[107]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__376__A (
    .DIODE(la_oen_mprj[108]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__377__A (
    .DIODE(la_oen_mprj[109]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__378__A (
    .DIODE(la_oen_mprj[110]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__379__A (
    .DIODE(la_oen_mprj[111]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__380__A (
    .DIODE(la_oen_mprj[112]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__381__A (
    .DIODE(la_oen_mprj[113]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__382__A (
    .DIODE(la_oen_mprj[114]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__383__A (
    .DIODE(la_oen_mprj[115]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__384__A (
    .DIODE(la_oen_mprj[116]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__385__A (
    .DIODE(la_oen_mprj[117]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__386__A (
    .DIODE(la_oen_mprj[118]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__387__A (
    .DIODE(la_oen_mprj[119]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__388__A (
    .DIODE(la_oen_mprj[120]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__389__A (
    .DIODE(la_oen_mprj[121]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__390__A (
    .DIODE(la_oen_mprj[122]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__391__A (
    .DIODE(la_oen_mprj[123]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__392__A (
    .DIODE(la_oen_mprj[124]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__393__A (
    .DIODE(la_oen_mprj[125]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__394__A (
    .DIODE(la_oen_mprj[126]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__395__A (
    .DIODE(la_oen_mprj[127]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__396__A (
    .DIODE(caravel_rstn),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__397__A (
    .DIODE(user_resetn),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__398__A (
    .DIODE(caravel_clk),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__399__A (
    .DIODE(caravel_clk2),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__400__A (
    .DIODE(mprj_cyc_o_core),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__401__A (
    .DIODE(mprj_stb_o_core),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__402__A (
    .DIODE(mprj_we_o_core),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__403__A (
    .DIODE(mprj_sel_o_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__404__A (
    .DIODE(mprj_sel_o_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__405__A (
    .DIODE(mprj_sel_o_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__406__A (
    .DIODE(mprj_sel_o_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__407__A (
    .DIODE(mprj_adr_o_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__408__A (
    .DIODE(mprj_adr_o_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__409__A (
    .DIODE(mprj_adr_o_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__410__A (
    .DIODE(mprj_adr_o_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__411__A (
    .DIODE(mprj_adr_o_core[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__412__A (
    .DIODE(mprj_adr_o_core[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__413__A (
    .DIODE(mprj_adr_o_core[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__414__A (
    .DIODE(mprj_adr_o_core[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__415__A (
    .DIODE(mprj_adr_o_core[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__416__A (
    .DIODE(mprj_adr_o_core[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__417__A (
    .DIODE(mprj_adr_o_core[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__418__A (
    .DIODE(mprj_adr_o_core[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__419__A (
    .DIODE(mprj_adr_o_core[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__420__A (
    .DIODE(mprj_adr_o_core[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__421__A (
    .DIODE(mprj_adr_o_core[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__422__A (
    .DIODE(mprj_adr_o_core[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__423__A (
    .DIODE(mprj_adr_o_core[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__424__A (
    .DIODE(mprj_adr_o_core[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__425__A (
    .DIODE(mprj_adr_o_core[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__426__A (
    .DIODE(mprj_adr_o_core[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__427__A (
    .DIODE(mprj_adr_o_core[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__428__A (
    .DIODE(mprj_adr_o_core[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__429__A (
    .DIODE(mprj_adr_o_core[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__430__A (
    .DIODE(mprj_adr_o_core[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__431__A (
    .DIODE(mprj_adr_o_core[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__432__A (
    .DIODE(mprj_adr_o_core[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__433__A (
    .DIODE(mprj_adr_o_core[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__434__A (
    .DIODE(mprj_adr_o_core[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__435__A (
    .DIODE(mprj_adr_o_core[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__436__A (
    .DIODE(mprj_adr_o_core[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__437__A (
    .DIODE(mprj_adr_o_core[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__438__A (
    .DIODE(mprj_adr_o_core[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__439__A (
    .DIODE(mprj_dat_o_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__440__A (
    .DIODE(mprj_dat_o_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__441__A (
    .DIODE(mprj_dat_o_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__442__A (
    .DIODE(mprj_dat_o_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__443__A (
    .DIODE(mprj_dat_o_core[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__444__A (
    .DIODE(mprj_dat_o_core[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__445__A (
    .DIODE(mprj_dat_o_core[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__446__A (
    .DIODE(mprj_dat_o_core[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__447__A (
    .DIODE(mprj_dat_o_core[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__448__A (
    .DIODE(mprj_dat_o_core[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__449__A (
    .DIODE(mprj_dat_o_core[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__450__A (
    .DIODE(mprj_dat_o_core[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__451__A (
    .DIODE(mprj_dat_o_core[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__452__A (
    .DIODE(mprj_dat_o_core[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__453__A (
    .DIODE(mprj_dat_o_core[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__454__A (
    .DIODE(mprj_dat_o_core[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__455__A (
    .DIODE(mprj_dat_o_core[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__456__A (
    .DIODE(mprj_dat_o_core[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__457__A (
    .DIODE(mprj_dat_o_core[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__458__A (
    .DIODE(mprj_dat_o_core[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__459__A (
    .DIODE(mprj_dat_o_core[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__460__A (
    .DIODE(mprj_dat_o_core[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__461__A (
    .DIODE(mprj_dat_o_core[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__462__A (
    .DIODE(mprj_dat_o_core[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__463__A (
    .DIODE(mprj_dat_o_core[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__464__A (
    .DIODE(mprj_dat_o_core[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__465__A (
    .DIODE(mprj_dat_o_core[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__466__A (
    .DIODE(mprj_dat_o_core[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__467__A (
    .DIODE(mprj_dat_o_core[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__468__A (
    .DIODE(mprj_dat_o_core[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__469__A (
    .DIODE(mprj_dat_o_core[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__470__A (
    .DIODE(mprj_dat_o_core[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__471__A (
    .DIODE(la_data_out_mprj[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__472__A (
    .DIODE(la_data_out_mprj[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__473__A (
    .DIODE(la_data_out_mprj[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__474__A (
    .DIODE(la_data_out_mprj[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__475__A (
    .DIODE(la_data_out_mprj[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__476__A (
    .DIODE(la_data_out_mprj[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__477__A (
    .DIODE(la_data_out_mprj[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__478__A (
    .DIODE(la_data_out_mprj[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__479__A (
    .DIODE(la_data_out_mprj[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__480__A (
    .DIODE(la_data_out_mprj[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__481__A (
    .DIODE(la_data_out_mprj[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__482__A (
    .DIODE(la_data_out_mprj[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__483__A (
    .DIODE(la_data_out_mprj[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__484__A (
    .DIODE(la_data_out_mprj[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__485__A (
    .DIODE(la_data_out_mprj[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__486__A (
    .DIODE(la_data_out_mprj[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__487__A (
    .DIODE(la_data_out_mprj[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__488__A (
    .DIODE(la_data_out_mprj[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__489__A (
    .DIODE(la_data_out_mprj[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__490__A (
    .DIODE(la_data_out_mprj[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__491__A (
    .DIODE(la_data_out_mprj[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__492__A (
    .DIODE(la_data_out_mprj[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__493__A (
    .DIODE(la_data_out_mprj[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__494__A (
    .DIODE(la_data_out_mprj[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__495__A (
    .DIODE(la_data_out_mprj[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__496__A (
    .DIODE(la_data_out_mprj[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__497__A (
    .DIODE(la_data_out_mprj[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__498__A (
    .DIODE(la_data_out_mprj[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__499__A (
    .DIODE(la_data_out_mprj[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__500__A (
    .DIODE(la_data_out_mprj[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__501__A (
    .DIODE(la_data_out_mprj[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__502__A (
    .DIODE(la_data_out_mprj[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__503__A (
    .DIODE(la_data_out_mprj[32]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__504__A (
    .DIODE(la_data_out_mprj[33]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__505__A (
    .DIODE(la_data_out_mprj[34]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__506__A (
    .DIODE(la_data_out_mprj[35]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__507__A (
    .DIODE(la_data_out_mprj[36]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__508__A (
    .DIODE(la_data_out_mprj[37]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__509__A (
    .DIODE(la_data_out_mprj[38]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__510__A (
    .DIODE(la_data_out_mprj[39]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__511__A (
    .DIODE(la_data_out_mprj[40]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__512__A (
    .DIODE(la_data_out_mprj[41]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__513__A (
    .DIODE(la_data_out_mprj[42]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__514__A (
    .DIODE(la_data_out_mprj[43]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__515__A (
    .DIODE(la_data_out_mprj[44]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__516__A (
    .DIODE(la_data_out_mprj[45]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__517__A (
    .DIODE(la_data_out_mprj[46]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__518__A (
    .DIODE(la_data_out_mprj[47]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__519__A (
    .DIODE(la_data_out_mprj[48]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__520__A (
    .DIODE(la_data_out_mprj[49]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__521__A (
    .DIODE(la_data_out_mprj[50]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__522__A (
    .DIODE(la_data_out_mprj[51]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__523__A (
    .DIODE(la_data_out_mprj[52]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__524__A (
    .DIODE(la_data_out_mprj[53]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__525__A (
    .DIODE(la_data_out_mprj[54]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__526__A (
    .DIODE(la_data_out_mprj[55]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__527__A (
    .DIODE(la_data_out_mprj[56]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__528__A (
    .DIODE(la_data_out_mprj[57]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__529__A (
    .DIODE(la_data_out_mprj[58]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__530__A (
    .DIODE(la_data_out_mprj[59]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__531__A (
    .DIODE(la_data_out_mprj[60]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__532__A (
    .DIODE(la_data_out_mprj[61]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__533__A (
    .DIODE(la_data_out_mprj[62]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__534__A (
    .DIODE(la_data_out_mprj[63]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__535__A (
    .DIODE(la_data_out_mprj[64]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__536__A (
    .DIODE(la_data_out_mprj[65]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__537__A (
    .DIODE(la_data_out_mprj[66]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__538__A (
    .DIODE(la_data_out_mprj[67]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__539__A (
    .DIODE(la_data_out_mprj[68]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__540__A (
    .DIODE(la_data_out_mprj[69]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__541__A (
    .DIODE(la_data_out_mprj[70]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__542__A (
    .DIODE(la_data_out_mprj[71]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__543__A (
    .DIODE(la_data_out_mprj[72]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__544__A (
    .DIODE(la_data_out_mprj[73]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__545__A (
    .DIODE(la_data_out_mprj[74]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__546__A (
    .DIODE(la_data_out_mprj[75]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__547__A (
    .DIODE(la_data_out_mprj[76]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__548__A (
    .DIODE(la_data_out_mprj[77]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__549__A (
    .DIODE(la_data_out_mprj[78]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__550__A (
    .DIODE(la_data_out_mprj[79]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__551__A (
    .DIODE(la_data_out_mprj[80]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__552__A (
    .DIODE(la_data_out_mprj[81]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__553__A (
    .DIODE(la_data_out_mprj[82]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__554__A (
    .DIODE(la_data_out_mprj[83]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__555__A (
    .DIODE(la_data_out_mprj[84]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__556__A (
    .DIODE(la_data_out_mprj[85]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__557__A (
    .DIODE(la_data_out_mprj[86]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__558__A (
    .DIODE(la_data_out_mprj[87]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__559__A (
    .DIODE(la_data_out_mprj[88]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__560__A (
    .DIODE(la_data_out_mprj[89]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__561__A (
    .DIODE(la_data_out_mprj[90]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__562__A (
    .DIODE(la_data_out_mprj[91]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__563__A (
    .DIODE(la_data_out_mprj[92]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__564__A (
    .DIODE(la_data_out_mprj[93]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__565__A (
    .DIODE(la_data_out_mprj[94]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__566__A (
    .DIODE(la_data_out_mprj[95]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__567__A (
    .DIODE(la_data_out_mprj[96]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__568__A (
    .DIODE(la_data_out_mprj[97]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__569__A (
    .DIODE(la_data_out_mprj[98]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__570__A (
    .DIODE(la_data_out_mprj[99]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__571__A (
    .DIODE(la_data_out_mprj[100]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__572__A (
    .DIODE(la_data_out_mprj[101]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__573__A (
    .DIODE(la_data_out_mprj[102]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__574__A (
    .DIODE(la_data_out_mprj[103]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__575__A (
    .DIODE(la_data_out_mprj[104]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__576__A (
    .DIODE(la_data_out_mprj[105]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__577__A (
    .DIODE(la_data_out_mprj[106]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__578__A (
    .DIODE(la_data_out_mprj[107]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__579__A (
    .DIODE(la_data_out_mprj[108]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__580__A (
    .DIODE(la_data_out_mprj[109]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__581__A (
    .DIODE(la_data_out_mprj[110]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__582__A (
    .DIODE(la_data_out_mprj[111]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__583__A (
    .DIODE(la_data_out_mprj[112]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__584__A (
    .DIODE(la_data_out_mprj[113]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__585__A (
    .DIODE(la_data_out_mprj[114]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__586__A (
    .DIODE(la_data_out_mprj[115]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__587__A (
    .DIODE(la_data_out_mprj[116]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__588__A (
    .DIODE(la_data_out_mprj[117]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__589__A (
    .DIODE(la_data_out_mprj[118]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__590__A (
    .DIODE(la_data_out_mprj[119]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__591__A (
    .DIODE(la_data_out_mprj[120]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__592__A (
    .DIODE(la_data_out_mprj[121]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__593__A (
    .DIODE(la_data_out_mprj[122]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__594__A (
    .DIODE(la_data_out_mprj[123]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__595__A (
    .DIODE(la_data_out_mprj[124]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__596__A (
    .DIODE(la_data_out_mprj[125]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__597__A (
    .DIODE(la_data_out_mprj[126]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__598__A (
    .DIODE(la_data_out_mprj[127]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__599__A (
    .DIODE(la_oen_mprj[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__600__A (
    .DIODE(la_oen_mprj[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__601__A (
    .DIODE(la_oen_mprj[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__602__A (
    .DIODE(la_oen_mprj[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__603__A (
    .DIODE(la_oen_mprj[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__604__A (
    .DIODE(la_oen_mprj[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__605__A (
    .DIODE(la_oen_mprj[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__606__A (
    .DIODE(la_oen_mprj[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__607__A (
    .DIODE(la_oen_mprj[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__608__A (
    .DIODE(la_oen_mprj[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__609__A (
    .DIODE(la_oen_mprj[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__610__A (
    .DIODE(la_oen_mprj[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__611__A (
    .DIODE(la_oen_mprj[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__612__A (
    .DIODE(la_oen_mprj[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__613__A (
    .DIODE(la_oen_mprj[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__614__A (
    .DIODE(la_oen_mprj[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__615__A (
    .DIODE(la_oen_mprj[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__616__A (
    .DIODE(la_oen_mprj[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__617__A (
    .DIODE(la_oen_mprj[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__618__A (
    .DIODE(la_oen_mprj[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__619__A (
    .DIODE(la_oen_mprj[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__620__A (
    .DIODE(la_oen_mprj[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__621__A (
    .DIODE(la_oen_mprj[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__622__A (
    .DIODE(la_oen_mprj[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__623__A (
    .DIODE(la_oen_mprj[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__624__A (
    .DIODE(la_oen_mprj[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__625__A (
    .DIODE(la_oen_mprj[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__626__A (
    .DIODE(la_oen_mprj[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__627__A (
    .DIODE(la_oen_mprj[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__628__A (
    .DIODE(la_oen_mprj[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__629__A (
    .DIODE(la_oen_mprj[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__630__A (
    .DIODE(la_oen_mprj[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__631__A (
    .DIODE(la_oen_mprj[32]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__632__A (
    .DIODE(la_oen_mprj[33]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__633__A (
    .DIODE(la_oen_mprj[34]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__634__A (
    .DIODE(la_oen_mprj[35]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__635__A (
    .DIODE(la_oen_mprj[36]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__636__A (
    .DIODE(la_oen_mprj[37]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__637__A (
    .DIODE(la_oen_mprj[38]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__638__A (
    .DIODE(la_oen_mprj[39]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__639__A (
    .DIODE(la_oen_mprj[40]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__640__A (
    .DIODE(la_oen_mprj[41]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__641__A (
    .DIODE(la_oen_mprj[42]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__642__A (
    .DIODE(la_oen_mprj[43]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__643__A (
    .DIODE(la_oen_mprj[44]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__644__A (
    .DIODE(la_oen_mprj[45]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__645__A (
    .DIODE(la_oen_mprj[46]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__646__A (
    .DIODE(la_oen_mprj[47]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__647__A (
    .DIODE(la_oen_mprj[48]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__648__A (
    .DIODE(la_oen_mprj[49]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__649__A (
    .DIODE(la_oen_mprj[50]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__650__A (
    .DIODE(la_oen_mprj[51]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__651__A (
    .DIODE(la_oen_mprj[52]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__652__A (
    .DIODE(la_oen_mprj[53]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__653__A (
    .DIODE(la_oen_mprj[54]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__654__A (
    .DIODE(la_oen_mprj[55]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__655__A (
    .DIODE(la_oen_mprj[56]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__656__A (
    .DIODE(la_oen_mprj[57]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__657__A (
    .DIODE(la_oen_mprj[58]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__658__A (
    .DIODE(la_oen_mprj[59]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__659__A (
    .DIODE(la_oen_mprj[60]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA__660__A (
    .DIODE(la_oen_mprj[61]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[0]_A  (
    .DIODE(_074_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[0]_TE  (
    .DIODE(\mprj_logic1[74] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[100]_A  (
    .DIODE(_075_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[100]_TE  (
    .DIODE(\mprj_logic1[174] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[101]_A  (
    .DIODE(_076_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[101]_TE  (
    .DIODE(\mprj_logic1[175] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[102]_A  (
    .DIODE(_077_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[102]_TE  (
    .DIODE(\mprj_logic1[176] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[103]_A  (
    .DIODE(_078_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[103]_TE  (
    .DIODE(\mprj_logic1[177] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[104]_A  (
    .DIODE(_079_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[104]_TE  (
    .DIODE(\mprj_logic1[178] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[105]_A  (
    .DIODE(_080_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[105]_TE  (
    .DIODE(\mprj_logic1[179] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[106]_A  (
    .DIODE(_081_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[106]_TE  (
    .DIODE(\mprj_logic1[180] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[107]_A  (
    .DIODE(_082_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[107]_TE  (
    .DIODE(\mprj_logic1[181] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[108]_A  (
    .DIODE(_083_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[108]_TE  (
    .DIODE(\mprj_logic1[182] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[109]_A  (
    .DIODE(_084_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[109]_TE  (
    .DIODE(\mprj_logic1[183] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[10]_A  (
    .DIODE(_085_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[10]_TE  (
    .DIODE(\mprj_logic1[84] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[110]_A  (
    .DIODE(_086_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[110]_TE  (
    .DIODE(\mprj_logic1[184] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[111]_A  (
    .DIODE(_087_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[111]_TE  (
    .DIODE(\mprj_logic1[185] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[112]_A  (
    .DIODE(_088_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[112]_TE  (
    .DIODE(\mprj_logic1[186] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[113]_A  (
    .DIODE(_089_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[113]_TE  (
    .DIODE(\mprj_logic1[187] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[114]_A  (
    .DIODE(_090_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[114]_TE  (
    .DIODE(\mprj_logic1[188] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[115]_A  (
    .DIODE(_091_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[115]_TE  (
    .DIODE(\mprj_logic1[189] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[116]_A  (
    .DIODE(_092_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[116]_TE  (
    .DIODE(\mprj_logic1[190] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[117]_A  (
    .DIODE(_093_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[117]_TE  (
    .DIODE(\mprj_logic1[191] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[118]_A  (
    .DIODE(_094_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[118]_TE  (
    .DIODE(\mprj_logic1[192] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[119]_A  (
    .DIODE(_095_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[119]_TE  (
    .DIODE(\mprj_logic1[193] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[11]_A  (
    .DIODE(_096_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[11]_TE  (
    .DIODE(\mprj_logic1[85] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[120]_A  (
    .DIODE(_097_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[120]_TE  (
    .DIODE(\mprj_logic1[194] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[121]_A  (
    .DIODE(_098_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[121]_TE  (
    .DIODE(\mprj_logic1[195] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[122]_A  (
    .DIODE(_099_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[122]_TE  (
    .DIODE(\mprj_logic1[196] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[123]_A  (
    .DIODE(_100_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[123]_TE  (
    .DIODE(\mprj_logic1[197] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[124]_A  (
    .DIODE(_101_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[124]_TE  (
    .DIODE(\mprj_logic1[198] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[125]_A  (
    .DIODE(_102_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[125]_TE  (
    .DIODE(\mprj_logic1[199] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[126]_A  (
    .DIODE(_103_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[126]_TE  (
    .DIODE(\mprj_logic1[200] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[127]_A  (
    .DIODE(_104_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[127]_TE  (
    .DIODE(\mprj_logic1[201] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[12]_A  (
    .DIODE(_105_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[12]_TE  (
    .DIODE(\mprj_logic1[86] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[13]_A  (
    .DIODE(_106_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[13]_TE  (
    .DIODE(\mprj_logic1[87] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[14]_A  (
    .DIODE(_107_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[14]_TE  (
    .DIODE(\mprj_logic1[88] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[15]_A  (
    .DIODE(_108_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[15]_TE  (
    .DIODE(\mprj_logic1[89] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[16]_A  (
    .DIODE(_109_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[16]_TE  (
    .DIODE(\mprj_logic1[90] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[17]_A  (
    .DIODE(_110_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[17]_TE  (
    .DIODE(\mprj_logic1[91] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[18]_A  (
    .DIODE(_111_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[18]_TE  (
    .DIODE(\mprj_logic1[92] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[19]_A  (
    .DIODE(_112_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[19]_TE  (
    .DIODE(\mprj_logic1[93] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[1]_A  (
    .DIODE(_113_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[1]_TE  (
    .DIODE(\mprj_logic1[75] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[20]_A  (
    .DIODE(_114_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[20]_TE  (
    .DIODE(\mprj_logic1[94] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[21]_A  (
    .DIODE(_115_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[21]_TE  (
    .DIODE(\mprj_logic1[95] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[22]_A  (
    .DIODE(_116_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[22]_TE  (
    .DIODE(\mprj_logic1[96] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[23]_A  (
    .DIODE(_117_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[23]_TE  (
    .DIODE(\mprj_logic1[97] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[24]_A  (
    .DIODE(_118_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[24]_TE  (
    .DIODE(\mprj_logic1[98] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[25]_A  (
    .DIODE(_119_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[25]_TE  (
    .DIODE(\mprj_logic1[99] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[26]_A  (
    .DIODE(_120_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[26]_TE  (
    .DIODE(\mprj_logic1[100] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[27]_A  (
    .DIODE(_121_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[27]_TE  (
    .DIODE(\mprj_logic1[101] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[28]_A  (
    .DIODE(_122_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[28]_TE  (
    .DIODE(\mprj_logic1[102] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[29]_A  (
    .DIODE(_123_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[29]_TE  (
    .DIODE(\mprj_logic1[103] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[2]_A  (
    .DIODE(_124_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[2]_TE  (
    .DIODE(\mprj_logic1[76] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[30]_A  (
    .DIODE(_125_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[30]_TE  (
    .DIODE(\mprj_logic1[104] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[31]_A  (
    .DIODE(_126_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[31]_TE  (
    .DIODE(\mprj_logic1[105] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[32]_A  (
    .DIODE(_127_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[32]_TE  (
    .DIODE(\mprj_logic1[106] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[33]_A  (
    .DIODE(_128_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[33]_TE  (
    .DIODE(\mprj_logic1[107] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[34]_A  (
    .DIODE(_129_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[34]_TE  (
    .DIODE(\mprj_logic1[108] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[35]_A  (
    .DIODE(_130_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[35]_TE  (
    .DIODE(\mprj_logic1[109] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[36]_A  (
    .DIODE(_131_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[36]_TE  (
    .DIODE(\mprj_logic1[110] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[37]_A  (
    .DIODE(_132_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[37]_TE  (
    .DIODE(\mprj_logic1[111] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[38]_A  (
    .DIODE(_133_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[38]_TE  (
    .DIODE(\mprj_logic1[112] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[39]_A  (
    .DIODE(_134_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[39]_TE  (
    .DIODE(\mprj_logic1[113] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[3]_A  (
    .DIODE(_135_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[3]_TE  (
    .DIODE(\mprj_logic1[77] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[40]_A  (
    .DIODE(_136_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[40]_TE  (
    .DIODE(\mprj_logic1[114] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[41]_A  (
    .DIODE(_137_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[41]_TE  (
    .DIODE(\mprj_logic1[115] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[42]_A  (
    .DIODE(_138_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[42]_TE  (
    .DIODE(\mprj_logic1[116] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[43]_A  (
    .DIODE(_139_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[43]_TE  (
    .DIODE(\mprj_logic1[117] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[44]_A  (
    .DIODE(_140_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[44]_TE  (
    .DIODE(\mprj_logic1[118] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[45]_A  (
    .DIODE(_141_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[45]_TE  (
    .DIODE(\mprj_logic1[119] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[46]_A  (
    .DIODE(_142_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[46]_TE  (
    .DIODE(\mprj_logic1[120] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[47]_A  (
    .DIODE(_143_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[47]_TE  (
    .DIODE(\mprj_logic1[121] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[48]_A  (
    .DIODE(_144_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[48]_TE  (
    .DIODE(\mprj_logic1[122] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[49]_A  (
    .DIODE(_145_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[49]_TE  (
    .DIODE(\mprj_logic1[123] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[4]_A  (
    .DIODE(_146_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[4]_TE  (
    .DIODE(\mprj_logic1[78] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[50]_A  (
    .DIODE(_147_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[50]_TE  (
    .DIODE(\mprj_logic1[124] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[51]_A  (
    .DIODE(_148_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[51]_TE  (
    .DIODE(\mprj_logic1[125] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[52]_A  (
    .DIODE(_149_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[52]_TE  (
    .DIODE(\mprj_logic1[126] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[53]_A  (
    .DIODE(_150_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[53]_TE  (
    .DIODE(\mprj_logic1[127] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[54]_A  (
    .DIODE(_151_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[54]_TE  (
    .DIODE(\mprj_logic1[128] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[55]_A  (
    .DIODE(_152_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[55]_TE  (
    .DIODE(\mprj_logic1[129] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[56]_A  (
    .DIODE(_153_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[56]_TE  (
    .DIODE(\mprj_logic1[130] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[57]_A  (
    .DIODE(_154_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[57]_TE  (
    .DIODE(\mprj_logic1[131] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[58]_A  (
    .DIODE(_155_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[58]_TE  (
    .DIODE(\mprj_logic1[132] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[59]_A  (
    .DIODE(_156_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[59]_TE  (
    .DIODE(\mprj_logic1[133] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[5]_A  (
    .DIODE(_157_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[5]_TE  (
    .DIODE(\mprj_logic1[79] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[60]_A  (
    .DIODE(_158_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[60]_TE  (
    .DIODE(\mprj_logic1[134] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[61]_A  (
    .DIODE(_159_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[61]_TE  (
    .DIODE(\mprj_logic1[135] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[62]_A  (
    .DIODE(_160_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[62]_TE  (
    .DIODE(\mprj_logic1[136] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[63]_A  (
    .DIODE(_161_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[63]_TE  (
    .DIODE(\mprj_logic1[137] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[64]_A  (
    .DIODE(_162_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[64]_TE  (
    .DIODE(\mprj_logic1[138] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[65]_A  (
    .DIODE(_163_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[65]_TE  (
    .DIODE(\mprj_logic1[139] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[66]_A  (
    .DIODE(_164_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[66]_TE  (
    .DIODE(\mprj_logic1[140] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[67]_A  (
    .DIODE(_165_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[67]_TE  (
    .DIODE(\mprj_logic1[141] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[68]_A  (
    .DIODE(_166_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[68]_TE  (
    .DIODE(\mprj_logic1[142] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[69]_A  (
    .DIODE(_167_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[69]_TE  (
    .DIODE(\mprj_logic1[143] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[6]_A  (
    .DIODE(_168_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[6]_TE  (
    .DIODE(\mprj_logic1[80] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[70]_A  (
    .DIODE(_169_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[70]_TE  (
    .DIODE(\mprj_logic1[144] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[71]_A  (
    .DIODE(_170_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[71]_TE  (
    .DIODE(\mprj_logic1[145] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[72]_A  (
    .DIODE(_171_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[72]_TE  (
    .DIODE(\mprj_logic1[146] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[73]_A  (
    .DIODE(_172_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[73]_TE  (
    .DIODE(\mprj_logic1[147] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[74]_A  (
    .DIODE(_173_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[74]_TE  (
    .DIODE(\mprj_logic1[148] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[75]_A  (
    .DIODE(_174_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[75]_TE  (
    .DIODE(\mprj_logic1[149] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[76]_A  (
    .DIODE(_175_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[76]_TE  (
    .DIODE(\mprj_logic1[150] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[77]_A  (
    .DIODE(_176_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[77]_TE  (
    .DIODE(\mprj_logic1[151] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[78]_A  (
    .DIODE(_177_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[78]_TE  (
    .DIODE(\mprj_logic1[152] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[79]_A  (
    .DIODE(_178_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[79]_TE  (
    .DIODE(\mprj_logic1[153] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[7]_A  (
    .DIODE(_179_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[7]_TE  (
    .DIODE(\mprj_logic1[81] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[80]_A  (
    .DIODE(_180_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[80]_TE  (
    .DIODE(\mprj_logic1[154] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[81]_A  (
    .DIODE(_181_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[81]_TE  (
    .DIODE(\mprj_logic1[155] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[82]_A  (
    .DIODE(_182_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[82]_TE  (
    .DIODE(\mprj_logic1[156] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[83]_A  (
    .DIODE(_183_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[83]_TE  (
    .DIODE(\mprj_logic1[157] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[84]_A  (
    .DIODE(_184_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[84]_TE  (
    .DIODE(\mprj_logic1[158] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[85]_A  (
    .DIODE(_185_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[85]_TE  (
    .DIODE(\mprj_logic1[159] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[86]_A  (
    .DIODE(_186_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[86]_TE  (
    .DIODE(\mprj_logic1[160] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[87]_A  (
    .DIODE(_187_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[87]_TE  (
    .DIODE(\mprj_logic1[161] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[88]_A  (
    .DIODE(_188_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[88]_TE  (
    .DIODE(\mprj_logic1[162] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[89]_A  (
    .DIODE(_189_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[89]_TE  (
    .DIODE(\mprj_logic1[163] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[8]_A  (
    .DIODE(_190_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[8]_TE  (
    .DIODE(\mprj_logic1[82] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[90]_A  (
    .DIODE(_191_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[90]_TE  (
    .DIODE(\mprj_logic1[164] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[91]_A  (
    .DIODE(_192_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[91]_TE  (
    .DIODE(\mprj_logic1[165] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[92]_A  (
    .DIODE(_193_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[92]_TE  (
    .DIODE(\mprj_logic1[166] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[93]_A  (
    .DIODE(_194_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[93]_TE  (
    .DIODE(\mprj_logic1[167] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[94]_A  (
    .DIODE(_195_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[94]_TE  (
    .DIODE(\mprj_logic1[168] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[95]_A  (
    .DIODE(_196_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[95]_TE  (
    .DIODE(\mprj_logic1[169] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[96]_A  (
    .DIODE(_197_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[96]_TE  (
    .DIODE(\mprj_logic1[170] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[97]_A  (
    .DIODE(_198_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[97]_TE  (
    .DIODE(\mprj_logic1[171] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[98]_A  (
    .DIODE(_199_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[98]_TE  (
    .DIODE(\mprj_logic1[172] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[99]_A  (
    .DIODE(_200_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[99]_TE  (
    .DIODE(\mprj_logic1[173] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[9]_A  (
    .DIODE(_201_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_la_buf[9]_TE  (
    .DIODE(\mprj_logic1[83] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj2_pwrgood_A (
    .DIODE(mprj2_logic1),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj2_vdd_pwrgood_A (
    .DIODE(mprj2_vdd_logic1),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[0]_A  (
    .DIODE(_010_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[0]_TE  (
    .DIODE(\mprj_logic1[10] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[10]_A  (
    .DIODE(_011_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[10]_TE  (
    .DIODE(\mprj_logic1[20] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[11]_A  (
    .DIODE(_012_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[11]_TE  (
    .DIODE(\mprj_logic1[21] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[12]_A  (
    .DIODE(_013_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[12]_TE  (
    .DIODE(\mprj_logic1[22] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[13]_A  (
    .DIODE(_014_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[13]_TE  (
    .DIODE(\mprj_logic1[23] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[14]_A  (
    .DIODE(_015_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[14]_TE  (
    .DIODE(\mprj_logic1[24] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[15]_A  (
    .DIODE(_016_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[15]_TE  (
    .DIODE(\mprj_logic1[25] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[16]_A  (
    .DIODE(_017_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[16]_TE  (
    .DIODE(\mprj_logic1[26] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[17]_A  (
    .DIODE(_018_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[17]_TE  (
    .DIODE(\mprj_logic1[27] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[18]_A  (
    .DIODE(_019_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[18]_TE  (
    .DIODE(\mprj_logic1[28] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[19]_A  (
    .DIODE(_020_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[19]_TE  (
    .DIODE(\mprj_logic1[29] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[1]_A  (
    .DIODE(_021_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[1]_TE  (
    .DIODE(\mprj_logic1[11] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[20]_A  (
    .DIODE(_022_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[20]_TE  (
    .DIODE(\mprj_logic1[30] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[21]_A  (
    .DIODE(_023_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[21]_TE  (
    .DIODE(\mprj_logic1[31] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[22]_A  (
    .DIODE(_024_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[22]_TE  (
    .DIODE(\mprj_logic1[32] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[23]_A  (
    .DIODE(_025_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[23]_TE  (
    .DIODE(\mprj_logic1[33] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[24]_A  (
    .DIODE(_026_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[24]_TE  (
    .DIODE(\mprj_logic1[34] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[25]_A  (
    .DIODE(_027_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[25]_TE  (
    .DIODE(\mprj_logic1[35] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[26]_A  (
    .DIODE(_028_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[26]_TE  (
    .DIODE(\mprj_logic1[36] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[27]_A  (
    .DIODE(_029_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[27]_TE  (
    .DIODE(\mprj_logic1[37] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[28]_A  (
    .DIODE(_030_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[28]_TE  (
    .DIODE(\mprj_logic1[38] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[29]_A  (
    .DIODE(_031_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[29]_TE  (
    .DIODE(\mprj_logic1[39] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[2]_A  (
    .DIODE(_032_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[2]_TE  (
    .DIODE(\mprj_logic1[12] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[30]_A  (
    .DIODE(_033_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[30]_TE  (
    .DIODE(\mprj_logic1[40] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[31]_A  (
    .DIODE(_034_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[31]_TE  (
    .DIODE(\mprj_logic1[41] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[3]_A  (
    .DIODE(_035_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[3]_TE  (
    .DIODE(\mprj_logic1[13] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[4]_A  (
    .DIODE(_036_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[4]_TE  (
    .DIODE(\mprj_logic1[14] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[5]_A  (
    .DIODE(_037_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[5]_TE  (
    .DIODE(\mprj_logic1[15] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[6]_A  (
    .DIODE(_038_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[6]_TE  (
    .DIODE(\mprj_logic1[16] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[7]_A  (
    .DIODE(_039_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[7]_TE  (
    .DIODE(\mprj_logic1[17] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[8]_A  (
    .DIODE(_040_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[8]_TE  (
    .DIODE(\mprj_logic1[18] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[9]_A  (
    .DIODE(_041_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_adr_buf[9]_TE  (
    .DIODE(\mprj_logic1[19] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_clk2_buf_A (
    .DIODE(_002_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_clk2_buf_TE (
    .DIODE(\mprj_logic1[2] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_clk_buf_A (
    .DIODE(_001_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_clk_buf_TE (
    .DIODE(\mprj_logic1[1] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_cyc_buf_A (
    .DIODE(_003_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_cyc_buf_TE (
    .DIODE(\mprj_logic1[3] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[0]_A  (
    .DIODE(_042_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[0]_TE  (
    .DIODE(\mprj_logic1[42] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[10]_A  (
    .DIODE(_043_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[10]_TE  (
    .DIODE(\mprj_logic1[52] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[11]_A  (
    .DIODE(_044_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[11]_TE  (
    .DIODE(\mprj_logic1[53] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[12]_A  (
    .DIODE(_045_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[12]_TE  (
    .DIODE(\mprj_logic1[54] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[13]_A  (
    .DIODE(_046_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[13]_TE  (
    .DIODE(\mprj_logic1[55] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[14]_A  (
    .DIODE(_047_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[14]_TE  (
    .DIODE(\mprj_logic1[56] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[15]_A  (
    .DIODE(_048_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[15]_TE  (
    .DIODE(\mprj_logic1[57] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[16]_A  (
    .DIODE(_049_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[16]_TE  (
    .DIODE(\mprj_logic1[58] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[17]_A  (
    .DIODE(_050_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[17]_TE  (
    .DIODE(\mprj_logic1[59] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[18]_A  (
    .DIODE(_051_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[18]_TE  (
    .DIODE(\mprj_logic1[60] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[19]_A  (
    .DIODE(_052_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[19]_TE  (
    .DIODE(\mprj_logic1[61] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[1]_A  (
    .DIODE(_053_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[1]_TE  (
    .DIODE(\mprj_logic1[43] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[20]_A  (
    .DIODE(_054_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[20]_TE  (
    .DIODE(\mprj_logic1[62] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[21]_A  (
    .DIODE(_055_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[21]_TE  (
    .DIODE(\mprj_logic1[63] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[22]_A  (
    .DIODE(_056_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[22]_TE  (
    .DIODE(\mprj_logic1[64] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[23]_A  (
    .DIODE(_057_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[23]_TE  (
    .DIODE(\mprj_logic1[65] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[24]_A  (
    .DIODE(_058_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[24]_TE  (
    .DIODE(\mprj_logic1[66] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[25]_A  (
    .DIODE(_059_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[25]_TE  (
    .DIODE(\mprj_logic1[67] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[26]_A  (
    .DIODE(_060_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[26]_TE  (
    .DIODE(\mprj_logic1[68] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[27]_A  (
    .DIODE(_061_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[27]_TE  (
    .DIODE(\mprj_logic1[69] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[28]_A  (
    .DIODE(_062_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[28]_TE  (
    .DIODE(\mprj_logic1[70] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[29]_A  (
    .DIODE(_063_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[29]_TE  (
    .DIODE(\mprj_logic1[71] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[2]_A  (
    .DIODE(_064_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[2]_TE  (
    .DIODE(\mprj_logic1[44] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[30]_A  (
    .DIODE(_065_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[30]_TE  (
    .DIODE(\mprj_logic1[72] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[31]_A  (
    .DIODE(_066_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[31]_TE  (
    .DIODE(\mprj_logic1[73] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[3]_A  (
    .DIODE(_067_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[3]_TE  (
    .DIODE(\mprj_logic1[45] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[4]_A  (
    .DIODE(_068_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[4]_TE  (
    .DIODE(\mprj_logic1[46] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[5]_A  (
    .DIODE(_069_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[5]_TE  (
    .DIODE(\mprj_logic1[47] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[6]_A  (
    .DIODE(_070_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[6]_TE  (
    .DIODE(\mprj_logic1[48] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[7]_A  (
    .DIODE(_071_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[7]_TE  (
    .DIODE(\mprj_logic1[49] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[8]_A  (
    .DIODE(_072_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[8]_TE  (
    .DIODE(\mprj_logic1[50] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[9]_A  (
    .DIODE(_073_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_dat_buf[9]_TE  (
    .DIODE(\mprj_logic1[51] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_pwrgood_A (
    .DIODE(\mprj_logic1[458] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_rstn_buf_A (
    .DIODE(_000_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_rstn_buf_TE (
    .DIODE(\mprj_logic1[0] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[0]_A  (
    .DIODE(_006_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[0]_TE  (
    .DIODE(\mprj_logic1[6] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[1]_A  (
    .DIODE(_007_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[1]_TE  (
    .DIODE(\mprj_logic1[7] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[2]_A  (
    .DIODE(_008_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[2]_TE  (
    .DIODE(\mprj_logic1[8] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[3]_A  (
    .DIODE(_009_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_mprj_sel_buf[3]_TE  (
    .DIODE(\mprj_logic1[9] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_stb_buf_A (
    .DIODE(_004_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_stb_buf_TE (
    .DIODE(\mprj_logic1[4] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_vdd_pwrgood_A (
    .DIODE(mprj_vdd_logic1),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_we_buf_A (
    .DIODE(_005_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_mprj_we_buf_TE (
    .DIODE(\mprj_logic1[5] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[0]_A  (
    .DIODE(\la_data_in_mprj_bar[0] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[100]_A  (
    .DIODE(\la_data_in_mprj_bar[100] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[101]_A  (
    .DIODE(\la_data_in_mprj_bar[101] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[102]_A  (
    .DIODE(\la_data_in_mprj_bar[102] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[103]_A  (
    .DIODE(\la_data_in_mprj_bar[103] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[104]_A  (
    .DIODE(\la_data_in_mprj_bar[104] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[105]_A  (
    .DIODE(\la_data_in_mprj_bar[105] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[106]_A  (
    .DIODE(\la_data_in_mprj_bar[106] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[107]_A  (
    .DIODE(\la_data_in_mprj_bar[107] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[108]_A  (
    .DIODE(\la_data_in_mprj_bar[108] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[109]_A  (
    .DIODE(\la_data_in_mprj_bar[109] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[10]_A  (
    .DIODE(\la_data_in_mprj_bar[10] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[110]_A  (
    .DIODE(\la_data_in_mprj_bar[110] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[111]_A  (
    .DIODE(\la_data_in_mprj_bar[111] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[112]_A  (
    .DIODE(\la_data_in_mprj_bar[112] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[113]_A  (
    .DIODE(\la_data_in_mprj_bar[113] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[114]_A  (
    .DIODE(\la_data_in_mprj_bar[114] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[115]_A  (
    .DIODE(\la_data_in_mprj_bar[115] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[116]_A  (
    .DIODE(\la_data_in_mprj_bar[116] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[117]_A  (
    .DIODE(\la_data_in_mprj_bar[117] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[118]_A  (
    .DIODE(\la_data_in_mprj_bar[118] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[119]_A  (
    .DIODE(\la_data_in_mprj_bar[119] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[11]_A  (
    .DIODE(\la_data_in_mprj_bar[11] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[120]_A  (
    .DIODE(\la_data_in_mprj_bar[120] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[121]_A  (
    .DIODE(\la_data_in_mprj_bar[121] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[122]_A  (
    .DIODE(\la_data_in_mprj_bar[122] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[123]_A  (
    .DIODE(\la_data_in_mprj_bar[123] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[124]_A  (
    .DIODE(\la_data_in_mprj_bar[124] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[125]_A  (
    .DIODE(\la_data_in_mprj_bar[125] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[126]_A  (
    .DIODE(\la_data_in_mprj_bar[126] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[127]_A  (
    .DIODE(\la_data_in_mprj_bar[127] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[12]_A  (
    .DIODE(\la_data_in_mprj_bar[12] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[13]_A  (
    .DIODE(\la_data_in_mprj_bar[13] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[14]_A  (
    .DIODE(\la_data_in_mprj_bar[14] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[15]_A  (
    .DIODE(\la_data_in_mprj_bar[15] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[16]_A  (
    .DIODE(\la_data_in_mprj_bar[16] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[17]_A  (
    .DIODE(\la_data_in_mprj_bar[17] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[18]_A  (
    .DIODE(\la_data_in_mprj_bar[18] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[19]_A  (
    .DIODE(\la_data_in_mprj_bar[19] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[1]_A  (
    .DIODE(\la_data_in_mprj_bar[1] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[20]_A  (
    .DIODE(\la_data_in_mprj_bar[20] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[21]_A  (
    .DIODE(\la_data_in_mprj_bar[21] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[22]_A  (
    .DIODE(\la_data_in_mprj_bar[22] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[23]_A  (
    .DIODE(\la_data_in_mprj_bar[23] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[24]_A  (
    .DIODE(\la_data_in_mprj_bar[24] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[25]_A  (
    .DIODE(\la_data_in_mprj_bar[25] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[26]_A  (
    .DIODE(\la_data_in_mprj_bar[26] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[27]_A  (
    .DIODE(\la_data_in_mprj_bar[27] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[28]_A  (
    .DIODE(\la_data_in_mprj_bar[28] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[29]_A  (
    .DIODE(\la_data_in_mprj_bar[29] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[2]_A  (
    .DIODE(\la_data_in_mprj_bar[2] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[30]_A  (
    .DIODE(\la_data_in_mprj_bar[30] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[31]_A  (
    .DIODE(\la_data_in_mprj_bar[31] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[32]_A  (
    .DIODE(\la_data_in_mprj_bar[32] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[33]_A  (
    .DIODE(\la_data_in_mprj_bar[33] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[34]_A  (
    .DIODE(\la_data_in_mprj_bar[34] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[35]_A  (
    .DIODE(\la_data_in_mprj_bar[35] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[36]_A  (
    .DIODE(\la_data_in_mprj_bar[36] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[37]_A  (
    .DIODE(\la_data_in_mprj_bar[37] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[38]_A  (
    .DIODE(\la_data_in_mprj_bar[38] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[39]_A  (
    .DIODE(\la_data_in_mprj_bar[39] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[3]_A  (
    .DIODE(\la_data_in_mprj_bar[3] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[40]_A  (
    .DIODE(\la_data_in_mprj_bar[40] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[41]_A  (
    .DIODE(\la_data_in_mprj_bar[41] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[42]_A  (
    .DIODE(\la_data_in_mprj_bar[42] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[43]_A  (
    .DIODE(\la_data_in_mprj_bar[43] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[44]_A  (
    .DIODE(\la_data_in_mprj_bar[44] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[45]_A  (
    .DIODE(\la_data_in_mprj_bar[45] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[46]_A  (
    .DIODE(\la_data_in_mprj_bar[46] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[47]_A  (
    .DIODE(\la_data_in_mprj_bar[47] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[48]_A  (
    .DIODE(\la_data_in_mprj_bar[48] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[49]_A  (
    .DIODE(\la_data_in_mprj_bar[49] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[4]_A  (
    .DIODE(\la_data_in_mprj_bar[4] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[50]_A  (
    .DIODE(\la_data_in_mprj_bar[50] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[51]_A  (
    .DIODE(\la_data_in_mprj_bar[51] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[52]_A  (
    .DIODE(\la_data_in_mprj_bar[52] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[53]_A  (
    .DIODE(\la_data_in_mprj_bar[53] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[54]_A  (
    .DIODE(\la_data_in_mprj_bar[54] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[55]_A  (
    .DIODE(\la_data_in_mprj_bar[55] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[56]_A  (
    .DIODE(\la_data_in_mprj_bar[56] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[57]_A  (
    .DIODE(\la_data_in_mprj_bar[57] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[58]_A  (
    .DIODE(\la_data_in_mprj_bar[58] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[59]_A  (
    .DIODE(\la_data_in_mprj_bar[59] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[5]_A  (
    .DIODE(\la_data_in_mprj_bar[5] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[60]_A  (
    .DIODE(\la_data_in_mprj_bar[60] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[61]_A  (
    .DIODE(\la_data_in_mprj_bar[61] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[62]_A  (
    .DIODE(\la_data_in_mprj_bar[62] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[63]_A  (
    .DIODE(\la_data_in_mprj_bar[63] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[64]_A  (
    .DIODE(\la_data_in_mprj_bar[64] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[65]_A  (
    .DIODE(\la_data_in_mprj_bar[65] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[66]_A  (
    .DIODE(\la_data_in_mprj_bar[66] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[67]_A  (
    .DIODE(\la_data_in_mprj_bar[67] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[68]_A  (
    .DIODE(\la_data_in_mprj_bar[68] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[69]_A  (
    .DIODE(\la_data_in_mprj_bar[69] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[6]_A  (
    .DIODE(\la_data_in_mprj_bar[6] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[70]_A  (
    .DIODE(\la_data_in_mprj_bar[70] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[71]_A  (
    .DIODE(\la_data_in_mprj_bar[71] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[72]_A  (
    .DIODE(\la_data_in_mprj_bar[72] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[73]_A  (
    .DIODE(\la_data_in_mprj_bar[73] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[74]_A  (
    .DIODE(\la_data_in_mprj_bar[74] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[75]_A  (
    .DIODE(\la_data_in_mprj_bar[75] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[76]_A  (
    .DIODE(\la_data_in_mprj_bar[76] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[77]_A  (
    .DIODE(\la_data_in_mprj_bar[77] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[78]_A  (
    .DIODE(\la_data_in_mprj_bar[78] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[79]_A  (
    .DIODE(\la_data_in_mprj_bar[79] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[7]_A  (
    .DIODE(\la_data_in_mprj_bar[7] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[80]_A  (
    .DIODE(\la_data_in_mprj_bar[80] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[81]_A  (
    .DIODE(\la_data_in_mprj_bar[81] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[82]_A  (
    .DIODE(\la_data_in_mprj_bar[82] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[83]_A  (
    .DIODE(\la_data_in_mprj_bar[83] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[84]_A  (
    .DIODE(\la_data_in_mprj_bar[84] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[85]_A  (
    .DIODE(\la_data_in_mprj_bar[85] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[86]_A  (
    .DIODE(\la_data_in_mprj_bar[86] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[87]_A  (
    .DIODE(\la_data_in_mprj_bar[87] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[88]_A  (
    .DIODE(\la_data_in_mprj_bar[88] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[89]_A  (
    .DIODE(\la_data_in_mprj_bar[89] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[8]_A  (
    .DIODE(\la_data_in_mprj_bar[8] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[90]_A  (
    .DIODE(\la_data_in_mprj_bar[90] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[91]_A  (
    .DIODE(\la_data_in_mprj_bar[91] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[92]_A  (
    .DIODE(\la_data_in_mprj_bar[92] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[93]_A  (
    .DIODE(\la_data_in_mprj_bar[93] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[94]_A  (
    .DIODE(\la_data_in_mprj_bar[94] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[95]_A  (
    .DIODE(\la_data_in_mprj_bar[95] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[96]_A  (
    .DIODE(\la_data_in_mprj_bar[96] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[97]_A  (
    .DIODE(\la_data_in_mprj_bar[97] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[98]_A  (
    .DIODE(\la_data_in_mprj_bar[98] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[99]_A  (
    .DIODE(\la_data_in_mprj_bar[99] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_buffers[9]_A  (
    .DIODE(\la_data_in_mprj_bar[9] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[0]_A  (
    .DIODE(la_data_out_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[0]_B  (
    .DIODE(\mprj_logic1[330] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[100]_A  (
    .DIODE(la_data_out_core[100]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[100]_B  (
    .DIODE(\mprj_logic1[430] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[101]_A  (
    .DIODE(la_data_out_core[101]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[101]_B  (
    .DIODE(\mprj_logic1[431] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[102]_A  (
    .DIODE(la_data_out_core[102]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[102]_B  (
    .DIODE(\mprj_logic1[432] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[103]_A  (
    .DIODE(la_data_out_core[103]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[103]_B  (
    .DIODE(\mprj_logic1[433] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[104]_A  (
    .DIODE(la_data_out_core[104]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[104]_B  (
    .DIODE(\mprj_logic1[434] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[105]_A  (
    .DIODE(la_data_out_core[105]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[105]_B  (
    .DIODE(\mprj_logic1[435] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[106]_A  (
    .DIODE(la_data_out_core[106]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[106]_B  (
    .DIODE(\mprj_logic1[436] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[107]_A  (
    .DIODE(la_data_out_core[107]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[107]_B  (
    .DIODE(\mprj_logic1[437] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[108]_A  (
    .DIODE(la_data_out_core[108]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[108]_B  (
    .DIODE(\mprj_logic1[438] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[109]_A  (
    .DIODE(la_data_out_core[109]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[109]_B  (
    .DIODE(\mprj_logic1[439] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[10]_A  (
    .DIODE(la_data_out_core[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[10]_B  (
    .DIODE(\mprj_logic1[340] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[110]_A  (
    .DIODE(la_data_out_core[110]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[110]_B  (
    .DIODE(\mprj_logic1[440] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[111]_A  (
    .DIODE(la_data_out_core[111]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[111]_B  (
    .DIODE(\mprj_logic1[441] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[112]_A  (
    .DIODE(la_data_out_core[112]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[112]_B  (
    .DIODE(\mprj_logic1[442] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[113]_A  (
    .DIODE(la_data_out_core[113]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[113]_B  (
    .DIODE(\mprj_logic1[443] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[114]_A  (
    .DIODE(la_data_out_core[114]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[114]_B  (
    .DIODE(\mprj_logic1[444] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[115]_A  (
    .DIODE(la_data_out_core[115]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[115]_B  (
    .DIODE(\mprj_logic1[445] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[116]_A  (
    .DIODE(la_data_out_core[116]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[116]_B  (
    .DIODE(\mprj_logic1[446] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[117]_A  (
    .DIODE(la_data_out_core[117]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[117]_B  (
    .DIODE(\mprj_logic1[447] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[118]_A  (
    .DIODE(la_data_out_core[118]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[118]_B  (
    .DIODE(\mprj_logic1[448] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[119]_A  (
    .DIODE(la_data_out_core[119]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[119]_B  (
    .DIODE(\mprj_logic1[449] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[11]_A  (
    .DIODE(la_data_out_core[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[11]_B  (
    .DIODE(\mprj_logic1[341] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[120]_A  (
    .DIODE(la_data_out_core[120]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[120]_B  (
    .DIODE(\mprj_logic1[450] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[121]_A  (
    .DIODE(la_data_out_core[121]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[121]_B  (
    .DIODE(\mprj_logic1[451] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[122]_A  (
    .DIODE(la_data_out_core[122]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[122]_B  (
    .DIODE(\mprj_logic1[452] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[123]_A  (
    .DIODE(la_data_out_core[123]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[123]_B  (
    .DIODE(\mprj_logic1[453] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[124]_A  (
    .DIODE(la_data_out_core[124]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[124]_B  (
    .DIODE(\mprj_logic1[454] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[125]_A  (
    .DIODE(la_data_out_core[125]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[125]_B  (
    .DIODE(\mprj_logic1[455] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[126]_A  (
    .DIODE(la_data_out_core[126]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[126]_B  (
    .DIODE(\mprj_logic1[456] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[127]_A  (
    .DIODE(la_data_out_core[127]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[127]_B  (
    .DIODE(\mprj_logic1[457] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[12]_A  (
    .DIODE(la_data_out_core[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[12]_B  (
    .DIODE(\mprj_logic1[342] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[13]_A  (
    .DIODE(la_data_out_core[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[13]_B  (
    .DIODE(\mprj_logic1[343] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[14]_A  (
    .DIODE(la_data_out_core[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[14]_B  (
    .DIODE(\mprj_logic1[344] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[15]_A  (
    .DIODE(la_data_out_core[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[15]_B  (
    .DIODE(\mprj_logic1[345] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[16]_A  (
    .DIODE(la_data_out_core[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[16]_B  (
    .DIODE(\mprj_logic1[346] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[17]_A  (
    .DIODE(la_data_out_core[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[17]_B  (
    .DIODE(\mprj_logic1[347] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[18]_A  (
    .DIODE(la_data_out_core[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[18]_B  (
    .DIODE(\mprj_logic1[348] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[19]_A  (
    .DIODE(la_data_out_core[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[19]_B  (
    .DIODE(\mprj_logic1[349] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[1]_A  (
    .DIODE(la_data_out_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[1]_B  (
    .DIODE(\mprj_logic1[331] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[20]_A  (
    .DIODE(la_data_out_core[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[20]_B  (
    .DIODE(\mprj_logic1[350] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[21]_A  (
    .DIODE(la_data_out_core[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[21]_B  (
    .DIODE(\mprj_logic1[351] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[22]_A  (
    .DIODE(la_data_out_core[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[22]_B  (
    .DIODE(\mprj_logic1[352] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[23]_A  (
    .DIODE(la_data_out_core[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[23]_B  (
    .DIODE(\mprj_logic1[353] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[24]_A  (
    .DIODE(la_data_out_core[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[24]_B  (
    .DIODE(\mprj_logic1[354] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[25]_A  (
    .DIODE(la_data_out_core[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[25]_B  (
    .DIODE(\mprj_logic1[355] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[26]_A  (
    .DIODE(la_data_out_core[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[26]_B  (
    .DIODE(\mprj_logic1[356] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[27]_A  (
    .DIODE(la_data_out_core[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[27]_B  (
    .DIODE(\mprj_logic1[357] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[28]_A  (
    .DIODE(la_data_out_core[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[28]_B  (
    .DIODE(\mprj_logic1[358] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[29]_A  (
    .DIODE(la_data_out_core[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[29]_B  (
    .DIODE(\mprj_logic1[359] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[2]_A  (
    .DIODE(la_data_out_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[2]_B  (
    .DIODE(\mprj_logic1[332] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[30]_A  (
    .DIODE(la_data_out_core[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[30]_B  (
    .DIODE(\mprj_logic1[360] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[31]_A  (
    .DIODE(la_data_out_core[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[31]_B  (
    .DIODE(\mprj_logic1[361] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[32]_A  (
    .DIODE(la_data_out_core[32]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[32]_B  (
    .DIODE(\mprj_logic1[362] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[33]_A  (
    .DIODE(la_data_out_core[33]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[33]_B  (
    .DIODE(\mprj_logic1[363] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[34]_A  (
    .DIODE(la_data_out_core[34]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[34]_B  (
    .DIODE(\mprj_logic1[364] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[35]_A  (
    .DIODE(la_data_out_core[35]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[35]_B  (
    .DIODE(\mprj_logic1[365] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[36]_A  (
    .DIODE(la_data_out_core[36]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[36]_B  (
    .DIODE(\mprj_logic1[366] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[37]_A  (
    .DIODE(la_data_out_core[37]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[37]_B  (
    .DIODE(\mprj_logic1[367] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[38]_A  (
    .DIODE(la_data_out_core[38]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[38]_B  (
    .DIODE(\mprj_logic1[368] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[39]_A  (
    .DIODE(la_data_out_core[39]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[39]_B  (
    .DIODE(\mprj_logic1[369] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[3]_A  (
    .DIODE(la_data_out_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[3]_B  (
    .DIODE(\mprj_logic1[333] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[40]_A  (
    .DIODE(la_data_out_core[40]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[40]_B  (
    .DIODE(\mprj_logic1[370] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[41]_A  (
    .DIODE(la_data_out_core[41]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[41]_B  (
    .DIODE(\mprj_logic1[371] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[42]_A  (
    .DIODE(la_data_out_core[42]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[42]_B  (
    .DIODE(\mprj_logic1[372] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[43]_A  (
    .DIODE(la_data_out_core[43]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[43]_B  (
    .DIODE(\mprj_logic1[373] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[44]_A  (
    .DIODE(la_data_out_core[44]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[44]_B  (
    .DIODE(\mprj_logic1[374] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[45]_A  (
    .DIODE(la_data_out_core[45]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[45]_B  (
    .DIODE(\mprj_logic1[375] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[46]_A  (
    .DIODE(la_data_out_core[46]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[46]_B  (
    .DIODE(\mprj_logic1[376] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[47]_A  (
    .DIODE(la_data_out_core[47]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[47]_B  (
    .DIODE(\mprj_logic1[377] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[48]_A  (
    .DIODE(la_data_out_core[48]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[48]_B  (
    .DIODE(\mprj_logic1[378] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[49]_A  (
    .DIODE(la_data_out_core[49]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[49]_B  (
    .DIODE(\mprj_logic1[379] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[4]_A  (
    .DIODE(la_data_out_core[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[4]_B  (
    .DIODE(\mprj_logic1[334] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[50]_A  (
    .DIODE(la_data_out_core[50]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[50]_B  (
    .DIODE(\mprj_logic1[380] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[51]_A  (
    .DIODE(la_data_out_core[51]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[51]_B  (
    .DIODE(\mprj_logic1[381] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[52]_A  (
    .DIODE(la_data_out_core[52]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[52]_B  (
    .DIODE(\mprj_logic1[382] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[53]_A  (
    .DIODE(la_data_out_core[53]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[53]_B  (
    .DIODE(\mprj_logic1[383] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[54]_A  (
    .DIODE(la_data_out_core[54]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[54]_B  (
    .DIODE(\mprj_logic1[384] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[55]_A  (
    .DIODE(la_data_out_core[55]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[55]_B  (
    .DIODE(\mprj_logic1[385] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[56]_A  (
    .DIODE(la_data_out_core[56]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[56]_B  (
    .DIODE(\mprj_logic1[386] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[57]_A  (
    .DIODE(la_data_out_core[57]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[57]_B  (
    .DIODE(\mprj_logic1[387] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[58]_A  (
    .DIODE(la_data_out_core[58]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[58]_B  (
    .DIODE(\mprj_logic1[388] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[59]_A  (
    .DIODE(la_data_out_core[59]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[59]_B  (
    .DIODE(\mprj_logic1[389] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[5]_A  (
    .DIODE(la_data_out_core[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[5]_B  (
    .DIODE(\mprj_logic1[335] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[60]_A  (
    .DIODE(la_data_out_core[60]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[60]_B  (
    .DIODE(\mprj_logic1[390] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[61]_A  (
    .DIODE(la_data_out_core[61]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[61]_B  (
    .DIODE(\mprj_logic1[391] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[62]_A  (
    .DIODE(la_data_out_core[62]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[62]_B  (
    .DIODE(\mprj_logic1[392] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[63]_A  (
    .DIODE(la_data_out_core[63]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[63]_B  (
    .DIODE(\mprj_logic1[393] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[64]_A  (
    .DIODE(la_data_out_core[64]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[64]_B  (
    .DIODE(\mprj_logic1[394] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[65]_A  (
    .DIODE(la_data_out_core[65]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[65]_B  (
    .DIODE(\mprj_logic1[395] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[66]_A  (
    .DIODE(la_data_out_core[66]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[66]_B  (
    .DIODE(\mprj_logic1[396] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[67]_A  (
    .DIODE(la_data_out_core[67]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[67]_B  (
    .DIODE(\mprj_logic1[397] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[68]_A  (
    .DIODE(la_data_out_core[68]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[68]_B  (
    .DIODE(\mprj_logic1[398] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[69]_A  (
    .DIODE(la_data_out_core[69]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[69]_B  (
    .DIODE(\mprj_logic1[399] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[6]_A  (
    .DIODE(la_data_out_core[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[6]_B  (
    .DIODE(\mprj_logic1[336] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[70]_A  (
    .DIODE(la_data_out_core[70]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[70]_B  (
    .DIODE(\mprj_logic1[400] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[71]_A  (
    .DIODE(la_data_out_core[71]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[71]_B  (
    .DIODE(\mprj_logic1[401] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[72]_A  (
    .DIODE(la_data_out_core[72]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[72]_B  (
    .DIODE(\mprj_logic1[402] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[73]_A  (
    .DIODE(la_data_out_core[73]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[73]_B  (
    .DIODE(\mprj_logic1[403] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[74]_A  (
    .DIODE(la_data_out_core[74]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[74]_B  (
    .DIODE(\mprj_logic1[404] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[75]_A  (
    .DIODE(la_data_out_core[75]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[75]_B  (
    .DIODE(\mprj_logic1[405] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[76]_A  (
    .DIODE(la_data_out_core[76]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[76]_B  (
    .DIODE(\mprj_logic1[406] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[77]_A  (
    .DIODE(la_data_out_core[77]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[77]_B  (
    .DIODE(\mprj_logic1[407] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[78]_A  (
    .DIODE(la_data_out_core[78]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[78]_B  (
    .DIODE(\mprj_logic1[408] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[79]_A  (
    .DIODE(la_data_out_core[79]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[79]_B  (
    .DIODE(\mprj_logic1[409] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[7]_A  (
    .DIODE(la_data_out_core[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[7]_B  (
    .DIODE(\mprj_logic1[337] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[80]_A  (
    .DIODE(la_data_out_core[80]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[80]_B  (
    .DIODE(\mprj_logic1[410] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[81]_A  (
    .DIODE(la_data_out_core[81]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[81]_B  (
    .DIODE(\mprj_logic1[411] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[82]_A  (
    .DIODE(la_data_out_core[82]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[82]_B  (
    .DIODE(\mprj_logic1[412] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[83]_A  (
    .DIODE(la_data_out_core[83]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[83]_B  (
    .DIODE(\mprj_logic1[413] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[84]_A  (
    .DIODE(la_data_out_core[84]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[84]_B  (
    .DIODE(\mprj_logic1[414] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[85]_A  (
    .DIODE(la_data_out_core[85]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[85]_B  (
    .DIODE(\mprj_logic1[415] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[86]_A  (
    .DIODE(la_data_out_core[86]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[86]_B  (
    .DIODE(\mprj_logic1[416] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[87]_A  (
    .DIODE(la_data_out_core[87]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[87]_B  (
    .DIODE(\mprj_logic1[417] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[88]_A  (
    .DIODE(la_data_out_core[88]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[88]_B  (
    .DIODE(\mprj_logic1[418] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[89]_A  (
    .DIODE(la_data_out_core[89]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[89]_B  (
    .DIODE(\mprj_logic1[419] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[8]_A  (
    .DIODE(la_data_out_core[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[8]_B  (
    .DIODE(\mprj_logic1[338] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[90]_A  (
    .DIODE(la_data_out_core[90]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[90]_B  (
    .DIODE(\mprj_logic1[420] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[91]_A  (
    .DIODE(la_data_out_core[91]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[91]_B  (
    .DIODE(\mprj_logic1[421] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[92]_A  (
    .DIODE(la_data_out_core[92]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[92]_B  (
    .DIODE(\mprj_logic1[422] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[93]_A  (
    .DIODE(la_data_out_core[93]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[93]_B  (
    .DIODE(\mprj_logic1[423] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[94]_A  (
    .DIODE(la_data_out_core[94]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[94]_B  (
    .DIODE(\mprj_logic1[424] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[95]_A  (
    .DIODE(la_data_out_core[95]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[95]_B  (
    .DIODE(\mprj_logic1[425] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[96]_A  (
    .DIODE(la_data_out_core[96]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[96]_B  (
    .DIODE(\mprj_logic1[426] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[97]_A  (
    .DIODE(la_data_out_core[97]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[97]_B  (
    .DIODE(\mprj_logic1[427] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[98]_A  (
    .DIODE(la_data_out_core[98]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[98]_B  (
    .DIODE(\mprj_logic1[428] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[99]_A  (
    .DIODE(la_data_out_core[99]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[99]_B  (
    .DIODE(\mprj_logic1[429] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[9]_A  (
    .DIODE(la_data_out_core[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[9]_B  (
    .DIODE(\mprj_logic1[339] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[0]_A  (
    .DIODE(_202_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[0]_TE  (
    .DIODE(\mprj_logic1[202] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[100]_A  (
    .DIODE(_203_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[100]_TE  (
    .DIODE(\mprj_logic1[302] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[101]_A  (
    .DIODE(_204_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[101]_TE  (
    .DIODE(\mprj_logic1[303] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[102]_A  (
    .DIODE(_205_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[102]_TE  (
    .DIODE(\mprj_logic1[304] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[103]_A  (
    .DIODE(_206_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[103]_TE  (
    .DIODE(\mprj_logic1[305] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[104]_A  (
    .DIODE(_207_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[104]_TE  (
    .DIODE(\mprj_logic1[306] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[105]_A  (
    .DIODE(_208_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[105]_TE  (
    .DIODE(\mprj_logic1[307] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[106]_A  (
    .DIODE(_209_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[106]_TE  (
    .DIODE(\mprj_logic1[308] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[107]_A  (
    .DIODE(_210_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[107]_TE  (
    .DIODE(\mprj_logic1[309] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[108]_A  (
    .DIODE(_211_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[108]_TE  (
    .DIODE(\mprj_logic1[310] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[109]_A  (
    .DIODE(_212_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[109]_TE  (
    .DIODE(\mprj_logic1[311] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[10]_A  (
    .DIODE(_213_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[10]_TE  (
    .DIODE(\mprj_logic1[212] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[110]_A  (
    .DIODE(_214_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[110]_TE  (
    .DIODE(\mprj_logic1[312] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[111]_A  (
    .DIODE(_215_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[111]_TE  (
    .DIODE(\mprj_logic1[313] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[112]_A  (
    .DIODE(_216_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[112]_TE  (
    .DIODE(\mprj_logic1[314] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[113]_A  (
    .DIODE(_217_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[113]_TE  (
    .DIODE(\mprj_logic1[315] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[114]_A  (
    .DIODE(_218_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[114]_TE  (
    .DIODE(\mprj_logic1[316] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[115]_A  (
    .DIODE(_219_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[115]_TE  (
    .DIODE(\mprj_logic1[317] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[116]_A  (
    .DIODE(_220_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[116]_TE  (
    .DIODE(\mprj_logic1[318] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[117]_A  (
    .DIODE(_221_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[117]_TE  (
    .DIODE(\mprj_logic1[319] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[118]_A  (
    .DIODE(_222_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[118]_TE  (
    .DIODE(\mprj_logic1[320] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[119]_A  (
    .DIODE(_223_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[119]_TE  (
    .DIODE(\mprj_logic1[321] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[11]_A  (
    .DIODE(_224_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[11]_TE  (
    .DIODE(\mprj_logic1[213] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[120]_A  (
    .DIODE(_225_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[120]_TE  (
    .DIODE(\mprj_logic1[322] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[121]_A  (
    .DIODE(_226_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[121]_TE  (
    .DIODE(\mprj_logic1[323] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[122]_A  (
    .DIODE(_227_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[122]_TE  (
    .DIODE(\mprj_logic1[324] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[123]_A  (
    .DIODE(_228_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[123]_TE  (
    .DIODE(\mprj_logic1[325] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[124]_A  (
    .DIODE(_229_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[124]_TE  (
    .DIODE(\mprj_logic1[326] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[125]_A  (
    .DIODE(_230_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[125]_TE  (
    .DIODE(\mprj_logic1[327] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[126]_A  (
    .DIODE(_231_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[126]_TE  (
    .DIODE(\mprj_logic1[328] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[127]_A  (
    .DIODE(_232_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[127]_TE  (
    .DIODE(\mprj_logic1[329] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[12]_A  (
    .DIODE(_233_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[12]_TE  (
    .DIODE(\mprj_logic1[214] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[13]_A  (
    .DIODE(_234_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[13]_TE  (
    .DIODE(\mprj_logic1[215] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[14]_A  (
    .DIODE(_235_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[14]_TE  (
    .DIODE(\mprj_logic1[216] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[15]_A  (
    .DIODE(_236_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[15]_TE  (
    .DIODE(\mprj_logic1[217] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[16]_A  (
    .DIODE(_237_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[16]_TE  (
    .DIODE(\mprj_logic1[218] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[17]_A  (
    .DIODE(_238_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[17]_TE  (
    .DIODE(\mprj_logic1[219] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[18]_A  (
    .DIODE(_239_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[18]_TE  (
    .DIODE(\mprj_logic1[220] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[19]_A  (
    .DIODE(_240_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[19]_TE  (
    .DIODE(\mprj_logic1[221] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[1]_A  (
    .DIODE(_241_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[1]_TE  (
    .DIODE(\mprj_logic1[203] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[20]_A  (
    .DIODE(_242_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[20]_TE  (
    .DIODE(\mprj_logic1[222] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[21]_A  (
    .DIODE(_243_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[21]_TE  (
    .DIODE(\mprj_logic1[223] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[22]_A  (
    .DIODE(_244_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[22]_TE  (
    .DIODE(\mprj_logic1[224] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[23]_A  (
    .DIODE(_245_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[23]_TE  (
    .DIODE(\mprj_logic1[225] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[24]_A  (
    .DIODE(_246_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[24]_TE  (
    .DIODE(\mprj_logic1[226] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[25]_A  (
    .DIODE(_247_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[25]_TE  (
    .DIODE(\mprj_logic1[227] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[26]_A  (
    .DIODE(_248_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[26]_TE  (
    .DIODE(\mprj_logic1[228] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[27]_A  (
    .DIODE(_249_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[27]_TE  (
    .DIODE(\mprj_logic1[229] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[28]_A  (
    .DIODE(_250_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[28]_TE  (
    .DIODE(\mprj_logic1[230] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[29]_A  (
    .DIODE(_251_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[29]_TE  (
    .DIODE(\mprj_logic1[231] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[2]_A  (
    .DIODE(_252_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[2]_TE  (
    .DIODE(\mprj_logic1[204] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[30]_A  (
    .DIODE(_253_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[30]_TE  (
    .DIODE(\mprj_logic1[232] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[31]_A  (
    .DIODE(_254_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[31]_TE  (
    .DIODE(\mprj_logic1[233] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[32]_A  (
    .DIODE(_255_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[32]_TE  (
    .DIODE(\mprj_logic1[234] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[33]_A  (
    .DIODE(_256_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[33]_TE  (
    .DIODE(\mprj_logic1[235] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[34]_A  (
    .DIODE(_257_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[34]_TE  (
    .DIODE(\mprj_logic1[236] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[35]_A  (
    .DIODE(_258_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[35]_TE  (
    .DIODE(\mprj_logic1[237] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[36]_A  (
    .DIODE(_259_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[36]_TE  (
    .DIODE(\mprj_logic1[238] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[37]_A  (
    .DIODE(_260_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[37]_TE  (
    .DIODE(\mprj_logic1[239] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[38]_A  (
    .DIODE(_261_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[38]_TE  (
    .DIODE(\mprj_logic1[240] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[39]_A  (
    .DIODE(_262_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[39]_TE  (
    .DIODE(\mprj_logic1[241] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[3]_A  (
    .DIODE(_263_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[3]_TE  (
    .DIODE(\mprj_logic1[205] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[40]_A  (
    .DIODE(_264_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[40]_TE  (
    .DIODE(\mprj_logic1[242] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[41]_A  (
    .DIODE(_265_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[41]_TE  (
    .DIODE(\mprj_logic1[243] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[42]_A  (
    .DIODE(_266_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[42]_TE  (
    .DIODE(\mprj_logic1[244] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[43]_A  (
    .DIODE(_267_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[43]_TE  (
    .DIODE(\mprj_logic1[245] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[44]_A  (
    .DIODE(_268_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[44]_TE  (
    .DIODE(\mprj_logic1[246] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[45]_A  (
    .DIODE(_269_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[45]_TE  (
    .DIODE(\mprj_logic1[247] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[46]_A  (
    .DIODE(_270_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[46]_TE  (
    .DIODE(\mprj_logic1[248] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[47]_A  (
    .DIODE(_271_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[47]_TE  (
    .DIODE(\mprj_logic1[249] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[48]_A  (
    .DIODE(_272_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[48]_TE  (
    .DIODE(\mprj_logic1[250] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[49]_A  (
    .DIODE(_273_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[49]_TE  (
    .DIODE(\mprj_logic1[251] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[4]_A  (
    .DIODE(_274_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[4]_TE  (
    .DIODE(\mprj_logic1[206] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[50]_A  (
    .DIODE(_275_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[50]_TE  (
    .DIODE(\mprj_logic1[252] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[51]_A  (
    .DIODE(_276_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[51]_TE  (
    .DIODE(\mprj_logic1[253] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[52]_A  (
    .DIODE(_277_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[52]_TE  (
    .DIODE(\mprj_logic1[254] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[53]_A  (
    .DIODE(_278_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[53]_TE  (
    .DIODE(\mprj_logic1[255] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[54]_A  (
    .DIODE(_279_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[54]_TE  (
    .DIODE(\mprj_logic1[256] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[55]_A  (
    .DIODE(_280_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[55]_TE  (
    .DIODE(\mprj_logic1[257] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[56]_A  (
    .DIODE(_281_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[56]_TE  (
    .DIODE(\mprj_logic1[258] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[57]_A  (
    .DIODE(_282_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[57]_TE  (
    .DIODE(\mprj_logic1[259] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[58]_A  (
    .DIODE(_283_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[58]_TE  (
    .DIODE(\mprj_logic1[260] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[59]_A  (
    .DIODE(_284_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[59]_TE  (
    .DIODE(\mprj_logic1[261] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[5]_A  (
    .DIODE(_285_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[5]_TE  (
    .DIODE(\mprj_logic1[207] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[60]_A  (
    .DIODE(_286_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[60]_TE  (
    .DIODE(\mprj_logic1[262] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[61]_A  (
    .DIODE(_287_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[61]_TE  (
    .DIODE(\mprj_logic1[263] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[62]_A  (
    .DIODE(_288_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[62]_TE  (
    .DIODE(\mprj_logic1[264] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[63]_A  (
    .DIODE(_289_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[63]_TE  (
    .DIODE(\mprj_logic1[265] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[64]_A  (
    .DIODE(_290_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[64]_TE  (
    .DIODE(\mprj_logic1[266] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[65]_A  (
    .DIODE(_291_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[65]_TE  (
    .DIODE(\mprj_logic1[267] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[66]_A  (
    .DIODE(_292_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[66]_TE  (
    .DIODE(\mprj_logic1[268] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[67]_A  (
    .DIODE(_293_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[67]_TE  (
    .DIODE(\mprj_logic1[269] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[68]_A  (
    .DIODE(_294_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[68]_TE  (
    .DIODE(\mprj_logic1[270] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[69]_A  (
    .DIODE(_295_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[69]_TE  (
    .DIODE(\mprj_logic1[271] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[6]_A  (
    .DIODE(_296_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[6]_TE  (
    .DIODE(\mprj_logic1[208] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[70]_A  (
    .DIODE(_297_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[70]_TE  (
    .DIODE(\mprj_logic1[272] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[71]_A  (
    .DIODE(_298_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[71]_TE  (
    .DIODE(\mprj_logic1[273] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[72]_A  (
    .DIODE(_299_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[72]_TE  (
    .DIODE(\mprj_logic1[274] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[73]_A  (
    .DIODE(_300_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[73]_TE  (
    .DIODE(\mprj_logic1[275] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[74]_A  (
    .DIODE(_301_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[74]_TE  (
    .DIODE(\mprj_logic1[276] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[75]_A  (
    .DIODE(_302_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[75]_TE  (
    .DIODE(\mprj_logic1[277] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[76]_A  (
    .DIODE(_303_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[76]_TE  (
    .DIODE(\mprj_logic1[278] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[77]_A  (
    .DIODE(_304_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[77]_TE  (
    .DIODE(\mprj_logic1[279] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[78]_A  (
    .DIODE(_305_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[78]_TE  (
    .DIODE(\mprj_logic1[280] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[79]_A  (
    .DIODE(_306_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[79]_TE  (
    .DIODE(\mprj_logic1[281] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[7]_A  (
    .DIODE(_307_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[7]_TE  (
    .DIODE(\mprj_logic1[209] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[80]_A  (
    .DIODE(_308_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[80]_TE  (
    .DIODE(\mprj_logic1[282] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[81]_A  (
    .DIODE(_309_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[81]_TE  (
    .DIODE(\mprj_logic1[283] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[82]_A  (
    .DIODE(_310_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[82]_TE  (
    .DIODE(\mprj_logic1[284] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[83]_A  (
    .DIODE(_311_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[83]_TE  (
    .DIODE(\mprj_logic1[285] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[84]_A  (
    .DIODE(_312_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[84]_TE  (
    .DIODE(\mprj_logic1[286] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[85]_A  (
    .DIODE(_313_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[85]_TE  (
    .DIODE(\mprj_logic1[287] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[86]_A  (
    .DIODE(_314_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[86]_TE  (
    .DIODE(\mprj_logic1[288] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[87]_A  (
    .DIODE(_315_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[87]_TE  (
    .DIODE(\mprj_logic1[289] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[88]_A  (
    .DIODE(_316_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[88]_TE  (
    .DIODE(\mprj_logic1[290] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[89]_A  (
    .DIODE(_317_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[89]_TE  (
    .DIODE(\mprj_logic1[291] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[8]_A  (
    .DIODE(_318_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[8]_TE  (
    .DIODE(\mprj_logic1[210] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[90]_A  (
    .DIODE(_319_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[90]_TE  (
    .DIODE(\mprj_logic1[292] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[91]_A  (
    .DIODE(_320_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[91]_TE  (
    .DIODE(\mprj_logic1[293] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[92]_A  (
    .DIODE(_321_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[92]_TE  (
    .DIODE(\mprj_logic1[294] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[93]_A  (
    .DIODE(_322_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[93]_TE  (
    .DIODE(\mprj_logic1[295] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[94]_A  (
    .DIODE(_323_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[94]_TE  (
    .DIODE(\mprj_logic1[296] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[95]_A  (
    .DIODE(_324_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[95]_TE  (
    .DIODE(\mprj_logic1[297] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[96]_A  (
    .DIODE(_325_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[96]_TE  (
    .DIODE(\mprj_logic1[298] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[97]_A  (
    .DIODE(_326_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[97]_TE  (
    .DIODE(\mprj_logic1[299] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[98]_A  (
    .DIODE(_327_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[98]_TE  (
    .DIODE(\mprj_logic1[300] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[99]_A  (
    .DIODE(_328_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[99]_TE  (
    .DIODE(\mprj_logic1[301] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[9]_A  (
    .DIODE(_329_),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_oen_buffers[9]_TE  (
    .DIODE(\mprj_logic1[211] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1007 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1019 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1050 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1081 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1093 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1124 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1143 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1155 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1162 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1174 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1193 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1205 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1248 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_125 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1255 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1286 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1298 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1310 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1317 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_1326 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_1346 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1348 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_137 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_149 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_156 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_168 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1780 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_1792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1797 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1809 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1821 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1828 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1840 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1852 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1859 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_187 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1871 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1883 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1890 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1902 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1914 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1933 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1945 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_195 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1952 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1964 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_1976 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1983 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_1995 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2007 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_201 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2045 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_205 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2057 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2076 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2088 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_2119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_2131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_2138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_218 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_232 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_261 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_54 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_58 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_63 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_630 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_659 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_666 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_678 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_690 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_728 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_740 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_75 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_752 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_759 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_771 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_783 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_790 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_802 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_814 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_821 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_83 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_833 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_845 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_852 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_864 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_87 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_876 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_883 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_895 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_907 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_914 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_926 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_938 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_94 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_945 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_957 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_969 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_976 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_988 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_1004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1020 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1051 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1063 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_1088 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1124 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1149 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_1161 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1167 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1170 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1174 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1188 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1238 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1252 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1264 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1295 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1307 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1311 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_1325 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1333 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1341 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1374 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1382 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_150 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_174 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1771 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1775 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1779 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1783 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1791 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_1815 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1870 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1882 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1894 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1919 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_1935 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1941 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_1977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_1992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2002 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_2038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_2068 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_2074 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_2077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_2082 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2086 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_2098 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_2105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_2133 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_2145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_251 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_312 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_317 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_321 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_325 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_329 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_333 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_337 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_341 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_345 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_351 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_354 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_361 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_371 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_383 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_395 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_417 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_430 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_434 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_455 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_463 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_467 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_475 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_481 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_485 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_497 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_505 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_509 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_513 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_532 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_536 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_539 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_55 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_551 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_555 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_570 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_578 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_625 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_629 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_662 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_673 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_678 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_690 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_71 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_715 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_725 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_748 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_760 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_773 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_785 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_804 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_808 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_820 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_83 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_845 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_857 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_869 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_880 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_928 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_940 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_959 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_96 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_971 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_983 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1007 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1011 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1017 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1021 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1027 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1030 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1035 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1060 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1064 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1091 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1097 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1152 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1158 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1210 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1214 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1221 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1225 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1240 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1252 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1264 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_127 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1274 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1278 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1287 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1301 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1338 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1351 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_139 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1394 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1402 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1404 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1429 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1433 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1437 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1441 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1449 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1453 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1462 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1468 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1472 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1476 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_151 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1544 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1553 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1557 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1561 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1565 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1572 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1584 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1597 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1601 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1610 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1627 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_163 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1646 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1666 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1674 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1682 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1690 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1706 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1713 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1717 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1725 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1742 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1749 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1753 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1765 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_1770 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1776 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1780 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1784 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_1788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1821 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1847 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1859 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1871 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_188 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_1883 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_1943 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_1953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1957 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1969 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1981 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_1993 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_2005 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_2009 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_2012 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_2022 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_2038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_2050 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_2067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_2093 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_2097 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_2103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_2107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_2111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_2123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_2136 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_232 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_240 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_251 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_278 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_290 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_297 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_311 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_322 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_326 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_332 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_347 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_391 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_397 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_400 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_409 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_413 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_417 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_423 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_426 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_432 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_436 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_439 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_447 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_455 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_480 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_484 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_507 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_511 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_523 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_535 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_554 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_585 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_600 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_629 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_633 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_645 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_657 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_669 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_672 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_680 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_685 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_716 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_720 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_728 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_74 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_748 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_752 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_764 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_772 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_798 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_802 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_810 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_815 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_842 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_846 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_849 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_853 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_86 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_861 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_865 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_897 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_901 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_914 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_920 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_928 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_11_933 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_938 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_950 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_962 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_975 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_98 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_981 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_996 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1017 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1021 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1035 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1039 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1044 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1048 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1060 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1073 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1085 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_1097 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1152 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1164 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1191 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1250 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1252 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1264 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1303 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1311 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1338 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1361 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1374 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1378 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1382 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1394 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1406 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1418 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1433 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1435 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_1440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_1448 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1454 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1458 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1462 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1466 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1478 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1486 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1491 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1499 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1503 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1527 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1535 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1539 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1547 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1552 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1557 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1561 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1588 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1592 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1596 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1600 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1610 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1614 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1627 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1631 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1646 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1656 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1660 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1664 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1669 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1673 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1677 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1679 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1683 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1687 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1693 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1701 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1720 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1732 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1735 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1740 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1756 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1780 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_1791 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1796 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_1855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1862 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1874 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1886 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_1898 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1923 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1927 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1954 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1966 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_1978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_1982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1984 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_1996 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_2008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_2040 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_2045 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_2057 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_2102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_2106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_2118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_2130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_2142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_233 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_253 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_265 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_291 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_325 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_337 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_349 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_361 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_373 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_385 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_422 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_441 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_453 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_457 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_465 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_474 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_486 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_491 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_503 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_515 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_532 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_546 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_558 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_565 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_585 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_597 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_607 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_617 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_628 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_632 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_640 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_664 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_669 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_673 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_685 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_689 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_693 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_701 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_71 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_715 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_723 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_734 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_748 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_752 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_760 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_764 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_772 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_776 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_800 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_815 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_83 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_833 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_849 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_861 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_873 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_886 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_890 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_894 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_919 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_927 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_938 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_959 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_967 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_12_986 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1017 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1021 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1048 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1052 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1084 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1088 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1096 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1143 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1155 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1177 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1199 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1203 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1207 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1211 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1255 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1364 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1368 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1376 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1402 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1404 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1408 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1418 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1424 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1431 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1454 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1458 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1465 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1477 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1481 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1484 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1498 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1502 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1515 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1566 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1570 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1574 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1578 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1591 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_1603 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1627 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1631 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1641 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1645 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1648 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1652 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1656 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1660 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1664 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1672 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1676 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1680 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1704 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1714 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1718 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1730 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1742 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1754 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1766 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1812 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1816 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_182 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_1820 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1829 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1867 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1912 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1935 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_1947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_1977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_1985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_1989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_2003 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_2009 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_2012 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2020 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2042 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_2046 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_2051 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_2073 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_2075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_2087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_2091 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_2136 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_291 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_302 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_309 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_317 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_329 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_339 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_345 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_371 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_383 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_395 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_407 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_413 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_432 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_444 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_448 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_452 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_472 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_476 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_507 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_511 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_523 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_527 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_554 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_566 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_585 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_590 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_594 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_602 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_620 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_624 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_636 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_655 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_659 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_66 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_669 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_69 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_699 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_707 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_719 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_13_727 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_73 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_752 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_756 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_760 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_777 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_781 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_806 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_837 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_850 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_859 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_871 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_883 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_895 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_899 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_911 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_92 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_929 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_941 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_96 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_13_965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_973 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1348 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1356 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1392 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1399 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1447 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1463 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_1475 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1500 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1504 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1510 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1514 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1518 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1521 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1525 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1529 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1533 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1537 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1547 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1559 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1571 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1591 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1608 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1650 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1662 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1673 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1692 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1696 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1716 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1724 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1750 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1762 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1772 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_1784 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_1787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1793 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1796 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1808 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1893 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_1905 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1915 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1927 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_194 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_1963 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_1982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_1986 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_2005 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_2009 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_2043 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_2092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_2096 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_2124 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_2136 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_219 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_247 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_259 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_271 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_310 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_322 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_359 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_363 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_375 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_395 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_432 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_444 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_45 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_452 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_456 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_483 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_491 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_495 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_509 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_514 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_518 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_532 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_551 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_563 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_590 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_602 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_14_610 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_615 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_627 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_76 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_88 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_127 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1344 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1356 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1368 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_1380 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_139 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1437 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1441 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1447 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1463 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1475 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1487 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_151 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1510 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1517 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1523 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1540 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1552 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1560 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1565 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1613 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1625 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_163 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1634 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1644 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1666 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1670 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1682 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1688 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1692 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_1695 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1701 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1730 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1734 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1746 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1754 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1786 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1791 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_1796 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1802 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1805 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_1817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1859 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1863 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1875 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1878 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1890 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1902 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1928 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_1932 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1943 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1956 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_1968 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_1988 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_1992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_1998 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_2000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_2006 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_2018 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_2030 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_2035 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_2039 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_2067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_2107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_2111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_2115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_234 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_281 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_324 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_328 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_332 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_361 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_384 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_408 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_412 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_415 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_419 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_423 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_15_432 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_478 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_498 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_502 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_525 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_529 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_15_543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_554 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_558 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_573 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_589 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_602 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_15_66 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_73 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_77 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_96 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_113 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1347 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1384 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1415 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1419 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1449 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1453 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1465 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1477 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_16_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1490 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_1502 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1525 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1537 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1541 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1555 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1585 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1589 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1601 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1616 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1628 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1640 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1644 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_16_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1663 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1669 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1711 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1714 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_1722 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_174 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_16_1750 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1758 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1770 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1807 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_1843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_1927 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1958 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_1966 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_1982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_2008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_2020 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_2031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_2069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_2073 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_2087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_210 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_233 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_16_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_289 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_293 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_303 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_308 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_320 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_326 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_374 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_394 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_431 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_439 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_444 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_463 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_475 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_487 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_508 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_536 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_558 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_568 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_597 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_16_75 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_88 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_108 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1402 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1405 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1424 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1457 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1461 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1473 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1485 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1497 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1509 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1516 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1541 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1545 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1549 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_156 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1570 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1573 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1580 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1584 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1603 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1607 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1619 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_1626 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1632 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1634 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1640 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1652 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1664 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_1676 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1684 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1713 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1717 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1729 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_1741 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1747 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_1756 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_176 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1761 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_1773 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1812 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1821 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1829 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1833 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1845 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1857 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1869 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_1878 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_188 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1883 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1905 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_1913 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_1929 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1935 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1957 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_1984 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_1996 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_2000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_2008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_2013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_2025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_2033 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_2047 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_2053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_2059 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_2073 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_2085 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_2088 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_2120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_235 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_253 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_302 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_310 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_321 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_346 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_17_35 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_350 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_353 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_391 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_403 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_413 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_462 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_466 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_478 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_484 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_507 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_511 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_523 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_527 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_530 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_547 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_574 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_580 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_583 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_597 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_66 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_96 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1384 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1404 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1408 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1439 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1463 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1467 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1479 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1494 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1510 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_152 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1529 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1533 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1541 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_1551 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_1556 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_158 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_1582 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1616 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_162 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1662 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1677 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_170 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1700 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1704 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1716 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1724 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_1738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1763 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1775 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1805 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1809 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_1872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1880 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1899 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1903 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1907 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_1945 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1964 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1968 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_1982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_1988 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_1994 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_2015 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_2027 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_2049 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_2073 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_2085 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_2126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_2138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_295 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_308 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_329 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_391 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_402 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_429 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_433 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_447 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_455 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_483 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_504 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_508 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_516 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_539 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_551 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_563 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_575 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_579 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_63 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_67 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_75 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_18_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_113 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1352 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1364 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1376 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_1388 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1403 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1417 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1446 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1475 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1479 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1491 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1503 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1536 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_1548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_157 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1573 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_1581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1591 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_1603 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1631 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1634 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1638 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1650 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1658 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1679 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1683 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_169 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1691 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1695 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1707 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_1721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_1725 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1728 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1742 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1746 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_1754 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1756 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1760 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_1772 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1797 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1801 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_181 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_1847 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_1868 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_1872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_1876 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1878 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1890 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1902 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_1930 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_1963 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_1975 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_2000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_2004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_2016 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_2040 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_2048 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_2051 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_2059 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_2077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_2126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_2138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_222 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_238 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_271 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_287 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_299 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_338 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_35 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_362 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_407 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_411 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_424 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_470 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_474 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_486 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_513 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_52 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_525 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_530 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_535 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_568 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_572 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_584 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_596 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_19_604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_19_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_84 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_92 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_95 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1006 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1018 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1043 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1055 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1153 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1165 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1177 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1189 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1201 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1211 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1214 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1238 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1250 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_1262 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1268 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_1271 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1287 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1292 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1296 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1308 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1317 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_1329 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_133 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1336 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1348 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_1384 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_157 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_169 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1780 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1804 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_181 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_1816 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1824 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1851 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1863 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1875 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1912 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1924 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1936 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1973 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_1985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_1989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2022 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2034 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2046 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2058 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_2079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_2128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_2132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_220 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_232 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_281 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_630 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_662 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_677 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_689 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_701 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_713 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_74 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_750 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_762 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_811 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_86 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_929 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_933 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_945 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_957 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_98 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_994 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_133 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_1352 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1384 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1400 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1419 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1494 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1518 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1530 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1551 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1589 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1601 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_1604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1625 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1629 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1641 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_1653 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1663 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1677 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1689 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1701 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1723 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1762 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1781 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1785 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_1811 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1852 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1864 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1876 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_1888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_1893 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1903 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1907 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1913 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1932 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1944 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_1956 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_1968 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_1978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_1983 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_2004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_2016 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_2031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_2043 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_2067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_2079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_2087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_2126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_2138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_300 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_312 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_324 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_337 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_354 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_366 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_378 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_20_386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_391 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_418 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_430 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_449 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_453 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_457 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_465 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_469 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_481 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_493 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_496 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_500 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_510 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_514 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_518 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_535 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_547 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_567 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_571 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_579 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_20_621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_75 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_79 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1352 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1364 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_1376 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1380 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1383 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1388 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1402 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1405 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_143 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1436 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1444 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1448 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1455 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1483 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1495 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1503 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1530 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1534 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1546 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1558 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1570 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1573 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1589 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1601 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1613 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1625 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1634 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_1638 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1662 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1666 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1678 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1682 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1695 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1699 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1720 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1741 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1745 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1756 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1764 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1769 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1781 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_179 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1793 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1801 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1804 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1812 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_1817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_182 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1842 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1854 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1864 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1876 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1878 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_1882 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1886 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1889 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1913 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1933 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_1937 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_1963 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_1989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_1993 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_2000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_2012 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_2024 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_2036 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_2044 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_2049 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_2057 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_21_2075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_210 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_2101 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_2105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_2109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_222 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_297 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_301 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_35 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_350 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_353 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_371 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_383 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_406 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_422 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_426 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_434 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_438 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_446 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_467 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_477 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_481 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_485 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_21_489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_493 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_523 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_21_527 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_542 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_546 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_21_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_565 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_58 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_21_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_589 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_598 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_21_623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_66 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_21_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_21_74 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_79 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_113 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_1352 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_1372 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1378 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1388 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1400 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_1404 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1408 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_1411 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1415 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1418 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1444 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1455 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1467 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1479 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_1494 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_150 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1502 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1522 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1526 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_1538 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_1555 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1559 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1578 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1590 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1602 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1616 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_1628 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1634 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1653 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_1657 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1663 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_1669 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_1677 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_1698 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1704 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_1718 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1722 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_1750 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1771 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_1775 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_1783 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1820 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1824 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_1836 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_1844 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_1880 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1886 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_1905 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1913 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1917 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_1929 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_198 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_1982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_2001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_2013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_2025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_2029 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_2031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_2039 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_2044 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_2092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_2096 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_2108 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_2120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_2132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_223 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_234 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_254 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_260 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_298 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_310 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_314 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_322 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_337 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_349 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_369 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_381 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_422 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_434 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_446 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_457 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_477 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_485 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_515 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_532 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_537 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_549 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_557 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_560 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_572 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_598 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_607 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_619 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_624 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_628 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_22_81 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_22_89 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1359 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1362 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1376 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_23_1382 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1394 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_23_1413 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1429 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1433 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1445 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1449 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1475 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1487 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1499 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1503 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1510 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_1512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1539 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_23_1569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1573 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1585 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1597 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_1621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1629 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_163 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1670 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1674 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1678 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1693 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1695 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1707 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_1719 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1725 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1728 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1742 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1754 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_1806 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1814 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1829 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1841 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1853 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1865 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_1915 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_1919 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_23_192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1937 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1963 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_197 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1975 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_1978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_1992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_1998 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_2000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_2012 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_2077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_2085 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_2106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_211 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_2120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_23_223 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_261 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_285 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_291 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_324 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_328 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_332 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_35 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_353 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_385 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_389 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_401 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_413 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_419 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_422 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_426 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_436 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_448 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_460 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_472 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_484 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_493 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_540 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_574 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_586 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_23_603 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_607 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_23_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_625 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_23_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_74 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_88 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_1387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_1397 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_1401 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1425 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1429 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_143 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1441 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1455 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1467 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1479 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_1486 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1494 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1498 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_151 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1522 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1526 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_1538 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_1543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1553 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1567 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1579 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1591 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1616 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1628 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1648 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1652 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_1656 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_1660 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1683 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1695 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1707 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1719 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1758 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1811 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1880 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_1886 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_1907 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1927 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_194 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1951 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1963 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_1994 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_2006 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_2018 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_2031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_2037 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_2040 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_2060 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_2064 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_2076 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_2090 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_2110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_2122 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_213 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_2134 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_219 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_225 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_250 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_262 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_274 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_307 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_311 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_337 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_349 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_361 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_369 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_381 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_393 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_418 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_438 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_450 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_483 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_24_491 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_24_516 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_531 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_543 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_555 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_567 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_579 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_24_589 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_24_594 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_602 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_612 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_616 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_90 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1019 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1023 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1035 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1047 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1051 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_1075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1096 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_1111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_1154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1158 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_1160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1164 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1176 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_1208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_1213 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1219 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1221 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_1229 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1241 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1261 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1265 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1291 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1295 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1307 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1315 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1337 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1341 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1347 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1359 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1371 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1383 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1395 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1422 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1426 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1438 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1450 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1462 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_1465 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1473 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1481 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1502 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_1506 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1526 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_1538 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1544 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1563 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1567 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_157 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_1579 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1585 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_1644 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1648 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1652 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1664 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_169 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1690 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1694 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1706 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_1745 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1749 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1770 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1786 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1798 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_1810 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1816 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_1819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1849 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1853 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1865 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1877 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_189 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_1892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_1899 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_1903 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1922 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1926 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1938 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_1950 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_1989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_201 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_2038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2044 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2056 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_2068 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_2123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_2136 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_222 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_232 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_281 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_289 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_303 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_324 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_328 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_336 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_339 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_353 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_373 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_405 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_409 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_421 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_446 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_450 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_469 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_473 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_485 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_524 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_544 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_548 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_554 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_558 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_563 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_575 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_607 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_619 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_638 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_66 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_25_666 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_670 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_693 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_730 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_746 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_750 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_762 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_25_794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_815 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_849 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_853 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_891 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_895 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_899 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_903 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_934 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_945 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_95 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_25_957 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_25_974 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1042 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_1054 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_1057 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1066 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_1077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_1082 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_1087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_1162 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1176 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1186 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1191 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1195 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_1233 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_1236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1241 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1247 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_125 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1270 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1286 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1298 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1310 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1313 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1321 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1345 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1369 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_137 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1374 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1406 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1418 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1430 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1435 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1447 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_149 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1514 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1526 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1538 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_1544 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1547 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_1555 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1557 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1569 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1605 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1646 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1650 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1662 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1670 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1674 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1679 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1691 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1715 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_172 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1727 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1740 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1748 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1752 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1764 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1776 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1801 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_1851 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_1859 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1862 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1874 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1886 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_1898 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_191 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_1918 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1923 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1935 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1959 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1971 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1984 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_1996 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2020 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_203 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2032 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2045 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2057 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2081 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2093 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_2130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_2142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_234 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_246 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_258 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_270 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_274 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_305 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_309 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_321 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_333 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_389 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_393 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_398 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_410 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_422 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_43 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_430 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_442 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_450 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_453 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_457 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_47 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_471 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_483 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_495 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_504 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_516 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_565 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_577 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_581 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_593 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_605 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_617 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_622 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_634 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_640 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_666 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_676 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_685 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_688 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_700 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_711 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_716 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_725 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_737 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_741 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_753 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_761 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_764 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_776 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_784 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_797 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_837 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_841 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_844 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_856 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_859 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_864 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_876 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_882 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_895 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_899 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_911 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_917 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_920 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_939 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_943 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_959 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_969 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_97 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_974 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_981 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_986 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_26_990 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_995 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_26_999 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1050 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1074 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1086 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1172 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_27_121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1221 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1233 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_1245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_27_1253 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1256 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1268 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_27_1280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1391 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1404 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1452 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1465 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1477 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1513 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1526 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1538 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1574 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1587 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1599 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1648 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1660 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1672 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1684 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1696 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_27_1721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_1745 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1749 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_1761 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1770 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1806 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1867 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1879 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1928 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1940 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_1989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2050 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_2123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_2136 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_218 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_281 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_293 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_354 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_391 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_403 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_415 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_452 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_464 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_476 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_513 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_525 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_537 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_562 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_574 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_586 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_598 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_27_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_623 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_659 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_672 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_684 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_696 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_708 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_720 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_745 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_757 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_769 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_781 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_798 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_802 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_806 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_81 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_810 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_822 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_834 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_846 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_85 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_27_855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_27_861 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_864 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_27_868 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_873 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_877 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_881 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_893 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_905 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_27_913 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_27_924 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_929 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_941 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_953 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_27_965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_97 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_27_973 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1005 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1017 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1024 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1036 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1048 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1055 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1086 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1098 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1148 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1172 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1179 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1191 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1203 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1210 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1222 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1234 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1241 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_125 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1253 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1265 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1272 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1296 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1303 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1315 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1327 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1346 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_137 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1377 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1389 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1396 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1408 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1420 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1427 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1439 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1451 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1458 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1470 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1482 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1489 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_149 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1513 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1532 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1544 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1551 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_156 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1563 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1575 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1582 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1594 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1613 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1625 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1637 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1644 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1656 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1668 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1675 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_168 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1687 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1699 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1706 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_28_1718 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_28_1726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1729 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_28_1735 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1737 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1749 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1761 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1780 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_28_180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1811 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1830 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1842 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1854 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1861 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_187 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1873 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1885 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1923 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1935 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1954 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1966 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_1978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_199 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_1997 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_2009 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2016 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_2040 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2047 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2059 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2078 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2090 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_2102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_211 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_2121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_2133 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_2140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_218 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_249 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_261 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_28_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_292 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_304 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_311 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_28_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_323 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_335 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_354 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_366 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_373 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_385 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_397 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_28_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_404 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_428 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_28_43 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_435 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_447 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_459 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_466 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_478 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_490 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_497 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_509 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_28_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_521 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_528 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_540 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_28_55 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_552 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_559 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_571 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_583 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_28_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_590 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_602 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_614 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_28_63 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_633 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_645 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_652 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_664 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_67 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_676 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_683 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_695 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_707 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_714 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_745 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_757 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_769 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_776 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_79 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_800 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_807 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_850 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_862 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_869 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_881 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_893 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_28_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_912 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_924 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_94 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_943 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_955 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_962 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_974 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_986 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_993 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1037 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1049 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1074 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1086 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1098 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_1208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_125 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1272 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_1295 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_1303 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_133 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1336 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1348 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1360 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1780 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_1792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1797 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1809 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1821 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1833 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1845 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1870 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1882 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1894 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1919 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1943 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1955 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1967 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_1998 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2022 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_2034 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_2077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2083 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_2095 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_2126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_2138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_251 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_286 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_610 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_622 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_659 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_671 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_68 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_683 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_696 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_708 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_720 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_732 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_757 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_769 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_781 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_793 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_805 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_830 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_842 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_854 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_866 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_879 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_887 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_899 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_911 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_923 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_936 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_940 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_952 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_964 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_976 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_988 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1009 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1029 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1043 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1055 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1140 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1153 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1183 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1197 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1203 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1207 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1214 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1219 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1225 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1254 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1266 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1283 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1295 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1307 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1315 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1320 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1324 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1328 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1332 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1336 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1347 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1351 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1355 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1359 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1371 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1383 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1768 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1772 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1776 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1788 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1805 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1834 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1846 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1870 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_188 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1880 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_1884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1910 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1922 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1930 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_1942 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_1973 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_1981 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_1997 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_2022 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2027 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2039 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_2051 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_2058 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_2062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_2079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2083 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2095 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_2132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_229 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_241 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_253 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_256 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_268 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_272 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_294 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_613 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_617 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_629 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_641 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_653 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_661 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_67 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_673 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_678 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_690 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_702 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_71 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_714 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_722 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_759 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_76 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_763 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_767 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_779 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_785 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_811 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_823 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_889 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_893 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_906 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_92 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_933 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_941 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_946 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_958 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_966 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_995 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_999 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1037 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1049 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1074 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1086 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1098 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1155 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1172 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1198 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1210 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1222 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1284 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1296 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1304 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1314 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1319 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1331 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1339 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1351 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1363 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_1379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_178 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_1786 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1795 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1800 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1806 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1830 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1835 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1847 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1870 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_1911 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1917 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_1919 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_1927 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1943 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1955 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1967 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1986 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_1998 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_2077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2084 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_2096 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_2100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_2126 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_2138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_218 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_242 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_612 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_624 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_632 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_659 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_671 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_68 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_693 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_696 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_708 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_720 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_732 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_744 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_766 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_790 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_802 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_814 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_830 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_836 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_846 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_4_870 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_879 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_891 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_895 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_905 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_933 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_973 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_997 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1006 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1018 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1035 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1047 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1055 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1067 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1127 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1143 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1151 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1153 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1165 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1173 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1176 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1180 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1199 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1205 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1209 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1221 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1255 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1267 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1287 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1291 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1298 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1302 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1336 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1340 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1349 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1353 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1362 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1374 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1377 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1389 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_165 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1771 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1775 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1779 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1791 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1797 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1800 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1812 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1844 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_1884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_1888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1908 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1920 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1934 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1946 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_1957 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_1977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1985 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_1989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_1993 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_200 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_2001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_2015 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_2027 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2036 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2040 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2045 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_2049 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_2069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2084 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_2088 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_2094 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_2097 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_2101 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_2104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_2116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_2128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_2132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_220 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_225 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_235 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_248 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_252 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_256 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_259 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_271 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_278 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_288 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_52 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_609 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_613 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_617 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_621 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_633 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_645 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_65 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_657 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_663 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_665 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_677 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_689 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_69 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_702 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_714 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_718 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_724 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_743 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_747 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_751 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_763 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_767 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_771 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_783 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_81 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_812 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_816 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_826 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_857 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_861 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_865 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_876 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_880 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_913 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_5_937 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_950 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_954 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_958 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_964 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_967 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_99 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_994 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_1013 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1017 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1037 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1058 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1062 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1074 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1082 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1094 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_1118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_1166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_1179 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_121 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1224 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1236 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1281 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1293 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_133 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1342 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1354 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1378 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_160 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_164 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_168 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_172 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_1790 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1797 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1801 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1821 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1856 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1870 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1882 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_1890 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1895 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1903 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1907 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_1915 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1919 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1935 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1947 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_1959 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_1971 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_1986 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_1993 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_2002 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2016 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_2072 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_2076 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2080 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_2092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_2098 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_2129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_2141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_2145 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_226 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_241 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_253 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_260 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_272 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_291 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_624 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_632 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_659 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_671 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_683 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_705 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_711 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_72 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_721 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_739 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_749 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_755 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_766 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_790 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_802 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_807 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_815 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_829 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_84 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_846 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_6_867 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_875 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_879 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_891 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_912 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_924 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_6_936 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_940 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_982 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_994 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1000 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1029 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1031 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1035 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1039 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1051 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1063 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1068 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1080 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1083 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1092 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_1131 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1148 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1153 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1158 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1170 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1182 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1194 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_1206 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1214 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1218 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1240 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1252 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1264 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1272 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1287 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1299 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1311 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1319 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1325 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_1329 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1336 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1347 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1351 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1363 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1375 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_155 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_161 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_165 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1794 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1804 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1808 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_181 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1834 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1850 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1854 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1862 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1866 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_1878 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_188 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1883 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_1888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1914 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1918 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1937 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1942 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1946 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1965 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_1969 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_1976 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_1992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_2004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_2008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_2022 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2033 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_204 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2045 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_2049 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_2061 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_2069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_2075 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2079 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2083 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_2087 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_2093 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_2097 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_212 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_2120 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_2128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_2132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_218 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_222 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_228 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_235 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_281 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_285 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_289 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_52 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_630 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_642 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_654 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_674 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_678 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_690 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_698 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_703 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_715 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_723 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_726 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_738 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_750 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_762 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_77 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_791 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_81 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_810 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_814 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_826 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_846 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_848 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_852 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_864 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_872 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_921 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_925 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_931 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_934 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_942 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_946 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_7_958 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_963 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_7_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_974 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_984 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_988 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_1001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1005 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_1008 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1020 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1024 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_1071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1086 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1098 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1161 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1173 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1181 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_1217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1221 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1265 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1268 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1280 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_129 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1292 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1304 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1318 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1330 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1345 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1357 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1387 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_141 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_154 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_166 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1771 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1775 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1787 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1795 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1800 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_1812 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1819 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1831 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1838 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1850 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_1858 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1867 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1879 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_1896 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_190 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1901 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_1909 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1922 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1934 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1946 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1958 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_1970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_1978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_1992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2004 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2016 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_202 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_2028 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_2032 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2041 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2053 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2065 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_2077 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_2090 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_2094 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_2100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_2102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_2130 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_2142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_215 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_227 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_251 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_263 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_276 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_289 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_49 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_53 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_606 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_618 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_630 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_635 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_65 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_655 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_667 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_679 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_691 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_696 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_706 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_718 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_730 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_742 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_754 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_757 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_769 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_77 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_781 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_793 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_830 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_851 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_863 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_875 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_879 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_8_89 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_891 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_903 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_915 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_937 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_966 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_978 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_981 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_8_991 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_999 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1001 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1005 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1017 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1025 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1030 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1036 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1042 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1048 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1060 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1072 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1076 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1082 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1085 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1097 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1099 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1127 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1138 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1142 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1146 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1158 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1169 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1173 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1179 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1192 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1197 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1209 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1217 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_123 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1230 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1234 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1238 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1246 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1258 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1262 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1273 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1277 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1282 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1286 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1292 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1304 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1316 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1328 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1338 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1343 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1347 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_135 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1352 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1362 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1366 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1374 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1378 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1382 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_147 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_159 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_167 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_171 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_175 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1774 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1778 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1786 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_179 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1795 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1799 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1805 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1809 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_1813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1818 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1822 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1827 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1839 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_184 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1851 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1856 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_1860 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1869 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1873 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1885 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1900 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1904 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1908 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1912 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_1920 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1924 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1928 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_1940 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1949 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_196 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1961 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1973 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_1980 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_1984 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_1996 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_2006 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_2010 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2014 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2026 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2038 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_2050 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_2059 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_2063 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_2069 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2071 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_208 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2083 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_2095 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_2108 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_2112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_2128 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_2132 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_2144 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_216 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_221 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_225 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_231 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_235 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_239 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_243 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_245 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_257 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_269 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_275 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_279 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_283 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_295 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_303 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_306 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_314 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_324 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_334 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_338 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_348 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_358 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_365 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_367 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_375 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_379 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_386 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_390 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_394 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_407 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_41 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_411 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_416 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_420 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_434 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_440 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_456 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_485 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_501 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_512 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_516 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_520 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_526 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_530 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_534 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_54 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_546 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_550 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_555 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_559 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_563 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_567 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_575 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_58 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_582 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_586 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_596 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_600 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_604 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_611 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_615 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_627 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_631 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_637 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_647 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_651 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_663 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_667 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_670 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_681 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_693 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_697 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_709 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_713 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_719 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_722 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_730 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_733 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_74 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_741 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_753 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_765 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_770 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_782 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_792 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_803 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_813 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_817 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_825 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_829 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_84 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_843 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_851 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_855 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_867 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_4 FILLER_9_88 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_884 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_888 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_8 FILLER_9_892 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_902 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_914 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_916 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_92 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_928 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_932 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_944 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_95 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_956 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_966 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_970 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_974 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_977 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_989 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_99 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__fill_2 FILLER_9_992 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_996 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_100 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_101 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_102 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_103 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_104 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_105 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_106 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_107 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_108 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_109 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_110 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_111 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_112 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_113 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_114 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_115 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_116 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_117 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_118 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_119 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_32 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_33 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_34 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_35 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_36 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_37 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_38 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_39 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_40 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_41 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_42 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_43 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_44 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_45 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_46 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_47 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_48 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_49 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_50 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_51 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_52 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_53 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_54 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_55 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_56 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_57 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_58 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_59 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_60 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_61 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_62 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_63 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_64 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_65 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_66 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_67 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_68 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_69 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_70 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_71 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_72 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_73 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_74 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_75 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_76 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_77 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_78 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_79 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_80 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_81 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_82 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_83 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_84 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_85 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_86 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_87 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_88 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_89 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_90 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_91 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_92 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_93 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 (
    .VGND(vssd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_94 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_95 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_96 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_97 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_98 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__decap_3 PHY_99 (
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd)
  );
  sky130_fd_sc_hd__inv_2 _330_ (
    .A(la_oen_mprj[62]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_288_)
  );
  sky130_fd_sc_hd__inv_2 _331_ (
    .A(la_oen_mprj[63]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_289_)
  );
  sky130_fd_sc_hd__inv_2 _332_ (
    .A(la_oen_mprj[64]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_290_)
  );
  sky130_fd_sc_hd__inv_2 _333_ (
    .A(la_oen_mprj[65]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_291_)
  );
  sky130_fd_sc_hd__inv_2 _334_ (
    .A(la_oen_mprj[66]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_292_)
  );
  sky130_fd_sc_hd__inv_2 _335_ (
    .A(la_oen_mprj[67]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_293_)
  );
  sky130_fd_sc_hd__inv_2 _336_ (
    .A(la_oen_mprj[68]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_294_)
  );
  sky130_fd_sc_hd__inv_2 _337_ (
    .A(la_oen_mprj[69]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_295_)
  );
  sky130_fd_sc_hd__inv_2 _338_ (
    .A(la_oen_mprj[70]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_297_)
  );
  sky130_fd_sc_hd__inv_2 _339_ (
    .A(la_oen_mprj[71]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_298_)
  );
  sky130_fd_sc_hd__inv_2 _340_ (
    .A(la_oen_mprj[72]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_299_)
  );
  sky130_fd_sc_hd__inv_2 _341_ (
    .A(la_oen_mprj[73]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_300_)
  );
  sky130_fd_sc_hd__inv_2 _342_ (
    .A(la_oen_mprj[74]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_301_)
  );
  sky130_fd_sc_hd__inv_2 _343_ (
    .A(la_oen_mprj[75]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_302_)
  );
  sky130_fd_sc_hd__inv_2 _344_ (
    .A(la_oen_mprj[76]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_303_)
  );
  sky130_fd_sc_hd__inv_2 _345_ (
    .A(la_oen_mprj[77]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_304_)
  );
  sky130_fd_sc_hd__inv_2 _346_ (
    .A(la_oen_mprj[78]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_305_)
  );
  sky130_fd_sc_hd__inv_2 _347_ (
    .A(la_oen_mprj[79]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_306_)
  );
  sky130_fd_sc_hd__inv_2 _348_ (
    .A(la_oen_mprj[80]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_308_)
  );
  sky130_fd_sc_hd__inv_2 _349_ (
    .A(la_oen_mprj[81]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_309_)
  );
  sky130_fd_sc_hd__inv_2 _350_ (
    .A(la_oen_mprj[82]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_310_)
  );
  sky130_fd_sc_hd__inv_2 _351_ (
    .A(la_oen_mprj[83]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_311_)
  );
  sky130_fd_sc_hd__inv_2 _352_ (
    .A(la_oen_mprj[84]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_312_)
  );
  sky130_fd_sc_hd__inv_2 _353_ (
    .A(la_oen_mprj[85]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_313_)
  );
  sky130_fd_sc_hd__inv_2 _354_ (
    .A(la_oen_mprj[86]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_314_)
  );
  sky130_fd_sc_hd__inv_2 _355_ (
    .A(la_oen_mprj[87]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_315_)
  );
  sky130_fd_sc_hd__inv_2 _356_ (
    .A(la_oen_mprj[88]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_316_)
  );
  sky130_fd_sc_hd__inv_2 _357_ (
    .A(la_oen_mprj[89]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_317_)
  );
  sky130_fd_sc_hd__inv_2 _358_ (
    .A(la_oen_mprj[90]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_319_)
  );
  sky130_fd_sc_hd__inv_2 _359_ (
    .A(la_oen_mprj[91]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_320_)
  );
  sky130_fd_sc_hd__inv_2 _360_ (
    .A(la_oen_mprj[92]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_321_)
  );
  sky130_fd_sc_hd__inv_2 _361_ (
    .A(la_oen_mprj[93]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_322_)
  );
  sky130_fd_sc_hd__inv_2 _362_ (
    .A(la_oen_mprj[94]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_323_)
  );
  sky130_fd_sc_hd__inv_2 _363_ (
    .A(la_oen_mprj[95]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_324_)
  );
  sky130_fd_sc_hd__inv_2 _364_ (
    .A(la_oen_mprj[96]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_325_)
  );
  sky130_fd_sc_hd__inv_2 _365_ (
    .A(la_oen_mprj[97]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_326_)
  );
  sky130_fd_sc_hd__inv_2 _366_ (
    .A(la_oen_mprj[98]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_327_)
  );
  sky130_fd_sc_hd__inv_2 _367_ (
    .A(la_oen_mprj[99]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_328_)
  );
  sky130_fd_sc_hd__inv_2 _368_ (
    .A(la_oen_mprj[100]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_203_)
  );
  sky130_fd_sc_hd__inv_2 _369_ (
    .A(la_oen_mprj[101]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_204_)
  );
  sky130_fd_sc_hd__inv_2 _370_ (
    .A(la_oen_mprj[102]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_205_)
  );
  sky130_fd_sc_hd__inv_2 _371_ (
    .A(la_oen_mprj[103]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_206_)
  );
  sky130_fd_sc_hd__inv_2 _372_ (
    .A(la_oen_mprj[104]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_207_)
  );
  sky130_fd_sc_hd__inv_2 _373_ (
    .A(la_oen_mprj[105]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_208_)
  );
  sky130_fd_sc_hd__inv_2 _374_ (
    .A(la_oen_mprj[106]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_209_)
  );
  sky130_fd_sc_hd__inv_2 _375_ (
    .A(la_oen_mprj[107]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_210_)
  );
  sky130_fd_sc_hd__inv_2 _376_ (
    .A(la_oen_mprj[108]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_211_)
  );
  sky130_fd_sc_hd__inv_2 _377_ (
    .A(la_oen_mprj[109]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_212_)
  );
  sky130_fd_sc_hd__inv_2 _378_ (
    .A(la_oen_mprj[110]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_214_)
  );
  sky130_fd_sc_hd__inv_2 _379_ (
    .A(la_oen_mprj[111]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_215_)
  );
  sky130_fd_sc_hd__inv_2 _380_ (
    .A(la_oen_mprj[112]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_216_)
  );
  sky130_fd_sc_hd__inv_2 _381_ (
    .A(la_oen_mprj[113]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_217_)
  );
  sky130_fd_sc_hd__inv_2 _382_ (
    .A(la_oen_mprj[114]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_218_)
  );
  sky130_fd_sc_hd__inv_2 _383_ (
    .A(la_oen_mprj[115]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_219_)
  );
  sky130_fd_sc_hd__inv_2 _384_ (
    .A(la_oen_mprj[116]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_220_)
  );
  sky130_fd_sc_hd__inv_2 _385_ (
    .A(la_oen_mprj[117]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_221_)
  );
  sky130_fd_sc_hd__inv_2 _386_ (
    .A(la_oen_mprj[118]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_222_)
  );
  sky130_fd_sc_hd__inv_2 _387_ (
    .A(la_oen_mprj[119]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_223_)
  );
  sky130_fd_sc_hd__inv_2 _388_ (
    .A(la_oen_mprj[120]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_225_)
  );
  sky130_fd_sc_hd__inv_2 _389_ (
    .A(la_oen_mprj[121]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_226_)
  );
  sky130_fd_sc_hd__inv_2 _390_ (
    .A(la_oen_mprj[122]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_227_)
  );
  sky130_fd_sc_hd__inv_2 _391_ (
    .A(la_oen_mprj[123]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_228_)
  );
  sky130_fd_sc_hd__inv_2 _392_ (
    .A(la_oen_mprj[124]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_229_)
  );
  sky130_fd_sc_hd__inv_2 _393_ (
    .A(la_oen_mprj[125]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_230_)
  );
  sky130_fd_sc_hd__inv_2 _394_ (
    .A(la_oen_mprj[126]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_231_)
  );
  sky130_fd_sc_hd__inv_2 _395_ (
    .A(la_oen_mprj[127]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_232_)
  );
  sky130_fd_sc_hd__inv_2 _396_ (
    .A(caravel_rstn),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_000_)
  );
  sky130_fd_sc_hd__inv_2 _397_ (
    .A(user_resetn),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(user_reset)
  );
  sky130_fd_sc_hd__inv_2 _398_ (
    .A(caravel_clk),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_001_)
  );
  sky130_fd_sc_hd__inv_2 _399_ (
    .A(caravel_clk2),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_002_)
  );
  sky130_fd_sc_hd__inv_2 _400_ (
    .A(mprj_cyc_o_core),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_003_)
  );
  sky130_fd_sc_hd__inv_2 _401_ (
    .A(mprj_stb_o_core),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_004_)
  );
  sky130_fd_sc_hd__inv_2 _402_ (
    .A(mprj_we_o_core),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_005_)
  );
  sky130_fd_sc_hd__inv_2 _403_ (
    .A(mprj_sel_o_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_006_)
  );
  sky130_fd_sc_hd__inv_2 _404_ (
    .A(mprj_sel_o_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_007_)
  );
  sky130_fd_sc_hd__inv_2 _405_ (
    .A(mprj_sel_o_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_008_)
  );
  sky130_fd_sc_hd__inv_2 _406_ (
    .A(mprj_sel_o_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_009_)
  );
  sky130_fd_sc_hd__inv_2 _407_ (
    .A(mprj_adr_o_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_010_)
  );
  sky130_fd_sc_hd__inv_2 _408_ (
    .A(mprj_adr_o_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_021_)
  );
  sky130_fd_sc_hd__inv_2 _409_ (
    .A(mprj_adr_o_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_032_)
  );
  sky130_fd_sc_hd__inv_2 _410_ (
    .A(mprj_adr_o_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_035_)
  );
  sky130_fd_sc_hd__inv_2 _411_ (
    .A(mprj_adr_o_core[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_036_)
  );
  sky130_fd_sc_hd__inv_2 _412_ (
    .A(mprj_adr_o_core[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_037_)
  );
  sky130_fd_sc_hd__inv_2 _413_ (
    .A(mprj_adr_o_core[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_038_)
  );
  sky130_fd_sc_hd__inv_2 _414_ (
    .A(mprj_adr_o_core[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_039_)
  );
  sky130_fd_sc_hd__inv_2 _415_ (
    .A(mprj_adr_o_core[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_040_)
  );
  sky130_fd_sc_hd__inv_2 _416_ (
    .A(mprj_adr_o_core[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_041_)
  );
  sky130_fd_sc_hd__inv_2 _417_ (
    .A(mprj_adr_o_core[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_011_)
  );
  sky130_fd_sc_hd__inv_2 _418_ (
    .A(mprj_adr_o_core[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_012_)
  );
  sky130_fd_sc_hd__inv_2 _419_ (
    .A(mprj_adr_o_core[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_013_)
  );
  sky130_fd_sc_hd__inv_2 _420_ (
    .A(mprj_adr_o_core[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_014_)
  );
  sky130_fd_sc_hd__inv_2 _421_ (
    .A(mprj_adr_o_core[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_015_)
  );
  sky130_fd_sc_hd__inv_2 _422_ (
    .A(mprj_adr_o_core[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_016_)
  );
  sky130_fd_sc_hd__inv_2 _423_ (
    .A(mprj_adr_o_core[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_017_)
  );
  sky130_fd_sc_hd__inv_2 _424_ (
    .A(mprj_adr_o_core[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_018_)
  );
  sky130_fd_sc_hd__inv_2 _425_ (
    .A(mprj_adr_o_core[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_019_)
  );
  sky130_fd_sc_hd__inv_2 _426_ (
    .A(mprj_adr_o_core[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_020_)
  );
  sky130_fd_sc_hd__inv_2 _427_ (
    .A(mprj_adr_o_core[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_022_)
  );
  sky130_fd_sc_hd__inv_2 _428_ (
    .A(mprj_adr_o_core[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_023_)
  );
  sky130_fd_sc_hd__inv_2 _429_ (
    .A(mprj_adr_o_core[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_024_)
  );
  sky130_fd_sc_hd__inv_2 _430_ (
    .A(mprj_adr_o_core[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_025_)
  );
  sky130_fd_sc_hd__inv_2 _431_ (
    .A(mprj_adr_o_core[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_026_)
  );
  sky130_fd_sc_hd__inv_2 _432_ (
    .A(mprj_adr_o_core[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_027_)
  );
  sky130_fd_sc_hd__inv_2 _433_ (
    .A(mprj_adr_o_core[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_028_)
  );
  sky130_fd_sc_hd__inv_2 _434_ (
    .A(mprj_adr_o_core[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_029_)
  );
  sky130_fd_sc_hd__inv_2 _435_ (
    .A(mprj_adr_o_core[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_030_)
  );
  sky130_fd_sc_hd__inv_2 _436_ (
    .A(mprj_adr_o_core[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_031_)
  );
  sky130_fd_sc_hd__inv_2 _437_ (
    .A(mprj_adr_o_core[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_033_)
  );
  sky130_fd_sc_hd__inv_2 _438_ (
    .A(mprj_adr_o_core[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_034_)
  );
  sky130_fd_sc_hd__inv_2 _439_ (
    .A(mprj_dat_o_core[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_042_)
  );
  sky130_fd_sc_hd__inv_2 _440_ (
    .A(mprj_dat_o_core[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_053_)
  );
  sky130_fd_sc_hd__inv_2 _441_ (
    .A(mprj_dat_o_core[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_064_)
  );
  sky130_fd_sc_hd__inv_2 _442_ (
    .A(mprj_dat_o_core[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_067_)
  );
  sky130_fd_sc_hd__inv_2 _443_ (
    .A(mprj_dat_o_core[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_068_)
  );
  sky130_fd_sc_hd__inv_2 _444_ (
    .A(mprj_dat_o_core[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_069_)
  );
  sky130_fd_sc_hd__inv_2 _445_ (
    .A(mprj_dat_o_core[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_070_)
  );
  sky130_fd_sc_hd__inv_2 _446_ (
    .A(mprj_dat_o_core[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_071_)
  );
  sky130_fd_sc_hd__inv_2 _447_ (
    .A(mprj_dat_o_core[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_072_)
  );
  sky130_fd_sc_hd__inv_2 _448_ (
    .A(mprj_dat_o_core[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_073_)
  );
  sky130_fd_sc_hd__inv_2 _449_ (
    .A(mprj_dat_o_core[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_043_)
  );
  sky130_fd_sc_hd__inv_2 _450_ (
    .A(mprj_dat_o_core[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_044_)
  );
  sky130_fd_sc_hd__inv_2 _451_ (
    .A(mprj_dat_o_core[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_045_)
  );
  sky130_fd_sc_hd__inv_2 _452_ (
    .A(mprj_dat_o_core[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_046_)
  );
  sky130_fd_sc_hd__inv_2 _453_ (
    .A(mprj_dat_o_core[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_047_)
  );
  sky130_fd_sc_hd__inv_2 _454_ (
    .A(mprj_dat_o_core[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_048_)
  );
  sky130_fd_sc_hd__inv_2 _455_ (
    .A(mprj_dat_o_core[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_049_)
  );
  sky130_fd_sc_hd__inv_2 _456_ (
    .A(mprj_dat_o_core[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_050_)
  );
  sky130_fd_sc_hd__inv_2 _457_ (
    .A(mprj_dat_o_core[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_051_)
  );
  sky130_fd_sc_hd__inv_2 _458_ (
    .A(mprj_dat_o_core[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_052_)
  );
  sky130_fd_sc_hd__inv_2 _459_ (
    .A(mprj_dat_o_core[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_054_)
  );
  sky130_fd_sc_hd__inv_2 _460_ (
    .A(mprj_dat_o_core[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_055_)
  );
  sky130_fd_sc_hd__inv_2 _461_ (
    .A(mprj_dat_o_core[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_056_)
  );
  sky130_fd_sc_hd__inv_2 _462_ (
    .A(mprj_dat_o_core[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_057_)
  );
  sky130_fd_sc_hd__inv_2 _463_ (
    .A(mprj_dat_o_core[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_058_)
  );
  sky130_fd_sc_hd__inv_2 _464_ (
    .A(mprj_dat_o_core[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_059_)
  );
  sky130_fd_sc_hd__inv_2 _465_ (
    .A(mprj_dat_o_core[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_060_)
  );
  sky130_fd_sc_hd__inv_2 _466_ (
    .A(mprj_dat_o_core[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_061_)
  );
  sky130_fd_sc_hd__inv_2 _467_ (
    .A(mprj_dat_o_core[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_062_)
  );
  sky130_fd_sc_hd__inv_2 _468_ (
    .A(mprj_dat_o_core[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_063_)
  );
  sky130_fd_sc_hd__inv_2 _469_ (
    .A(mprj_dat_o_core[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_065_)
  );
  sky130_fd_sc_hd__inv_2 _470_ (
    .A(mprj_dat_o_core[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_066_)
  );
  sky130_fd_sc_hd__inv_2 _471_ (
    .A(la_data_out_mprj[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_074_)
  );
  sky130_fd_sc_hd__inv_2 _472_ (
    .A(la_data_out_mprj[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_113_)
  );
  sky130_fd_sc_hd__inv_2 _473_ (
    .A(la_data_out_mprj[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_124_)
  );
  sky130_fd_sc_hd__inv_2 _474_ (
    .A(la_data_out_mprj[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_135_)
  );
  sky130_fd_sc_hd__inv_2 _475_ (
    .A(la_data_out_mprj[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_146_)
  );
  sky130_fd_sc_hd__inv_2 _476_ (
    .A(la_data_out_mprj[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_157_)
  );
  sky130_fd_sc_hd__inv_2 _477_ (
    .A(la_data_out_mprj[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_168_)
  );
  sky130_fd_sc_hd__inv_2 _478_ (
    .A(la_data_out_mprj[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_179_)
  );
  sky130_fd_sc_hd__inv_2 _479_ (
    .A(la_data_out_mprj[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_190_)
  );
  sky130_fd_sc_hd__inv_2 _480_ (
    .A(la_data_out_mprj[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_201_)
  );
  sky130_fd_sc_hd__inv_2 _481_ (
    .A(la_data_out_mprj[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_085_)
  );
  sky130_fd_sc_hd__inv_2 _482_ (
    .A(la_data_out_mprj[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_096_)
  );
  sky130_fd_sc_hd__inv_2 _483_ (
    .A(la_data_out_mprj[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_105_)
  );
  sky130_fd_sc_hd__inv_2 _484_ (
    .A(la_data_out_mprj[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_106_)
  );
  sky130_fd_sc_hd__inv_2 _485_ (
    .A(la_data_out_mprj[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_107_)
  );
  sky130_fd_sc_hd__inv_2 _486_ (
    .A(la_data_out_mprj[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_108_)
  );
  sky130_fd_sc_hd__inv_2 _487_ (
    .A(la_data_out_mprj[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_109_)
  );
  sky130_fd_sc_hd__inv_2 _488_ (
    .A(la_data_out_mprj[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_110_)
  );
  sky130_fd_sc_hd__inv_2 _489_ (
    .A(la_data_out_mprj[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_111_)
  );
  sky130_fd_sc_hd__inv_2 _490_ (
    .A(la_data_out_mprj[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_112_)
  );
  sky130_fd_sc_hd__inv_2 _491_ (
    .A(la_data_out_mprj[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_114_)
  );
  sky130_fd_sc_hd__inv_2 _492_ (
    .A(la_data_out_mprj[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_115_)
  );
  sky130_fd_sc_hd__inv_2 _493_ (
    .A(la_data_out_mprj[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_116_)
  );
  sky130_fd_sc_hd__inv_2 _494_ (
    .A(la_data_out_mprj[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_117_)
  );
  sky130_fd_sc_hd__inv_2 _495_ (
    .A(la_data_out_mprj[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_118_)
  );
  sky130_fd_sc_hd__inv_2 _496_ (
    .A(la_data_out_mprj[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_119_)
  );
  sky130_fd_sc_hd__inv_2 _497_ (
    .A(la_data_out_mprj[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_120_)
  );
  sky130_fd_sc_hd__inv_2 _498_ (
    .A(la_data_out_mprj[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_121_)
  );
  sky130_fd_sc_hd__inv_2 _499_ (
    .A(la_data_out_mprj[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_122_)
  );
  sky130_fd_sc_hd__inv_2 _500_ (
    .A(la_data_out_mprj[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_123_)
  );
  sky130_fd_sc_hd__inv_2 _501_ (
    .A(la_data_out_mprj[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_125_)
  );
  sky130_fd_sc_hd__inv_2 _502_ (
    .A(la_data_out_mprj[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_126_)
  );
  sky130_fd_sc_hd__inv_2 _503_ (
    .A(la_data_out_mprj[32]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_127_)
  );
  sky130_fd_sc_hd__inv_2 _504_ (
    .A(la_data_out_mprj[33]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_128_)
  );
  sky130_fd_sc_hd__inv_2 _505_ (
    .A(la_data_out_mprj[34]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_129_)
  );
  sky130_fd_sc_hd__inv_2 _506_ (
    .A(la_data_out_mprj[35]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_130_)
  );
  sky130_fd_sc_hd__inv_2 _507_ (
    .A(la_data_out_mprj[36]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_131_)
  );
  sky130_fd_sc_hd__inv_2 _508_ (
    .A(la_data_out_mprj[37]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_132_)
  );
  sky130_fd_sc_hd__inv_2 _509_ (
    .A(la_data_out_mprj[38]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_133_)
  );
  sky130_fd_sc_hd__inv_2 _510_ (
    .A(la_data_out_mprj[39]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_134_)
  );
  sky130_fd_sc_hd__inv_2 _511_ (
    .A(la_data_out_mprj[40]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_136_)
  );
  sky130_fd_sc_hd__inv_2 _512_ (
    .A(la_data_out_mprj[41]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_137_)
  );
  sky130_fd_sc_hd__inv_2 _513_ (
    .A(la_data_out_mprj[42]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_138_)
  );
  sky130_fd_sc_hd__inv_2 _514_ (
    .A(la_data_out_mprj[43]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_139_)
  );
  sky130_fd_sc_hd__inv_2 _515_ (
    .A(la_data_out_mprj[44]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_140_)
  );
  sky130_fd_sc_hd__inv_2 _516_ (
    .A(la_data_out_mprj[45]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_141_)
  );
  sky130_fd_sc_hd__inv_2 _517_ (
    .A(la_data_out_mprj[46]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_142_)
  );
  sky130_fd_sc_hd__inv_2 _518_ (
    .A(la_data_out_mprj[47]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_143_)
  );
  sky130_fd_sc_hd__inv_2 _519_ (
    .A(la_data_out_mprj[48]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_144_)
  );
  sky130_fd_sc_hd__inv_2 _520_ (
    .A(la_data_out_mprj[49]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_145_)
  );
  sky130_fd_sc_hd__inv_2 _521_ (
    .A(la_data_out_mprj[50]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_147_)
  );
  sky130_fd_sc_hd__inv_2 _522_ (
    .A(la_data_out_mprj[51]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_148_)
  );
  sky130_fd_sc_hd__inv_2 _523_ (
    .A(la_data_out_mprj[52]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_149_)
  );
  sky130_fd_sc_hd__inv_2 _524_ (
    .A(la_data_out_mprj[53]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_150_)
  );
  sky130_fd_sc_hd__inv_2 _525_ (
    .A(la_data_out_mprj[54]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_151_)
  );
  sky130_fd_sc_hd__inv_2 _526_ (
    .A(la_data_out_mprj[55]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_152_)
  );
  sky130_fd_sc_hd__inv_2 _527_ (
    .A(la_data_out_mprj[56]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_153_)
  );
  sky130_fd_sc_hd__inv_2 _528_ (
    .A(la_data_out_mprj[57]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_154_)
  );
  sky130_fd_sc_hd__inv_2 _529_ (
    .A(la_data_out_mprj[58]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_155_)
  );
  sky130_fd_sc_hd__inv_2 _530_ (
    .A(la_data_out_mprj[59]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_156_)
  );
  sky130_fd_sc_hd__inv_2 _531_ (
    .A(la_data_out_mprj[60]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_158_)
  );
  sky130_fd_sc_hd__inv_2 _532_ (
    .A(la_data_out_mprj[61]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_159_)
  );
  sky130_fd_sc_hd__inv_2 _533_ (
    .A(la_data_out_mprj[62]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_160_)
  );
  sky130_fd_sc_hd__inv_2 _534_ (
    .A(la_data_out_mprj[63]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_161_)
  );
  sky130_fd_sc_hd__inv_2 _535_ (
    .A(la_data_out_mprj[64]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_162_)
  );
  sky130_fd_sc_hd__inv_2 _536_ (
    .A(la_data_out_mprj[65]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_163_)
  );
  sky130_fd_sc_hd__inv_2 _537_ (
    .A(la_data_out_mprj[66]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_164_)
  );
  sky130_fd_sc_hd__inv_2 _538_ (
    .A(la_data_out_mprj[67]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_165_)
  );
  sky130_fd_sc_hd__inv_2 _539_ (
    .A(la_data_out_mprj[68]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_166_)
  );
  sky130_fd_sc_hd__inv_2 _540_ (
    .A(la_data_out_mprj[69]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_167_)
  );
  sky130_fd_sc_hd__inv_2 _541_ (
    .A(la_data_out_mprj[70]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_169_)
  );
  sky130_fd_sc_hd__inv_2 _542_ (
    .A(la_data_out_mprj[71]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_170_)
  );
  sky130_fd_sc_hd__inv_2 _543_ (
    .A(la_data_out_mprj[72]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_171_)
  );
  sky130_fd_sc_hd__inv_2 _544_ (
    .A(la_data_out_mprj[73]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_172_)
  );
  sky130_fd_sc_hd__inv_2 _545_ (
    .A(la_data_out_mprj[74]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_173_)
  );
  sky130_fd_sc_hd__inv_2 _546_ (
    .A(la_data_out_mprj[75]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_174_)
  );
  sky130_fd_sc_hd__inv_2 _547_ (
    .A(la_data_out_mprj[76]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_175_)
  );
  sky130_fd_sc_hd__inv_2 _548_ (
    .A(la_data_out_mprj[77]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_176_)
  );
  sky130_fd_sc_hd__inv_2 _549_ (
    .A(la_data_out_mprj[78]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_177_)
  );
  sky130_fd_sc_hd__inv_2 _550_ (
    .A(la_data_out_mprj[79]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_178_)
  );
  sky130_fd_sc_hd__inv_2 _551_ (
    .A(la_data_out_mprj[80]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_180_)
  );
  sky130_fd_sc_hd__inv_2 _552_ (
    .A(la_data_out_mprj[81]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_181_)
  );
  sky130_fd_sc_hd__inv_2 _553_ (
    .A(la_data_out_mprj[82]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_182_)
  );
  sky130_fd_sc_hd__inv_2 _554_ (
    .A(la_data_out_mprj[83]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_183_)
  );
  sky130_fd_sc_hd__inv_2 _555_ (
    .A(la_data_out_mprj[84]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_184_)
  );
  sky130_fd_sc_hd__inv_2 _556_ (
    .A(la_data_out_mprj[85]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_185_)
  );
  sky130_fd_sc_hd__inv_2 _557_ (
    .A(la_data_out_mprj[86]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_186_)
  );
  sky130_fd_sc_hd__inv_2 _558_ (
    .A(la_data_out_mprj[87]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_187_)
  );
  sky130_fd_sc_hd__inv_2 _559_ (
    .A(la_data_out_mprj[88]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_188_)
  );
  sky130_fd_sc_hd__inv_2 _560_ (
    .A(la_data_out_mprj[89]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_189_)
  );
  sky130_fd_sc_hd__inv_2 _561_ (
    .A(la_data_out_mprj[90]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_191_)
  );
  sky130_fd_sc_hd__inv_2 _562_ (
    .A(la_data_out_mprj[91]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_192_)
  );
  sky130_fd_sc_hd__inv_2 _563_ (
    .A(la_data_out_mprj[92]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_193_)
  );
  sky130_fd_sc_hd__inv_2 _564_ (
    .A(la_data_out_mprj[93]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_194_)
  );
  sky130_fd_sc_hd__inv_2 _565_ (
    .A(la_data_out_mprj[94]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_195_)
  );
  sky130_fd_sc_hd__inv_2 _566_ (
    .A(la_data_out_mprj[95]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_196_)
  );
  sky130_fd_sc_hd__inv_2 _567_ (
    .A(la_data_out_mprj[96]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_197_)
  );
  sky130_fd_sc_hd__inv_2 _568_ (
    .A(la_data_out_mprj[97]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_198_)
  );
  sky130_fd_sc_hd__inv_2 _569_ (
    .A(la_data_out_mprj[98]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_199_)
  );
  sky130_fd_sc_hd__inv_2 _570_ (
    .A(la_data_out_mprj[99]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_200_)
  );
  sky130_fd_sc_hd__inv_2 _571_ (
    .A(la_data_out_mprj[100]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_075_)
  );
  sky130_fd_sc_hd__inv_2 _572_ (
    .A(la_data_out_mprj[101]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_076_)
  );
  sky130_fd_sc_hd__inv_2 _573_ (
    .A(la_data_out_mprj[102]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_077_)
  );
  sky130_fd_sc_hd__inv_2 _574_ (
    .A(la_data_out_mprj[103]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_078_)
  );
  sky130_fd_sc_hd__inv_2 _575_ (
    .A(la_data_out_mprj[104]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_079_)
  );
  sky130_fd_sc_hd__inv_2 _576_ (
    .A(la_data_out_mprj[105]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_080_)
  );
  sky130_fd_sc_hd__inv_2 _577_ (
    .A(la_data_out_mprj[106]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_081_)
  );
  sky130_fd_sc_hd__inv_2 _578_ (
    .A(la_data_out_mprj[107]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_082_)
  );
  sky130_fd_sc_hd__inv_2 _579_ (
    .A(la_data_out_mprj[108]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_083_)
  );
  sky130_fd_sc_hd__inv_2 _580_ (
    .A(la_data_out_mprj[109]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_084_)
  );
  sky130_fd_sc_hd__inv_2 _581_ (
    .A(la_data_out_mprj[110]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_086_)
  );
  sky130_fd_sc_hd__inv_2 _582_ (
    .A(la_data_out_mprj[111]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_087_)
  );
  sky130_fd_sc_hd__inv_2 _583_ (
    .A(la_data_out_mprj[112]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_088_)
  );
  sky130_fd_sc_hd__inv_2 _584_ (
    .A(la_data_out_mprj[113]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_089_)
  );
  sky130_fd_sc_hd__inv_2 _585_ (
    .A(la_data_out_mprj[114]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_090_)
  );
  sky130_fd_sc_hd__inv_2 _586_ (
    .A(la_data_out_mprj[115]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_091_)
  );
  sky130_fd_sc_hd__inv_2 _587_ (
    .A(la_data_out_mprj[116]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_092_)
  );
  sky130_fd_sc_hd__inv_2 _588_ (
    .A(la_data_out_mprj[117]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_093_)
  );
  sky130_fd_sc_hd__inv_2 _589_ (
    .A(la_data_out_mprj[118]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_094_)
  );
  sky130_fd_sc_hd__inv_2 _590_ (
    .A(la_data_out_mprj[119]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_095_)
  );
  sky130_fd_sc_hd__inv_2 _591_ (
    .A(la_data_out_mprj[120]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_097_)
  );
  sky130_fd_sc_hd__inv_2 _592_ (
    .A(la_data_out_mprj[121]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_098_)
  );
  sky130_fd_sc_hd__inv_2 _593_ (
    .A(la_data_out_mprj[122]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_099_)
  );
  sky130_fd_sc_hd__inv_2 _594_ (
    .A(la_data_out_mprj[123]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_100_)
  );
  sky130_fd_sc_hd__inv_2 _595_ (
    .A(la_data_out_mprj[124]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_101_)
  );
  sky130_fd_sc_hd__inv_2 _596_ (
    .A(la_data_out_mprj[125]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_102_)
  );
  sky130_fd_sc_hd__inv_2 _597_ (
    .A(la_data_out_mprj[126]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_103_)
  );
  sky130_fd_sc_hd__inv_2 _598_ (
    .A(la_data_out_mprj[127]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_104_)
  );
  sky130_fd_sc_hd__inv_2 _599_ (
    .A(la_oen_mprj[0]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_202_)
  );
  sky130_fd_sc_hd__inv_2 _600_ (
    .A(la_oen_mprj[1]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_241_)
  );
  sky130_fd_sc_hd__inv_2 _601_ (
    .A(la_oen_mprj[2]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_252_)
  );
  sky130_fd_sc_hd__inv_2 _602_ (
    .A(la_oen_mprj[3]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_263_)
  );
  sky130_fd_sc_hd__inv_2 _603_ (
    .A(la_oen_mprj[4]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_274_)
  );
  sky130_fd_sc_hd__inv_2 _604_ (
    .A(la_oen_mprj[5]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_285_)
  );
  sky130_fd_sc_hd__inv_2 _605_ (
    .A(la_oen_mprj[6]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_296_)
  );
  sky130_fd_sc_hd__inv_2 _606_ (
    .A(la_oen_mprj[7]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_307_)
  );
  sky130_fd_sc_hd__inv_2 _607_ (
    .A(la_oen_mprj[8]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_318_)
  );
  sky130_fd_sc_hd__inv_2 _608_ (
    .A(la_oen_mprj[9]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_329_)
  );
  sky130_fd_sc_hd__inv_2 _609_ (
    .A(la_oen_mprj[10]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_213_)
  );
  sky130_fd_sc_hd__inv_2 _610_ (
    .A(la_oen_mprj[11]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_224_)
  );
  sky130_fd_sc_hd__inv_2 _611_ (
    .A(la_oen_mprj[12]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_233_)
  );
  sky130_fd_sc_hd__inv_2 _612_ (
    .A(la_oen_mprj[13]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_234_)
  );
  sky130_fd_sc_hd__inv_2 _613_ (
    .A(la_oen_mprj[14]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_235_)
  );
  sky130_fd_sc_hd__inv_2 _614_ (
    .A(la_oen_mprj[15]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_236_)
  );
  sky130_fd_sc_hd__inv_2 _615_ (
    .A(la_oen_mprj[16]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_237_)
  );
  sky130_fd_sc_hd__inv_2 _616_ (
    .A(la_oen_mprj[17]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_238_)
  );
  sky130_fd_sc_hd__inv_2 _617_ (
    .A(la_oen_mprj[18]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_239_)
  );
  sky130_fd_sc_hd__inv_2 _618_ (
    .A(la_oen_mprj[19]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_240_)
  );
  sky130_fd_sc_hd__inv_2 _619_ (
    .A(la_oen_mprj[20]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_242_)
  );
  sky130_fd_sc_hd__inv_2 _620_ (
    .A(la_oen_mprj[21]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_243_)
  );
  sky130_fd_sc_hd__inv_2 _621_ (
    .A(la_oen_mprj[22]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_244_)
  );
  sky130_fd_sc_hd__inv_2 _622_ (
    .A(la_oen_mprj[23]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_245_)
  );
  sky130_fd_sc_hd__inv_2 _623_ (
    .A(la_oen_mprj[24]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_246_)
  );
  sky130_fd_sc_hd__inv_2 _624_ (
    .A(la_oen_mprj[25]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_247_)
  );
  sky130_fd_sc_hd__inv_2 _625_ (
    .A(la_oen_mprj[26]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_248_)
  );
  sky130_fd_sc_hd__inv_2 _626_ (
    .A(la_oen_mprj[27]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_249_)
  );
  sky130_fd_sc_hd__inv_2 _627_ (
    .A(la_oen_mprj[28]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_250_)
  );
  sky130_fd_sc_hd__inv_2 _628_ (
    .A(la_oen_mprj[29]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_251_)
  );
  sky130_fd_sc_hd__inv_2 _629_ (
    .A(la_oen_mprj[30]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_253_)
  );
  sky130_fd_sc_hd__inv_2 _630_ (
    .A(la_oen_mprj[31]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_254_)
  );
  sky130_fd_sc_hd__inv_2 _631_ (
    .A(la_oen_mprj[32]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_255_)
  );
  sky130_fd_sc_hd__inv_2 _632_ (
    .A(la_oen_mprj[33]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_256_)
  );
  sky130_fd_sc_hd__inv_2 _633_ (
    .A(la_oen_mprj[34]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_257_)
  );
  sky130_fd_sc_hd__inv_2 _634_ (
    .A(la_oen_mprj[35]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_258_)
  );
  sky130_fd_sc_hd__inv_2 _635_ (
    .A(la_oen_mprj[36]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_259_)
  );
  sky130_fd_sc_hd__inv_2 _636_ (
    .A(la_oen_mprj[37]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_260_)
  );
  sky130_fd_sc_hd__inv_2 _637_ (
    .A(la_oen_mprj[38]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_261_)
  );
  sky130_fd_sc_hd__inv_2 _638_ (
    .A(la_oen_mprj[39]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_262_)
  );
  sky130_fd_sc_hd__inv_2 _639_ (
    .A(la_oen_mprj[40]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_264_)
  );
  sky130_fd_sc_hd__inv_2 _640_ (
    .A(la_oen_mprj[41]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_265_)
  );
  sky130_fd_sc_hd__inv_2 _641_ (
    .A(la_oen_mprj[42]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_266_)
  );
  sky130_fd_sc_hd__inv_2 _642_ (
    .A(la_oen_mprj[43]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_267_)
  );
  sky130_fd_sc_hd__inv_2 _643_ (
    .A(la_oen_mprj[44]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_268_)
  );
  sky130_fd_sc_hd__inv_2 _644_ (
    .A(la_oen_mprj[45]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_269_)
  );
  sky130_fd_sc_hd__inv_2 _645_ (
    .A(la_oen_mprj[46]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_270_)
  );
  sky130_fd_sc_hd__inv_2 _646_ (
    .A(la_oen_mprj[47]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_271_)
  );
  sky130_fd_sc_hd__inv_2 _647_ (
    .A(la_oen_mprj[48]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_272_)
  );
  sky130_fd_sc_hd__inv_2 _648_ (
    .A(la_oen_mprj[49]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_273_)
  );
  sky130_fd_sc_hd__inv_2 _649_ (
    .A(la_oen_mprj[50]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_275_)
  );
  sky130_fd_sc_hd__inv_2 _650_ (
    .A(la_oen_mprj[51]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_276_)
  );
  sky130_fd_sc_hd__inv_2 _651_ (
    .A(la_oen_mprj[52]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_277_)
  );
  sky130_fd_sc_hd__inv_2 _652_ (
    .A(la_oen_mprj[53]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_278_)
  );
  sky130_fd_sc_hd__inv_2 _653_ (
    .A(la_oen_mprj[54]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_279_)
  );
  sky130_fd_sc_hd__inv_2 _654_ (
    .A(la_oen_mprj[55]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_280_)
  );
  sky130_fd_sc_hd__inv_2 _655_ (
    .A(la_oen_mprj[56]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_281_)
  );
  sky130_fd_sc_hd__inv_2 _656_ (
    .A(la_oen_mprj[57]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_282_)
  );
  sky130_fd_sc_hd__inv_2 _657_ (
    .A(la_oen_mprj[58]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_283_)
  );
  sky130_fd_sc_hd__inv_2 _658_ (
    .A(la_oen_mprj[59]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_284_)
  );
  sky130_fd_sc_hd__inv_2 _659_ (
    .A(la_oen_mprj[60]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_286_)
  );
  sky130_fd_sc_hd__inv_2 _660_ (
    .A(la_oen_mprj[61]),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(_287_)
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[0]  (
    .A(_074_),
    .TE(\mprj_logic1[74] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[0])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[100]  (
    .A(_075_),
    .TE(\mprj_logic1[174] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[100])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[101]  (
    .A(_076_),
    .TE(\mprj_logic1[175] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[101])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[102]  (
    .A(_077_),
    .TE(\mprj_logic1[176] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[102])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[103]  (
    .A(_078_),
    .TE(\mprj_logic1[177] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[103])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[104]  (
    .A(_079_),
    .TE(\mprj_logic1[178] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[104])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[105]  (
    .A(_080_),
    .TE(\mprj_logic1[179] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[105])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[106]  (
    .A(_081_),
    .TE(\mprj_logic1[180] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[106])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[107]  (
    .A(_082_),
    .TE(\mprj_logic1[181] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[107])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[108]  (
    .A(_083_),
    .TE(\mprj_logic1[182] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[108])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[109]  (
    .A(_084_),
    .TE(\mprj_logic1[183] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[109])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[10]  (
    .A(_085_),
    .TE(\mprj_logic1[84] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[10])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[110]  (
    .A(_086_),
    .TE(\mprj_logic1[184] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[110])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[111]  (
    .A(_087_),
    .TE(\mprj_logic1[185] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[111])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[112]  (
    .A(_088_),
    .TE(\mprj_logic1[186] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[112])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[113]  (
    .A(_089_),
    .TE(\mprj_logic1[187] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[113])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[114]  (
    .A(_090_),
    .TE(\mprj_logic1[188] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[114])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[115]  (
    .A(_091_),
    .TE(\mprj_logic1[189] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[115])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[116]  (
    .A(_092_),
    .TE(\mprj_logic1[190] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[116])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[117]  (
    .A(_093_),
    .TE(\mprj_logic1[191] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[117])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[118]  (
    .A(_094_),
    .TE(\mprj_logic1[192] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[118])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[119]  (
    .A(_095_),
    .TE(\mprj_logic1[193] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[119])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[11]  (
    .A(_096_),
    .TE(\mprj_logic1[85] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[11])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[120]  (
    .A(_097_),
    .TE(\mprj_logic1[194] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[120])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[121]  (
    .A(_098_),
    .TE(\mprj_logic1[195] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[121])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[122]  (
    .A(_099_),
    .TE(\mprj_logic1[196] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[122])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[123]  (
    .A(_100_),
    .TE(\mprj_logic1[197] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[123])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[124]  (
    .A(_101_),
    .TE(\mprj_logic1[198] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[124])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[125]  (
    .A(_102_),
    .TE(\mprj_logic1[199] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[125])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[126]  (
    .A(_103_),
    .TE(\mprj_logic1[200] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[126])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[127]  (
    .A(_104_),
    .TE(\mprj_logic1[201] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[127])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[12]  (
    .A(_105_),
    .TE(\mprj_logic1[86] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[12])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[13]  (
    .A(_106_),
    .TE(\mprj_logic1[87] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[13])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[14]  (
    .A(_107_),
    .TE(\mprj_logic1[88] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[14])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[15]  (
    .A(_108_),
    .TE(\mprj_logic1[89] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[15])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[16]  (
    .A(_109_),
    .TE(\mprj_logic1[90] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[16])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[17]  (
    .A(_110_),
    .TE(\mprj_logic1[91] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[17])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[18]  (
    .A(_111_),
    .TE(\mprj_logic1[92] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[18])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[19]  (
    .A(_112_),
    .TE(\mprj_logic1[93] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[19])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[1]  (
    .A(_113_),
    .TE(\mprj_logic1[75] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[1])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[20]  (
    .A(_114_),
    .TE(\mprj_logic1[94] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[20])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[21]  (
    .A(_115_),
    .TE(\mprj_logic1[95] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[21])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[22]  (
    .A(_116_),
    .TE(\mprj_logic1[96] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[22])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[23]  (
    .A(_117_),
    .TE(\mprj_logic1[97] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[23])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[24]  (
    .A(_118_),
    .TE(\mprj_logic1[98] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[24])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[25]  (
    .A(_119_),
    .TE(\mprj_logic1[99] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[25])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[26]  (
    .A(_120_),
    .TE(\mprj_logic1[100] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[26])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[27]  (
    .A(_121_),
    .TE(\mprj_logic1[101] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[27])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[28]  (
    .A(_122_),
    .TE(\mprj_logic1[102] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[28])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[29]  (
    .A(_123_),
    .TE(\mprj_logic1[103] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[29])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[2]  (
    .A(_124_),
    .TE(\mprj_logic1[76] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[2])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[30]  (
    .A(_125_),
    .TE(\mprj_logic1[104] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[30])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[31]  (
    .A(_126_),
    .TE(\mprj_logic1[105] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[31])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[32]  (
    .A(_127_),
    .TE(\mprj_logic1[106] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[32])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[33]  (
    .A(_128_),
    .TE(\mprj_logic1[107] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[33])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[34]  (
    .A(_129_),
    .TE(\mprj_logic1[108] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[34])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[35]  (
    .A(_130_),
    .TE(\mprj_logic1[109] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[35])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[36]  (
    .A(_131_),
    .TE(\mprj_logic1[110] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[36])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[37]  (
    .A(_132_),
    .TE(\mprj_logic1[111] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[37])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[38]  (
    .A(_133_),
    .TE(\mprj_logic1[112] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[38])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[39]  (
    .A(_134_),
    .TE(\mprj_logic1[113] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[39])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[3]  (
    .A(_135_),
    .TE(\mprj_logic1[77] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[3])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[40]  (
    .A(_136_),
    .TE(\mprj_logic1[114] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[40])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[41]  (
    .A(_137_),
    .TE(\mprj_logic1[115] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[41])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[42]  (
    .A(_138_),
    .TE(\mprj_logic1[116] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[42])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[43]  (
    .A(_139_),
    .TE(\mprj_logic1[117] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[43])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[44]  (
    .A(_140_),
    .TE(\mprj_logic1[118] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[44])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[45]  (
    .A(_141_),
    .TE(\mprj_logic1[119] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[45])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[46]  (
    .A(_142_),
    .TE(\mprj_logic1[120] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[46])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[47]  (
    .A(_143_),
    .TE(\mprj_logic1[121] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[47])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[48]  (
    .A(_144_),
    .TE(\mprj_logic1[122] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[48])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[49]  (
    .A(_145_),
    .TE(\mprj_logic1[123] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[49])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[4]  (
    .A(_146_),
    .TE(\mprj_logic1[78] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[4])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[50]  (
    .A(_147_),
    .TE(\mprj_logic1[124] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[50])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[51]  (
    .A(_148_),
    .TE(\mprj_logic1[125] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[51])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[52]  (
    .A(_149_),
    .TE(\mprj_logic1[126] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[52])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[53]  (
    .A(_150_),
    .TE(\mprj_logic1[127] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[53])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[54]  (
    .A(_151_),
    .TE(\mprj_logic1[128] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[54])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[55]  (
    .A(_152_),
    .TE(\mprj_logic1[129] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[55])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[56]  (
    .A(_153_),
    .TE(\mprj_logic1[130] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[56])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[57]  (
    .A(_154_),
    .TE(\mprj_logic1[131] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[57])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[58]  (
    .A(_155_),
    .TE(\mprj_logic1[132] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[58])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[59]  (
    .A(_156_),
    .TE(\mprj_logic1[133] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[59])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[5]  (
    .A(_157_),
    .TE(\mprj_logic1[79] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[5])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[60]  (
    .A(_158_),
    .TE(\mprj_logic1[134] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[60])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[61]  (
    .A(_159_),
    .TE(\mprj_logic1[135] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[61])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[62]  (
    .A(_160_),
    .TE(\mprj_logic1[136] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[62])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[63]  (
    .A(_161_),
    .TE(\mprj_logic1[137] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[63])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[64]  (
    .A(_162_),
    .TE(\mprj_logic1[138] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[64])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[65]  (
    .A(_163_),
    .TE(\mprj_logic1[139] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[65])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[66]  (
    .A(_164_),
    .TE(\mprj_logic1[140] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[66])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[67]  (
    .A(_165_),
    .TE(\mprj_logic1[141] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[67])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[68]  (
    .A(_166_),
    .TE(\mprj_logic1[142] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[68])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[69]  (
    .A(_167_),
    .TE(\mprj_logic1[143] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[69])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[6]  (
    .A(_168_),
    .TE(\mprj_logic1[80] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[6])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[70]  (
    .A(_169_),
    .TE(\mprj_logic1[144] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[70])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[71]  (
    .A(_170_),
    .TE(\mprj_logic1[145] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[71])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[72]  (
    .A(_171_),
    .TE(\mprj_logic1[146] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[72])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[73]  (
    .A(_172_),
    .TE(\mprj_logic1[147] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[73])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[74]  (
    .A(_173_),
    .TE(\mprj_logic1[148] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[74])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[75]  (
    .A(_174_),
    .TE(\mprj_logic1[149] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[75])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[76]  (
    .A(_175_),
    .TE(\mprj_logic1[150] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[76])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[77]  (
    .A(_176_),
    .TE(\mprj_logic1[151] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[77])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[78]  (
    .A(_177_),
    .TE(\mprj_logic1[152] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[78])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[79]  (
    .A(_178_),
    .TE(\mprj_logic1[153] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[79])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[7]  (
    .A(_179_),
    .TE(\mprj_logic1[81] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[7])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[80]  (
    .A(_180_),
    .TE(\mprj_logic1[154] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[80])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[81]  (
    .A(_181_),
    .TE(\mprj_logic1[155] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[81])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[82]  (
    .A(_182_),
    .TE(\mprj_logic1[156] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[82])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[83]  (
    .A(_183_),
    .TE(\mprj_logic1[157] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[83])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[84]  (
    .A(_184_),
    .TE(\mprj_logic1[158] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[84])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[85]  (
    .A(_185_),
    .TE(\mprj_logic1[159] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[85])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[86]  (
    .A(_186_),
    .TE(\mprj_logic1[160] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[86])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[87]  (
    .A(_187_),
    .TE(\mprj_logic1[161] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[87])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[88]  (
    .A(_188_),
    .TE(\mprj_logic1[162] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[88])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[89]  (
    .A(_189_),
    .TE(\mprj_logic1[163] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[89])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[8]  (
    .A(_190_),
    .TE(\mprj_logic1[82] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[8])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[90]  (
    .A(_191_),
    .TE(\mprj_logic1[164] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[90])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[91]  (
    .A(_192_),
    .TE(\mprj_logic1[165] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[91])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[92]  (
    .A(_193_),
    .TE(\mprj_logic1[166] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[92])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[93]  (
    .A(_194_),
    .TE(\mprj_logic1[167] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[93])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[94]  (
    .A(_195_),
    .TE(\mprj_logic1[168] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[94])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[95]  (
    .A(_196_),
    .TE(\mprj_logic1[169] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[95])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[96]  (
    .A(_197_),
    .TE(\mprj_logic1[170] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[96])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[97]  (
    .A(_198_),
    .TE(\mprj_logic1[171] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[97])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[98]  (
    .A(_199_),
    .TE(\mprj_logic1[172] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[98])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[99]  (
    .A(_200_),
    .TE(\mprj_logic1[173] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[99])
  );
  sky130_fd_sc_hd__einvp_8 \la_buf[9]  (
    .A(_201_),
    .TE(\mprj_logic1[83] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_data_in_core[9])
  );
  mprj2_logic_high mprj2_logic_high_inst (
    .HI(mprj2_logic1),
    .vccd2(vccd2),
    .vssd2(vssd2)
  );
  sky130_fd_sc_hd__buf_8 mprj2_pwrgood (
    .A(mprj2_logic1),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .X(user2_vcc_powergood)
  );
  sky130_fd_sc_hd__buf_8 mprj2_vdd_pwrgood (
    .A(mprj2_vdd_logic1),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .X(user2_vdd_powergood)
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[0]  (
    .A(_010_),
    .TE(\mprj_logic1[10] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[0])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[10]  (
    .A(_011_),
    .TE(\mprj_logic1[20] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[10])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[11]  (
    .A(_012_),
    .TE(\mprj_logic1[21] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[11])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[12]  (
    .A(_013_),
    .TE(\mprj_logic1[22] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[12])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[13]  (
    .A(_014_),
    .TE(\mprj_logic1[23] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[13])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[14]  (
    .A(_015_),
    .TE(\mprj_logic1[24] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[14])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[15]  (
    .A(_016_),
    .TE(\mprj_logic1[25] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[15])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[16]  (
    .A(_017_),
    .TE(\mprj_logic1[26] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[16])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[17]  (
    .A(_018_),
    .TE(\mprj_logic1[27] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[17])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[18]  (
    .A(_019_),
    .TE(\mprj_logic1[28] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[18])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[19]  (
    .A(_020_),
    .TE(\mprj_logic1[29] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[19])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[1]  (
    .A(_021_),
    .TE(\mprj_logic1[11] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[1])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[20]  (
    .A(_022_),
    .TE(\mprj_logic1[30] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[20])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[21]  (
    .A(_023_),
    .TE(\mprj_logic1[31] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[21])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[22]  (
    .A(_024_),
    .TE(\mprj_logic1[32] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[22])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[23]  (
    .A(_025_),
    .TE(\mprj_logic1[33] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[23])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[24]  (
    .A(_026_),
    .TE(\mprj_logic1[34] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[24])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[25]  (
    .A(_027_),
    .TE(\mprj_logic1[35] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[25])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[26]  (
    .A(_028_),
    .TE(\mprj_logic1[36] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[26])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[27]  (
    .A(_029_),
    .TE(\mprj_logic1[37] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[27])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[28]  (
    .A(_030_),
    .TE(\mprj_logic1[38] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[28])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[29]  (
    .A(_031_),
    .TE(\mprj_logic1[39] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[29])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[2]  (
    .A(_032_),
    .TE(\mprj_logic1[12] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[2])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[30]  (
    .A(_033_),
    .TE(\mprj_logic1[40] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[30])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[31]  (
    .A(_034_),
    .TE(\mprj_logic1[41] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[31])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[3]  (
    .A(_035_),
    .TE(\mprj_logic1[13] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[3])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[4]  (
    .A(_036_),
    .TE(\mprj_logic1[14] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[4])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[5]  (
    .A(_037_),
    .TE(\mprj_logic1[15] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[5])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[6]  (
    .A(_038_),
    .TE(\mprj_logic1[16] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[6])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[7]  (
    .A(_039_),
    .TE(\mprj_logic1[17] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[7])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[8]  (
    .A(_040_),
    .TE(\mprj_logic1[18] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[8])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_adr_buf[9]  (
    .A(_041_),
    .TE(\mprj_logic1[19] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_adr_o_user[9])
  );
  sky130_fd_sc_hd__einvp_8 mprj_clk2_buf (
    .A(_002_),
    .TE(\mprj_logic1[2] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(user_clock2)
  );
  sky130_fd_sc_hd__einvp_8 mprj_clk_buf (
    .A(_001_),
    .TE(\mprj_logic1[1] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(user_clock)
  );
  sky130_fd_sc_hd__einvp_8 mprj_cyc_buf (
    .A(_003_),
    .TE(\mprj_logic1[3] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_cyc_o_user)
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[0]  (
    .A(_042_),
    .TE(\mprj_logic1[42] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[0])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[10]  (
    .A(_043_),
    .TE(\mprj_logic1[52] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[10])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[11]  (
    .A(_044_),
    .TE(\mprj_logic1[53] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[11])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[12]  (
    .A(_045_),
    .TE(\mprj_logic1[54] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[12])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[13]  (
    .A(_046_),
    .TE(\mprj_logic1[55] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[13])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[14]  (
    .A(_047_),
    .TE(\mprj_logic1[56] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[14])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[15]  (
    .A(_048_),
    .TE(\mprj_logic1[57] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[15])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[16]  (
    .A(_049_),
    .TE(\mprj_logic1[58] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[16])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[17]  (
    .A(_050_),
    .TE(\mprj_logic1[59] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[17])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[18]  (
    .A(_051_),
    .TE(\mprj_logic1[60] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[18])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[19]  (
    .A(_052_),
    .TE(\mprj_logic1[61] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[19])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[1]  (
    .A(_053_),
    .TE(\mprj_logic1[43] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[1])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[20]  (
    .A(_054_),
    .TE(\mprj_logic1[62] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[20])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[21]  (
    .A(_055_),
    .TE(\mprj_logic1[63] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[21])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[22]  (
    .A(_056_),
    .TE(\mprj_logic1[64] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[22])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[23]  (
    .A(_057_),
    .TE(\mprj_logic1[65] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[23])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[24]  (
    .A(_058_),
    .TE(\mprj_logic1[66] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[24])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[25]  (
    .A(_059_),
    .TE(\mprj_logic1[67] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[25])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[26]  (
    .A(_060_),
    .TE(\mprj_logic1[68] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[26])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[27]  (
    .A(_061_),
    .TE(\mprj_logic1[69] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[27])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[28]  (
    .A(_062_),
    .TE(\mprj_logic1[70] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[28])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[29]  (
    .A(_063_),
    .TE(\mprj_logic1[71] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[29])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[2]  (
    .A(_064_),
    .TE(\mprj_logic1[44] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[2])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[30]  (
    .A(_065_),
    .TE(\mprj_logic1[72] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[30])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[31]  (
    .A(_066_),
    .TE(\mprj_logic1[73] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[31])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[3]  (
    .A(_067_),
    .TE(\mprj_logic1[45] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[3])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[4]  (
    .A(_068_),
    .TE(\mprj_logic1[46] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[4])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[5]  (
    .A(_069_),
    .TE(\mprj_logic1[47] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[5])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[6]  (
    .A(_070_),
    .TE(\mprj_logic1[48] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[6])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[7]  (
    .A(_071_),
    .TE(\mprj_logic1[49] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[7])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[8]  (
    .A(_072_),
    .TE(\mprj_logic1[50] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[8])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_dat_buf[9]  (
    .A(_073_),
    .TE(\mprj_logic1[51] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_dat_o_user[9])
  );
  mprj_logic_high mprj_logic_high_inst (
    .HI({ \mprj_logic1[458] , \mprj_logic1[457] , \mprj_logic1[456] , \mprj_logic1[455] , \mprj_logic1[454] , \mprj_logic1[453] , \mprj_logic1[452] , \mprj_logic1[451] , \mprj_logic1[450] , \mprj_logic1[449] , \mprj_logic1[448] , \mprj_logic1[447] , \mprj_logic1[446] , \mprj_logic1[445] , \mprj_logic1[444] , \mprj_logic1[443] , \mprj_logic1[442] , \mprj_logic1[441] , \mprj_logic1[440] , \mprj_logic1[439] , \mprj_logic1[438] , \mprj_logic1[437] , \mprj_logic1[436] , \mprj_logic1[435] , \mprj_logic1[434] , \mprj_logic1[433] , \mprj_logic1[432] , \mprj_logic1[431] , \mprj_logic1[430] , \mprj_logic1[429] , \mprj_logic1[428] , \mprj_logic1[427] , \mprj_logic1[426] , \mprj_logic1[425] , \mprj_logic1[424] , \mprj_logic1[423] , \mprj_logic1[422] , \mprj_logic1[421] , \mprj_logic1[420] , \mprj_logic1[419] , \mprj_logic1[418] , \mprj_logic1[417] , \mprj_logic1[416] , \mprj_logic1[415] , \mprj_logic1[414] , \mprj_logic1[413] , \mprj_logic1[412] , \mprj_logic1[411] , \mprj_logic1[410] , \mprj_logic1[409] , \mprj_logic1[408] , \mprj_logic1[407] , \mprj_logic1[406] , \mprj_logic1[405] , \mprj_logic1[404] , \mprj_logic1[403] , \mprj_logic1[402] , \mprj_logic1[401] , \mprj_logic1[400] , \mprj_logic1[399] , \mprj_logic1[398] , \mprj_logic1[397] , \mprj_logic1[396] , \mprj_logic1[395] , \mprj_logic1[394] , \mprj_logic1[393] , \mprj_logic1[392] , \mprj_logic1[391] , \mprj_logic1[390] , \mprj_logic1[389] , \mprj_logic1[388] , \mprj_logic1[387] , \mprj_logic1[386] , \mprj_logic1[385] , \mprj_logic1[384] , \mprj_logic1[383] , \mprj_logic1[382] , \mprj_logic1[381] , \mprj_logic1[380] , \mprj_logic1[379] , \mprj_logic1[378] , \mprj_logic1[377] , \mprj_logic1[376] , \mprj_logic1[375] , \mprj_logic1[374] , \mprj_logic1[373] , \mprj_logic1[372] , \mprj_logic1[371] , \mprj_logic1[370] , \mprj_logic1[369] , \mprj_logic1[368] , \mprj_logic1[367] , \mprj_logic1[366] , \mprj_logic1[365] , \mprj_logic1[364] , \mprj_logic1[363] , \mprj_logic1[362] , \mprj_logic1[361] , \mprj_logic1[360] , \mprj_logic1[359] , \mprj_logic1[358] , \mprj_logic1[357] , \mprj_logic1[356] , \mprj_logic1[355] , \mprj_logic1[354] , \mprj_logic1[353] , \mprj_logic1[352] , \mprj_logic1[351] , \mprj_logic1[350] , \mprj_logic1[349] , \mprj_logic1[348] , \mprj_logic1[347] , \mprj_logic1[346] , \mprj_logic1[345] , \mprj_logic1[344] , \mprj_logic1[343] , \mprj_logic1[342] , \mprj_logic1[341] , \mprj_logic1[340] , \mprj_logic1[339] , \mprj_logic1[338] , \mprj_logic1[337] , \mprj_logic1[336] , \mprj_logic1[335] , \mprj_logic1[334] , \mprj_logic1[333] , \mprj_logic1[332] , \mprj_logic1[331] , \mprj_logic1[330] , \mprj_logic1[329] , \mprj_logic1[328] , \mprj_logic1[327] , \mprj_logic1[326] , \mprj_logic1[325] , \mprj_logic1[324] , \mprj_logic1[323] , \mprj_logic1[322] , \mprj_logic1[321] , \mprj_logic1[320] , \mprj_logic1[319] , \mprj_logic1[318] , \mprj_logic1[317] , \mprj_logic1[316] , \mprj_logic1[315] , \mprj_logic1[314] , \mprj_logic1[313] , \mprj_logic1[312] , \mprj_logic1[311] , \mprj_logic1[310] , \mprj_logic1[309] , \mprj_logic1[308] , \mprj_logic1[307] , \mprj_logic1[306] , \mprj_logic1[305] , \mprj_logic1[304] , \mprj_logic1[303] , \mprj_logic1[302] , \mprj_logic1[301] , \mprj_logic1[300] , \mprj_logic1[299] , \mprj_logic1[298] , \mprj_logic1[297] , \mprj_logic1[296] , \mprj_logic1[295] , \mprj_logic1[294] , \mprj_logic1[293] , \mprj_logic1[292] , \mprj_logic1[291] , \mprj_logic1[290] , \mprj_logic1[289] , \mprj_logic1[288] , \mprj_logic1[287] , \mprj_logic1[286] , \mprj_logic1[285] , \mprj_logic1[284] , \mprj_logic1[283] , \mprj_logic1[282] , \mprj_logic1[281] , \mprj_logic1[280] , \mprj_logic1[279] , \mprj_logic1[278] , \mprj_logic1[277] , \mprj_logic1[276] , \mprj_logic1[275] , \mprj_logic1[274] , \mprj_logic1[273] , \mprj_logic1[272] , \mprj_logic1[271] , \mprj_logic1[270] , \mprj_logic1[269] , \mprj_logic1[268] , \mprj_logic1[267] , \mprj_logic1[266] , \mprj_logic1[265] , \mprj_logic1[264] , \mprj_logic1[263] , \mprj_logic1[262] , \mprj_logic1[261] , \mprj_logic1[260] , \mprj_logic1[259] , \mprj_logic1[258] , \mprj_logic1[257] , \mprj_logic1[256] , \mprj_logic1[255] , \mprj_logic1[254] , \mprj_logic1[253] , \mprj_logic1[252] , \mprj_logic1[251] , \mprj_logic1[250] , \mprj_logic1[249] , \mprj_logic1[248] , \mprj_logic1[247] , \mprj_logic1[246] , \mprj_logic1[245] , \mprj_logic1[244] , \mprj_logic1[243] , \mprj_logic1[242] , \mprj_logic1[241] , \mprj_logic1[240] , \mprj_logic1[239] , \mprj_logic1[238] , \mprj_logic1[237] , \mprj_logic1[236] , \mprj_logic1[235] , \mprj_logic1[234] , \mprj_logic1[233] , \mprj_logic1[232] , \mprj_logic1[231] , \mprj_logic1[230] , \mprj_logic1[229] , \mprj_logic1[228] , \mprj_logic1[227] , \mprj_logic1[226] , \mprj_logic1[225] , \mprj_logic1[224] , \mprj_logic1[223] , \mprj_logic1[222] , \mprj_logic1[221] , \mprj_logic1[220] , \mprj_logic1[219] , \mprj_logic1[218] , \mprj_logic1[217] , \mprj_logic1[216] , \mprj_logic1[215] , \mprj_logic1[214] , \mprj_logic1[213] , \mprj_logic1[212] , \mprj_logic1[211] , \mprj_logic1[210] , \mprj_logic1[209] , \mprj_logic1[208] , \mprj_logic1[207] , \mprj_logic1[206] , \mprj_logic1[205] , \mprj_logic1[204] , \mprj_logic1[203] , \mprj_logic1[202] , \mprj_logic1[201] , \mprj_logic1[200] , \mprj_logic1[199] , \mprj_logic1[198] , \mprj_logic1[197] , \mprj_logic1[196] , \mprj_logic1[195] , \mprj_logic1[194] , \mprj_logic1[193] , \mprj_logic1[192] , \mprj_logic1[191] , \mprj_logic1[190] , \mprj_logic1[189] , \mprj_logic1[188] , \mprj_logic1[187] , \mprj_logic1[186] , \mprj_logic1[185] , \mprj_logic1[184] , \mprj_logic1[183] , \mprj_logic1[182] , \mprj_logic1[181] , \mprj_logic1[180] , \mprj_logic1[179] , \mprj_logic1[178] , \mprj_logic1[177] , \mprj_logic1[176] , \mprj_logic1[175] , \mprj_logic1[174] , \mprj_logic1[173] , \mprj_logic1[172] , \mprj_logic1[171] , \mprj_logic1[170] , \mprj_logic1[169] , \mprj_logic1[168] , \mprj_logic1[167] , \mprj_logic1[166] , \mprj_logic1[165] , \mprj_logic1[164] , \mprj_logic1[163] , \mprj_logic1[162] , \mprj_logic1[161] , \mprj_logic1[160] , \mprj_logic1[159] , \mprj_logic1[158] , \mprj_logic1[157] , \mprj_logic1[156] , \mprj_logic1[155] , \mprj_logic1[154] , \mprj_logic1[153] , \mprj_logic1[152] , \mprj_logic1[151] , \mprj_logic1[150] , \mprj_logic1[149] , \mprj_logic1[148] , \mprj_logic1[147] , \mprj_logic1[146] , \mprj_logic1[145] , \mprj_logic1[144] , \mprj_logic1[143] , \mprj_logic1[142] , \mprj_logic1[141] , \mprj_logic1[140] , \mprj_logic1[139] , \mprj_logic1[138] , \mprj_logic1[137] , \mprj_logic1[136] , \mprj_logic1[135] , \mprj_logic1[134] , \mprj_logic1[133] , \mprj_logic1[132] , \mprj_logic1[131] , \mprj_logic1[130] , \mprj_logic1[129] , \mprj_logic1[128] , \mprj_logic1[127] , \mprj_logic1[126] , \mprj_logic1[125] , \mprj_logic1[124] , \mprj_logic1[123] , \mprj_logic1[122] , \mprj_logic1[121] , \mprj_logic1[120] , \mprj_logic1[119] , \mprj_logic1[118] , \mprj_logic1[117] , \mprj_logic1[116] , \mprj_logic1[115] , \mprj_logic1[114] , \mprj_logic1[113] , \mprj_logic1[112] , \mprj_logic1[111] , \mprj_logic1[110] , \mprj_logic1[109] , \mprj_logic1[108] , \mprj_logic1[107] , \mprj_logic1[106] , \mprj_logic1[105] , \mprj_logic1[104] , \mprj_logic1[103] , \mprj_logic1[102] , \mprj_logic1[101] , \mprj_logic1[100] , \mprj_logic1[99] , \mprj_logic1[98] , \mprj_logic1[97] , \mprj_logic1[96] , \mprj_logic1[95] , \mprj_logic1[94] , \mprj_logic1[93] , \mprj_logic1[92] , \mprj_logic1[91] , \mprj_logic1[90] , \mprj_logic1[89] , \mprj_logic1[88] , \mprj_logic1[87] , \mprj_logic1[86] , \mprj_logic1[85] , \mprj_logic1[84] , \mprj_logic1[83] , \mprj_logic1[82] , \mprj_logic1[81] , \mprj_logic1[80] , \mprj_logic1[79] , \mprj_logic1[78] , \mprj_logic1[77] , \mprj_logic1[76] , \mprj_logic1[75] , \mprj_logic1[74] , \mprj_logic1[73] , \mprj_logic1[72] , \mprj_logic1[71] , \mprj_logic1[70] , \mprj_logic1[69] , \mprj_logic1[68] , \mprj_logic1[67] , \mprj_logic1[66] , \mprj_logic1[65] , \mprj_logic1[64] , \mprj_logic1[63] , \mprj_logic1[62] , \mprj_logic1[61] , \mprj_logic1[60] , \mprj_logic1[59] , \mprj_logic1[58] , \mprj_logic1[57] , \mprj_logic1[56] , \mprj_logic1[55] , \mprj_logic1[54] , \mprj_logic1[53] , \mprj_logic1[52] , \mprj_logic1[51] , \mprj_logic1[50] , \mprj_logic1[49] , \mprj_logic1[48] , \mprj_logic1[47] , \mprj_logic1[46] , \mprj_logic1[45] , \mprj_logic1[44] , \mprj_logic1[43] , \mprj_logic1[42] , \mprj_logic1[41] , \mprj_logic1[40] , \mprj_logic1[39] , \mprj_logic1[38] , \mprj_logic1[37] , \mprj_logic1[36] , \mprj_logic1[35] , \mprj_logic1[34] , \mprj_logic1[33] , \mprj_logic1[32] , \mprj_logic1[31] , \mprj_logic1[30] , \mprj_logic1[29] , \mprj_logic1[28] , \mprj_logic1[27] , \mprj_logic1[26] , \mprj_logic1[25] , \mprj_logic1[24] , \mprj_logic1[23] , \mprj_logic1[22] , \mprj_logic1[21] , \mprj_logic1[20] , \mprj_logic1[19] , \mprj_logic1[18] , \mprj_logic1[17] , \mprj_logic1[16] , \mprj_logic1[15] , \mprj_logic1[14] , \mprj_logic1[13] , \mprj_logic1[12] , \mprj_logic1[11] , \mprj_logic1[10] , \mprj_logic1[9] , \mprj_logic1[8] , \mprj_logic1[7] , \mprj_logic1[6] , \mprj_logic1[5] , \mprj_logic1[4] , \mprj_logic1[3] , \mprj_logic1[2] , \mprj_logic1[1] , \mprj_logic1[0]  }),
    .vccd1(vccd1),
    .vssd1(vssd1)
  );
  sky130_fd_sc_hd__buf_8 mprj_pwrgood (
    .A(\mprj_logic1[458] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .X(user1_vcc_powergood)
  );
  sky130_fd_sc_hd__einvp_8 mprj_rstn_buf (
    .A(_000_),
    .TE(\mprj_logic1[0] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(user_resetn)
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[0]  (
    .A(_006_),
    .TE(\mprj_logic1[6] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_sel_o_user[0])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[1]  (
    .A(_007_),
    .TE(\mprj_logic1[7] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_sel_o_user[1])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[2]  (
    .A(_008_),
    .TE(\mprj_logic1[8] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_sel_o_user[2])
  );
  sky130_fd_sc_hd__einvp_8 \mprj_sel_buf[3]  (
    .A(_009_),
    .TE(\mprj_logic1[9] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_sel_o_user[3])
  );
  sky130_fd_sc_hd__einvp_8 mprj_stb_buf (
    .A(_004_),
    .TE(\mprj_logic1[4] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_stb_o_user)
  );
  sky130_fd_sc_hd__buf_8 mprj_vdd_pwrgood (
    .A(mprj_vdd_logic1),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .X(user1_vdd_powergood)
  );
  sky130_fd_sc_hd__einvp_8 mprj_we_buf (
    .A(_005_),
    .TE(\mprj_logic1[5] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(mprj_we_o_user)
  );
  mgmt_protect_hv powergood_check (
    .mprj2_vdd_logic1(mprj2_vdd_logic1),
    .mprj_vdd_logic1(mprj_vdd_logic1),
    .vccd(vccd),
    .vdda1(vdda1),
    .vdda2(vdda2),
    .vssa1(vssa1),
    .vssa2(vssa2),
    .vssd(vssd)
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[0]  (
    .A(\la_data_in_mprj_bar[0] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[0])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[100]  (
    .A(\la_data_in_mprj_bar[100] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[100])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[101]  (
    .A(\la_data_in_mprj_bar[101] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[101])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[102]  (
    .A(\la_data_in_mprj_bar[102] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[102])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[103]  (
    .A(\la_data_in_mprj_bar[103] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[103])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[104]  (
    .A(\la_data_in_mprj_bar[104] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[104])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[105]  (
    .A(\la_data_in_mprj_bar[105] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[105])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[106]  (
    .A(\la_data_in_mprj_bar[106] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[106])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[107]  (
    .A(\la_data_in_mprj_bar[107] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[107])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[108]  (
    .A(\la_data_in_mprj_bar[108] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[108])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[109]  (
    .A(\la_data_in_mprj_bar[109] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[109])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[10]  (
    .A(\la_data_in_mprj_bar[10] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[10])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[110]  (
    .A(\la_data_in_mprj_bar[110] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[110])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[111]  (
    .A(\la_data_in_mprj_bar[111] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[111])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[112]  (
    .A(\la_data_in_mprj_bar[112] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[112])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[113]  (
    .A(\la_data_in_mprj_bar[113] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[113])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[114]  (
    .A(\la_data_in_mprj_bar[114] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[114])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[115]  (
    .A(\la_data_in_mprj_bar[115] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[115])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[116]  (
    .A(\la_data_in_mprj_bar[116] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[116])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[117]  (
    .A(\la_data_in_mprj_bar[117] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[117])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[118]  (
    .A(\la_data_in_mprj_bar[118] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[118])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[119]  (
    .A(\la_data_in_mprj_bar[119] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[119])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[11]  (
    .A(\la_data_in_mprj_bar[11] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[11])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[120]  (
    .A(\la_data_in_mprj_bar[120] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[120])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[121]  (
    .A(\la_data_in_mprj_bar[121] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[121])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[122]  (
    .A(\la_data_in_mprj_bar[122] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[122])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[123]  (
    .A(\la_data_in_mprj_bar[123] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[123])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[124]  (
    .A(\la_data_in_mprj_bar[124] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[124])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[125]  (
    .A(\la_data_in_mprj_bar[125] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[125])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[126]  (
    .A(\la_data_in_mprj_bar[126] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[126])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[127]  (
    .A(\la_data_in_mprj_bar[127] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[127])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[12]  (
    .A(\la_data_in_mprj_bar[12] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[12])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[13]  (
    .A(\la_data_in_mprj_bar[13] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[13])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[14]  (
    .A(\la_data_in_mprj_bar[14] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[14])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[15]  (
    .A(\la_data_in_mprj_bar[15] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[15])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[16]  (
    .A(\la_data_in_mprj_bar[16] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[16])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[17]  (
    .A(\la_data_in_mprj_bar[17] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[17])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[18]  (
    .A(\la_data_in_mprj_bar[18] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[18])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[19]  (
    .A(\la_data_in_mprj_bar[19] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[19])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[1]  (
    .A(\la_data_in_mprj_bar[1] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[1])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[20]  (
    .A(\la_data_in_mprj_bar[20] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[20])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[21]  (
    .A(\la_data_in_mprj_bar[21] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[21])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[22]  (
    .A(\la_data_in_mprj_bar[22] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[22])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[23]  (
    .A(\la_data_in_mprj_bar[23] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[23])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[24]  (
    .A(\la_data_in_mprj_bar[24] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[24])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[25]  (
    .A(\la_data_in_mprj_bar[25] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[25])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[26]  (
    .A(\la_data_in_mprj_bar[26] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[26])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[27]  (
    .A(\la_data_in_mprj_bar[27] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[27])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[28]  (
    .A(\la_data_in_mprj_bar[28] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[28])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[29]  (
    .A(\la_data_in_mprj_bar[29] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[29])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[2]  (
    .A(\la_data_in_mprj_bar[2] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[2])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[30]  (
    .A(\la_data_in_mprj_bar[30] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[30])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[31]  (
    .A(\la_data_in_mprj_bar[31] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[31])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[32]  (
    .A(\la_data_in_mprj_bar[32] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[32])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[33]  (
    .A(\la_data_in_mprj_bar[33] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[33])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[34]  (
    .A(\la_data_in_mprj_bar[34] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[34])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[35]  (
    .A(\la_data_in_mprj_bar[35] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[35])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[36]  (
    .A(\la_data_in_mprj_bar[36] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[36])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[37]  (
    .A(\la_data_in_mprj_bar[37] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[37])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[38]  (
    .A(\la_data_in_mprj_bar[38] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[38])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[39]  (
    .A(\la_data_in_mprj_bar[39] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[39])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[3]  (
    .A(\la_data_in_mprj_bar[3] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[3])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[40]  (
    .A(\la_data_in_mprj_bar[40] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[40])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[41]  (
    .A(\la_data_in_mprj_bar[41] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[41])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[42]  (
    .A(\la_data_in_mprj_bar[42] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[42])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[43]  (
    .A(\la_data_in_mprj_bar[43] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[43])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[44]  (
    .A(\la_data_in_mprj_bar[44] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[44])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[45]  (
    .A(\la_data_in_mprj_bar[45] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[45])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[46]  (
    .A(\la_data_in_mprj_bar[46] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[46])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[47]  (
    .A(\la_data_in_mprj_bar[47] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[47])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[48]  (
    .A(\la_data_in_mprj_bar[48] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[48])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[49]  (
    .A(\la_data_in_mprj_bar[49] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[49])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[4]  (
    .A(\la_data_in_mprj_bar[4] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[4])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[50]  (
    .A(\la_data_in_mprj_bar[50] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[50])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[51]  (
    .A(\la_data_in_mprj_bar[51] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[51])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[52]  (
    .A(\la_data_in_mprj_bar[52] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[52])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[53]  (
    .A(\la_data_in_mprj_bar[53] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[53])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[54]  (
    .A(\la_data_in_mprj_bar[54] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[54])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[55]  (
    .A(\la_data_in_mprj_bar[55] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[55])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[56]  (
    .A(\la_data_in_mprj_bar[56] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[56])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[57]  (
    .A(\la_data_in_mprj_bar[57] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[57])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[58]  (
    .A(\la_data_in_mprj_bar[58] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[58])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[59]  (
    .A(\la_data_in_mprj_bar[59] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[59])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[5]  (
    .A(\la_data_in_mprj_bar[5] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[5])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[60]  (
    .A(\la_data_in_mprj_bar[60] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[60])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[61]  (
    .A(\la_data_in_mprj_bar[61] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[61])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[62]  (
    .A(\la_data_in_mprj_bar[62] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[62])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[63]  (
    .A(\la_data_in_mprj_bar[63] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[63])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[64]  (
    .A(\la_data_in_mprj_bar[64] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[64])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[65]  (
    .A(\la_data_in_mprj_bar[65] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[65])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[66]  (
    .A(\la_data_in_mprj_bar[66] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[66])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[67]  (
    .A(\la_data_in_mprj_bar[67] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[67])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[68]  (
    .A(\la_data_in_mprj_bar[68] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[68])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[69]  (
    .A(\la_data_in_mprj_bar[69] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[69])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[6]  (
    .A(\la_data_in_mprj_bar[6] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[6])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[70]  (
    .A(\la_data_in_mprj_bar[70] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[70])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[71]  (
    .A(\la_data_in_mprj_bar[71] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[71])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[72]  (
    .A(\la_data_in_mprj_bar[72] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[72])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[73]  (
    .A(\la_data_in_mprj_bar[73] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[73])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[74]  (
    .A(\la_data_in_mprj_bar[74] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[74])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[75]  (
    .A(\la_data_in_mprj_bar[75] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[75])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[76]  (
    .A(\la_data_in_mprj_bar[76] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[76])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[77]  (
    .A(\la_data_in_mprj_bar[77] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[77])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[78]  (
    .A(\la_data_in_mprj_bar[78] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[78])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[79]  (
    .A(\la_data_in_mprj_bar[79] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[79])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[7]  (
    .A(\la_data_in_mprj_bar[7] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[7])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[80]  (
    .A(\la_data_in_mprj_bar[80] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[80])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[81]  (
    .A(\la_data_in_mprj_bar[81] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[81])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[82]  (
    .A(\la_data_in_mprj_bar[82] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[82])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[83]  (
    .A(\la_data_in_mprj_bar[83] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[83])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[84]  (
    .A(\la_data_in_mprj_bar[84] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[84])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[85]  (
    .A(\la_data_in_mprj_bar[85] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[85])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[86]  (
    .A(\la_data_in_mprj_bar[86] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[86])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[87]  (
    .A(\la_data_in_mprj_bar[87] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[87])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[88]  (
    .A(\la_data_in_mprj_bar[88] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[88])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[89]  (
    .A(\la_data_in_mprj_bar[89] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[89])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[8]  (
    .A(\la_data_in_mprj_bar[8] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[8])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[90]  (
    .A(\la_data_in_mprj_bar[90] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[90])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[91]  (
    .A(\la_data_in_mprj_bar[91] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[91])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[92]  (
    .A(\la_data_in_mprj_bar[92] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[92])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[93]  (
    .A(\la_data_in_mprj_bar[93] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[93])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[94]  (
    .A(\la_data_in_mprj_bar[94] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[94])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[95]  (
    .A(\la_data_in_mprj_bar[95] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[95])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[96]  (
    .A(\la_data_in_mprj_bar[96] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[96])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[97]  (
    .A(\la_data_in_mprj_bar[97] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[97])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[98]  (
    .A(\la_data_in_mprj_bar[98] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[98])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[99]  (
    .A(\la_data_in_mprj_bar[99] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[99])
  );
  sky130_fd_sc_hd__inv_8 \user_to_mprj_in_buffers[9]  (
    .A(\la_data_in_mprj_bar[9] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(la_data_in_mprj[9])
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[0]  (
    .A(la_data_out_core[0]),
    .B(\mprj_logic1[330] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[0] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[100]  (
    .A(la_data_out_core[100]),
    .B(\mprj_logic1[430] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[100] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[101]  (
    .A(la_data_out_core[101]),
    .B(\mprj_logic1[431] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[101] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[102]  (
    .A(la_data_out_core[102]),
    .B(\mprj_logic1[432] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[102] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[103]  (
    .A(la_data_out_core[103]),
    .B(\mprj_logic1[433] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[103] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[104]  (
    .A(la_data_out_core[104]),
    .B(\mprj_logic1[434] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[104] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[105]  (
    .A(la_data_out_core[105]),
    .B(\mprj_logic1[435] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[105] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[106]  (
    .A(la_data_out_core[106]),
    .B(\mprj_logic1[436] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[106] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[107]  (
    .A(la_data_out_core[107]),
    .B(\mprj_logic1[437] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[107] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[108]  (
    .A(la_data_out_core[108]),
    .B(\mprj_logic1[438] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[108] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[109]  (
    .A(la_data_out_core[109]),
    .B(\mprj_logic1[439] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[109] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[10]  (
    .A(la_data_out_core[10]),
    .B(\mprj_logic1[340] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[10] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[110]  (
    .A(la_data_out_core[110]),
    .B(\mprj_logic1[440] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[110] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[111]  (
    .A(la_data_out_core[111]),
    .B(\mprj_logic1[441] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[111] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[112]  (
    .A(la_data_out_core[112]),
    .B(\mprj_logic1[442] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[112] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[113]  (
    .A(la_data_out_core[113]),
    .B(\mprj_logic1[443] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[113] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[114]  (
    .A(la_data_out_core[114]),
    .B(\mprj_logic1[444] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[114] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[115]  (
    .A(la_data_out_core[115]),
    .B(\mprj_logic1[445] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[115] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[116]  (
    .A(la_data_out_core[116]),
    .B(\mprj_logic1[446] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[116] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[117]  (
    .A(la_data_out_core[117]),
    .B(\mprj_logic1[447] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[117] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[118]  (
    .A(la_data_out_core[118]),
    .B(\mprj_logic1[448] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[118] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[119]  (
    .A(la_data_out_core[119]),
    .B(\mprj_logic1[449] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[119] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[11]  (
    .A(la_data_out_core[11]),
    .B(\mprj_logic1[341] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[11] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[120]  (
    .A(la_data_out_core[120]),
    .B(\mprj_logic1[450] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[120] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[121]  (
    .A(la_data_out_core[121]),
    .B(\mprj_logic1[451] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[121] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[122]  (
    .A(la_data_out_core[122]),
    .B(\mprj_logic1[452] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[122] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[123]  (
    .A(la_data_out_core[123]),
    .B(\mprj_logic1[453] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[123] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[124]  (
    .A(la_data_out_core[124]),
    .B(\mprj_logic1[454] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[124] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[125]  (
    .A(la_data_out_core[125]),
    .B(\mprj_logic1[455] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[125] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[126]  (
    .A(la_data_out_core[126]),
    .B(\mprj_logic1[456] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[126] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[127]  (
    .A(la_data_out_core[127]),
    .B(\mprj_logic1[457] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[127] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[12]  (
    .A(la_data_out_core[12]),
    .B(\mprj_logic1[342] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[12] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[13]  (
    .A(la_data_out_core[13]),
    .B(\mprj_logic1[343] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[13] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[14]  (
    .A(la_data_out_core[14]),
    .B(\mprj_logic1[344] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[14] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[15]  (
    .A(la_data_out_core[15]),
    .B(\mprj_logic1[345] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[15] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[16]  (
    .A(la_data_out_core[16]),
    .B(\mprj_logic1[346] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[16] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[17]  (
    .A(la_data_out_core[17]),
    .B(\mprj_logic1[347] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[17] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[18]  (
    .A(la_data_out_core[18]),
    .B(\mprj_logic1[348] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[18] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[19]  (
    .A(la_data_out_core[19]),
    .B(\mprj_logic1[349] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[19] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[1]  (
    .A(la_data_out_core[1]),
    .B(\mprj_logic1[331] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[1] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[20]  (
    .A(la_data_out_core[20]),
    .B(\mprj_logic1[350] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[20] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[21]  (
    .A(la_data_out_core[21]),
    .B(\mprj_logic1[351] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[21] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[22]  (
    .A(la_data_out_core[22]),
    .B(\mprj_logic1[352] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[22] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[23]  (
    .A(la_data_out_core[23]),
    .B(\mprj_logic1[353] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[23] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[24]  (
    .A(la_data_out_core[24]),
    .B(\mprj_logic1[354] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[24] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[25]  (
    .A(la_data_out_core[25]),
    .B(\mprj_logic1[355] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[25] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[26]  (
    .A(la_data_out_core[26]),
    .B(\mprj_logic1[356] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[26] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[27]  (
    .A(la_data_out_core[27]),
    .B(\mprj_logic1[357] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[27] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[28]  (
    .A(la_data_out_core[28]),
    .B(\mprj_logic1[358] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[28] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[29]  (
    .A(la_data_out_core[29]),
    .B(\mprj_logic1[359] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[29] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[2]  (
    .A(la_data_out_core[2]),
    .B(\mprj_logic1[332] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[2] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[30]  (
    .A(la_data_out_core[30]),
    .B(\mprj_logic1[360] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[30] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[31]  (
    .A(la_data_out_core[31]),
    .B(\mprj_logic1[361] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[31] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[32]  (
    .A(la_data_out_core[32]),
    .B(\mprj_logic1[362] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[32] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[33]  (
    .A(la_data_out_core[33]),
    .B(\mprj_logic1[363] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[33] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[34]  (
    .A(la_data_out_core[34]),
    .B(\mprj_logic1[364] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[34] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[35]  (
    .A(la_data_out_core[35]),
    .B(\mprj_logic1[365] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[35] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[36]  (
    .A(la_data_out_core[36]),
    .B(\mprj_logic1[366] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[36] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[37]  (
    .A(la_data_out_core[37]),
    .B(\mprj_logic1[367] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[37] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[38]  (
    .A(la_data_out_core[38]),
    .B(\mprj_logic1[368] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[38] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[39]  (
    .A(la_data_out_core[39]),
    .B(\mprj_logic1[369] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[39] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[3]  (
    .A(la_data_out_core[3]),
    .B(\mprj_logic1[333] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[3] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[40]  (
    .A(la_data_out_core[40]),
    .B(\mprj_logic1[370] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[40] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[41]  (
    .A(la_data_out_core[41]),
    .B(\mprj_logic1[371] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[41] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[42]  (
    .A(la_data_out_core[42]),
    .B(\mprj_logic1[372] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[42] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[43]  (
    .A(la_data_out_core[43]),
    .B(\mprj_logic1[373] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[43] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[44]  (
    .A(la_data_out_core[44]),
    .B(\mprj_logic1[374] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[44] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[45]  (
    .A(la_data_out_core[45]),
    .B(\mprj_logic1[375] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[45] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[46]  (
    .A(la_data_out_core[46]),
    .B(\mprj_logic1[376] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[46] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[47]  (
    .A(la_data_out_core[47]),
    .B(\mprj_logic1[377] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[47] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[48]  (
    .A(la_data_out_core[48]),
    .B(\mprj_logic1[378] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[48] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[49]  (
    .A(la_data_out_core[49]),
    .B(\mprj_logic1[379] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[49] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[4]  (
    .A(la_data_out_core[4]),
    .B(\mprj_logic1[334] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[4] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[50]  (
    .A(la_data_out_core[50]),
    .B(\mprj_logic1[380] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[50] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[51]  (
    .A(la_data_out_core[51]),
    .B(\mprj_logic1[381] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[51] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[52]  (
    .A(la_data_out_core[52]),
    .B(\mprj_logic1[382] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[52] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[53]  (
    .A(la_data_out_core[53]),
    .B(\mprj_logic1[383] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[53] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[54]  (
    .A(la_data_out_core[54]),
    .B(\mprj_logic1[384] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[54] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[55]  (
    .A(la_data_out_core[55]),
    .B(\mprj_logic1[385] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[55] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[56]  (
    .A(la_data_out_core[56]),
    .B(\mprj_logic1[386] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[56] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[57]  (
    .A(la_data_out_core[57]),
    .B(\mprj_logic1[387] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[57] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[58]  (
    .A(la_data_out_core[58]),
    .B(\mprj_logic1[388] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[58] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[59]  (
    .A(la_data_out_core[59]),
    .B(\mprj_logic1[389] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[59] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[5]  (
    .A(la_data_out_core[5]),
    .B(\mprj_logic1[335] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[5] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[60]  (
    .A(la_data_out_core[60]),
    .B(\mprj_logic1[390] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[60] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[61]  (
    .A(la_data_out_core[61]),
    .B(\mprj_logic1[391] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[61] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[62]  (
    .A(la_data_out_core[62]),
    .B(\mprj_logic1[392] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[62] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[63]  (
    .A(la_data_out_core[63]),
    .B(\mprj_logic1[393] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[63] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[64]  (
    .A(la_data_out_core[64]),
    .B(\mprj_logic1[394] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[64] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[65]  (
    .A(la_data_out_core[65]),
    .B(\mprj_logic1[395] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[65] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[66]  (
    .A(la_data_out_core[66]),
    .B(\mprj_logic1[396] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[66] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[67]  (
    .A(la_data_out_core[67]),
    .B(\mprj_logic1[397] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[67] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[68]  (
    .A(la_data_out_core[68]),
    .B(\mprj_logic1[398] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[68] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[69]  (
    .A(la_data_out_core[69]),
    .B(\mprj_logic1[399] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[69] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[6]  (
    .A(la_data_out_core[6]),
    .B(\mprj_logic1[336] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[6] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[70]  (
    .A(la_data_out_core[70]),
    .B(\mprj_logic1[400] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[70] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[71]  (
    .A(la_data_out_core[71]),
    .B(\mprj_logic1[401] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[71] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[72]  (
    .A(la_data_out_core[72]),
    .B(\mprj_logic1[402] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[72] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[73]  (
    .A(la_data_out_core[73]),
    .B(\mprj_logic1[403] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[73] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[74]  (
    .A(la_data_out_core[74]),
    .B(\mprj_logic1[404] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[74] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[75]  (
    .A(la_data_out_core[75]),
    .B(\mprj_logic1[405] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[75] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[76]  (
    .A(la_data_out_core[76]),
    .B(\mprj_logic1[406] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[76] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[77]  (
    .A(la_data_out_core[77]),
    .B(\mprj_logic1[407] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[77] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[78]  (
    .A(la_data_out_core[78]),
    .B(\mprj_logic1[408] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[78] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[79]  (
    .A(la_data_out_core[79]),
    .B(\mprj_logic1[409] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[79] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[7]  (
    .A(la_data_out_core[7]),
    .B(\mprj_logic1[337] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[7] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[80]  (
    .A(la_data_out_core[80]),
    .B(\mprj_logic1[410] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[80] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[81]  (
    .A(la_data_out_core[81]),
    .B(\mprj_logic1[411] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[81] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[82]  (
    .A(la_data_out_core[82]),
    .B(\mprj_logic1[412] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[82] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[83]  (
    .A(la_data_out_core[83]),
    .B(\mprj_logic1[413] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[83] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[84]  (
    .A(la_data_out_core[84]),
    .B(\mprj_logic1[414] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[84] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[85]  (
    .A(la_data_out_core[85]),
    .B(\mprj_logic1[415] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[85] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[86]  (
    .A(la_data_out_core[86]),
    .B(\mprj_logic1[416] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[86] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[87]  (
    .A(la_data_out_core[87]),
    .B(\mprj_logic1[417] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[87] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[88]  (
    .A(la_data_out_core[88]),
    .B(\mprj_logic1[418] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[88] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[89]  (
    .A(la_data_out_core[89]),
    .B(\mprj_logic1[419] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[89] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[8]  (
    .A(la_data_out_core[8]),
    .B(\mprj_logic1[338] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[8] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[90]  (
    .A(la_data_out_core[90]),
    .B(\mprj_logic1[420] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[90] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[91]  (
    .A(la_data_out_core[91]),
    .B(\mprj_logic1[421] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[91] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[92]  (
    .A(la_data_out_core[92]),
    .B(\mprj_logic1[422] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[92] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[93]  (
    .A(la_data_out_core[93]),
    .B(\mprj_logic1[423] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[93] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[94]  (
    .A(la_data_out_core[94]),
    .B(\mprj_logic1[424] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[94] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[95]  (
    .A(la_data_out_core[95]),
    .B(\mprj_logic1[425] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[95] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[96]  (
    .A(la_data_out_core[96]),
    .B(\mprj_logic1[426] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[96] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[97]  (
    .A(la_data_out_core[97]),
    .B(\mprj_logic1[427] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[97] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[98]  (
    .A(la_data_out_core[98]),
    .B(\mprj_logic1[428] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[98] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[99]  (
    .A(la_data_out_core[99]),
    .B(\mprj_logic1[429] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[99] )
  );
  sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[9]  (
    .A(la_data_out_core[9]),
    .B(\mprj_logic1[339] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Y(\la_data_in_mprj_bar[9] )
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[0]  (
    .A(_202_),
    .TE(\mprj_logic1[202] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[0])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[100]  (
    .A(_203_),
    .TE(\mprj_logic1[302] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[100])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[101]  (
    .A(_204_),
    .TE(\mprj_logic1[303] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[101])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[102]  (
    .A(_205_),
    .TE(\mprj_logic1[304] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[102])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[103]  (
    .A(_206_),
    .TE(\mprj_logic1[305] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[103])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[104]  (
    .A(_207_),
    .TE(\mprj_logic1[306] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[104])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[105]  (
    .A(_208_),
    .TE(\mprj_logic1[307] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[105])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[106]  (
    .A(_209_),
    .TE(\mprj_logic1[308] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[106])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[107]  (
    .A(_210_),
    .TE(\mprj_logic1[309] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[107])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[108]  (
    .A(_211_),
    .TE(\mprj_logic1[310] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[108])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[109]  (
    .A(_212_),
    .TE(\mprj_logic1[311] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[109])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[10]  (
    .A(_213_),
    .TE(\mprj_logic1[212] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[10])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[110]  (
    .A(_214_),
    .TE(\mprj_logic1[312] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[110])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[111]  (
    .A(_215_),
    .TE(\mprj_logic1[313] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[111])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[112]  (
    .A(_216_),
    .TE(\mprj_logic1[314] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[112])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[113]  (
    .A(_217_),
    .TE(\mprj_logic1[315] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[113])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[114]  (
    .A(_218_),
    .TE(\mprj_logic1[316] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[114])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[115]  (
    .A(_219_),
    .TE(\mprj_logic1[317] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[115])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[116]  (
    .A(_220_),
    .TE(\mprj_logic1[318] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[116])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[117]  (
    .A(_221_),
    .TE(\mprj_logic1[319] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[117])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[118]  (
    .A(_222_),
    .TE(\mprj_logic1[320] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[118])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[119]  (
    .A(_223_),
    .TE(\mprj_logic1[321] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[119])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[11]  (
    .A(_224_),
    .TE(\mprj_logic1[213] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[11])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[120]  (
    .A(_225_),
    .TE(\mprj_logic1[322] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[120])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[121]  (
    .A(_226_),
    .TE(\mprj_logic1[323] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[121])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[122]  (
    .A(_227_),
    .TE(\mprj_logic1[324] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[122])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[123]  (
    .A(_228_),
    .TE(\mprj_logic1[325] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[123])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[124]  (
    .A(_229_),
    .TE(\mprj_logic1[326] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[124])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[125]  (
    .A(_230_),
    .TE(\mprj_logic1[327] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[125])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[126]  (
    .A(_231_),
    .TE(\mprj_logic1[328] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[126])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[127]  (
    .A(_232_),
    .TE(\mprj_logic1[329] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[127])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[12]  (
    .A(_233_),
    .TE(\mprj_logic1[214] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[12])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[13]  (
    .A(_234_),
    .TE(\mprj_logic1[215] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[13])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[14]  (
    .A(_235_),
    .TE(\mprj_logic1[216] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[14])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[15]  (
    .A(_236_),
    .TE(\mprj_logic1[217] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[15])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[16]  (
    .A(_237_),
    .TE(\mprj_logic1[218] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[16])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[17]  (
    .A(_238_),
    .TE(\mprj_logic1[219] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[17])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[18]  (
    .A(_239_),
    .TE(\mprj_logic1[220] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[18])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[19]  (
    .A(_240_),
    .TE(\mprj_logic1[221] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[19])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[1]  (
    .A(_241_),
    .TE(\mprj_logic1[203] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[1])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[20]  (
    .A(_242_),
    .TE(\mprj_logic1[222] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[20])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[21]  (
    .A(_243_),
    .TE(\mprj_logic1[223] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[21])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[22]  (
    .A(_244_),
    .TE(\mprj_logic1[224] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[22])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[23]  (
    .A(_245_),
    .TE(\mprj_logic1[225] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[23])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[24]  (
    .A(_246_),
    .TE(\mprj_logic1[226] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[24])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[25]  (
    .A(_247_),
    .TE(\mprj_logic1[227] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[25])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[26]  (
    .A(_248_),
    .TE(\mprj_logic1[228] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[26])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[27]  (
    .A(_249_),
    .TE(\mprj_logic1[229] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[27])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[28]  (
    .A(_250_),
    .TE(\mprj_logic1[230] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[28])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[29]  (
    .A(_251_),
    .TE(\mprj_logic1[231] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[29])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[2]  (
    .A(_252_),
    .TE(\mprj_logic1[204] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[2])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[30]  (
    .A(_253_),
    .TE(\mprj_logic1[232] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[30])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[31]  (
    .A(_254_),
    .TE(\mprj_logic1[233] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[31])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[32]  (
    .A(_255_),
    .TE(\mprj_logic1[234] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[32])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[33]  (
    .A(_256_),
    .TE(\mprj_logic1[235] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[33])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[34]  (
    .A(_257_),
    .TE(\mprj_logic1[236] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[34])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[35]  (
    .A(_258_),
    .TE(\mprj_logic1[237] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[35])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[36]  (
    .A(_259_),
    .TE(\mprj_logic1[238] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[36])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[37]  (
    .A(_260_),
    .TE(\mprj_logic1[239] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[37])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[38]  (
    .A(_261_),
    .TE(\mprj_logic1[240] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[38])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[39]  (
    .A(_262_),
    .TE(\mprj_logic1[241] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[39])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[3]  (
    .A(_263_),
    .TE(\mprj_logic1[205] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[3])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[40]  (
    .A(_264_),
    .TE(\mprj_logic1[242] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[40])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[41]  (
    .A(_265_),
    .TE(\mprj_logic1[243] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[41])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[42]  (
    .A(_266_),
    .TE(\mprj_logic1[244] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[42])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[43]  (
    .A(_267_),
    .TE(\mprj_logic1[245] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[43])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[44]  (
    .A(_268_),
    .TE(\mprj_logic1[246] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[44])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[45]  (
    .A(_269_),
    .TE(\mprj_logic1[247] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[45])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[46]  (
    .A(_270_),
    .TE(\mprj_logic1[248] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[46])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[47]  (
    .A(_271_),
    .TE(\mprj_logic1[249] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[47])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[48]  (
    .A(_272_),
    .TE(\mprj_logic1[250] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[48])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[49]  (
    .A(_273_),
    .TE(\mprj_logic1[251] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[49])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[4]  (
    .A(_274_),
    .TE(\mprj_logic1[206] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[4])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[50]  (
    .A(_275_),
    .TE(\mprj_logic1[252] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[50])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[51]  (
    .A(_276_),
    .TE(\mprj_logic1[253] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[51])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[52]  (
    .A(_277_),
    .TE(\mprj_logic1[254] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[52])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[53]  (
    .A(_278_),
    .TE(\mprj_logic1[255] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[53])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[54]  (
    .A(_279_),
    .TE(\mprj_logic1[256] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[54])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[55]  (
    .A(_280_),
    .TE(\mprj_logic1[257] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[55])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[56]  (
    .A(_281_),
    .TE(\mprj_logic1[258] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[56])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[57]  (
    .A(_282_),
    .TE(\mprj_logic1[259] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[57])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[58]  (
    .A(_283_),
    .TE(\mprj_logic1[260] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[58])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[59]  (
    .A(_284_),
    .TE(\mprj_logic1[261] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[59])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[5]  (
    .A(_285_),
    .TE(\mprj_logic1[207] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[5])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[60]  (
    .A(_286_),
    .TE(\mprj_logic1[262] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[60])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[61]  (
    .A(_287_),
    .TE(\mprj_logic1[263] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[61])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[62]  (
    .A(_288_),
    .TE(\mprj_logic1[264] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[62])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[63]  (
    .A(_289_),
    .TE(\mprj_logic1[265] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[63])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[64]  (
    .A(_290_),
    .TE(\mprj_logic1[266] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[64])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[65]  (
    .A(_291_),
    .TE(\mprj_logic1[267] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[65])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[66]  (
    .A(_292_),
    .TE(\mprj_logic1[268] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[66])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[67]  (
    .A(_293_),
    .TE(\mprj_logic1[269] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[67])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[68]  (
    .A(_294_),
    .TE(\mprj_logic1[270] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[68])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[69]  (
    .A(_295_),
    .TE(\mprj_logic1[271] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[69])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[6]  (
    .A(_296_),
    .TE(\mprj_logic1[208] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[6])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[70]  (
    .A(_297_),
    .TE(\mprj_logic1[272] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[70])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[71]  (
    .A(_298_),
    .TE(\mprj_logic1[273] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[71])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[72]  (
    .A(_299_),
    .TE(\mprj_logic1[274] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[72])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[73]  (
    .A(_300_),
    .TE(\mprj_logic1[275] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[73])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[74]  (
    .A(_301_),
    .TE(\mprj_logic1[276] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[74])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[75]  (
    .A(_302_),
    .TE(\mprj_logic1[277] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[75])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[76]  (
    .A(_303_),
    .TE(\mprj_logic1[278] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[76])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[77]  (
    .A(_304_),
    .TE(\mprj_logic1[279] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[77])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[78]  (
    .A(_305_),
    .TE(\mprj_logic1[280] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[78])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[79]  (
    .A(_306_),
    .TE(\mprj_logic1[281] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[79])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[7]  (
    .A(_307_),
    .TE(\mprj_logic1[209] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[7])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[80]  (
    .A(_308_),
    .TE(\mprj_logic1[282] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[80])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[81]  (
    .A(_309_),
    .TE(\mprj_logic1[283] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[81])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[82]  (
    .A(_310_),
    .TE(\mprj_logic1[284] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[82])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[83]  (
    .A(_311_),
    .TE(\mprj_logic1[285] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[83])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[84]  (
    .A(_312_),
    .TE(\mprj_logic1[286] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[84])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[85]  (
    .A(_313_),
    .TE(\mprj_logic1[287] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[85])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[86]  (
    .A(_314_),
    .TE(\mprj_logic1[288] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[86])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[87]  (
    .A(_315_),
    .TE(\mprj_logic1[289] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[87])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[88]  (
    .A(_316_),
    .TE(\mprj_logic1[290] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[88])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[89]  (
    .A(_317_),
    .TE(\mprj_logic1[291] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[89])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[8]  (
    .A(_318_),
    .TE(\mprj_logic1[210] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[8])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[90]  (
    .A(_319_),
    .TE(\mprj_logic1[292] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[90])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[91]  (
    .A(_320_),
    .TE(\mprj_logic1[293] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[91])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[92]  (
    .A(_321_),
    .TE(\mprj_logic1[294] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[92])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[93]  (
    .A(_322_),
    .TE(\mprj_logic1[295] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[93])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[94]  (
    .A(_323_),
    .TE(\mprj_logic1[296] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[94])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[95]  (
    .A(_324_),
    .TE(\mprj_logic1[297] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[95])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[96]  (
    .A(_325_),
    .TE(\mprj_logic1[298] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[96])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[97]  (
    .A(_326_),
    .TE(\mprj_logic1[299] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[97])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[98]  (
    .A(_327_),
    .TE(\mprj_logic1[300] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[98])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[99]  (
    .A(_328_),
    .TE(\mprj_logic1[301] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[99])
  );
  sky130_fd_sc_hd__einvp_8 \user_to_mprj_oen_buffers[9]  (
    .A(_329_),
    .TE(\mprj_logic1[211] ),
    .VGND(vssd),
    .VNB(vssd),
    .VPB(vccd),
    .VPWR(vccd),
    .Z(la_oen_core[9])
  );
endmodule
