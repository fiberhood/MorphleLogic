magic
tech sky130A
magscale 1 2
timestamp 1608074286
<< nwell >>
rect 1066 296741 1340 297307
rect 298660 296741 298854 297307
rect 1066 295653 1340 296219
rect 298660 295653 298854 296219
rect 1066 294565 1340 295131
rect 298660 294565 298854 295131
rect 1066 293477 1340 294043
rect 298660 293477 298854 294043
rect 1066 292389 1340 292955
rect 298660 292389 298854 292955
rect 1066 291301 1340 291867
rect 298660 291301 298854 291867
rect 1066 290213 1340 290779
rect 298660 290213 298854 290779
rect 1066 289125 1340 289691
rect 298660 289125 298854 289691
rect 1066 288037 1340 288603
rect 298660 288037 298854 288603
rect 1066 286949 1340 287515
rect 298660 286949 298854 287515
rect 1066 285861 1340 286427
rect 298660 285861 298854 286427
rect 1066 284773 1340 285339
rect 298660 284773 298854 285339
rect 1066 283685 1340 284251
rect 298660 283685 298854 284251
rect 1066 282597 1340 283163
rect 298660 282597 298854 283163
rect 1066 281509 1340 282075
rect 298660 281509 298854 282075
rect 1066 280421 1340 280987
rect 298660 280421 298854 280987
rect 1066 279333 1340 279899
rect 298660 279333 298854 279899
rect 1066 278245 1340 278811
rect 298660 278245 298854 278811
rect 1066 277157 1340 277723
rect 298660 277157 298854 277723
rect 1066 276069 1340 276635
rect 298660 276069 298854 276635
rect 1066 274981 1340 275547
rect 298660 274981 298854 275547
rect 1066 273893 1340 274459
rect 298660 273893 298854 274459
rect 1066 272805 1340 273371
rect 298660 272805 298854 273371
rect 1066 271717 1340 272283
rect 298660 271717 298854 272283
rect 1066 270629 1340 271195
rect 298660 270629 298854 271195
rect 1066 269541 1340 270107
rect 298660 269541 298854 270107
rect 1066 268453 1340 269019
rect 298660 268453 298854 269019
rect 1066 267365 1340 267931
rect 298660 267365 298854 267931
rect 1066 266277 1340 266843
rect 298660 266277 298854 266843
rect 1066 265189 1340 265755
rect 298660 265189 298854 265755
rect 1066 264101 1340 264667
rect 298660 264101 298854 264667
rect 1066 263013 1340 263579
rect 298660 263013 298854 263579
rect 1066 261925 1340 262491
rect 298660 261925 298854 262491
rect 1066 260837 1340 261403
rect 298660 260837 298854 261403
rect 1066 259749 1340 260315
rect 298660 259749 298854 260315
rect 1066 258661 1340 259227
rect 298660 258661 298854 259227
rect 1066 257573 1340 258139
rect 298660 257573 298854 258139
rect 1066 256485 1340 257051
rect 298660 256485 298854 257051
rect 1066 255397 1340 255963
rect 298660 255397 298854 255963
rect 1066 254309 1340 254875
rect 298660 254309 298854 254875
rect 1066 253221 1340 253787
rect 298660 253221 298854 253787
rect 1066 252133 1340 252699
rect 298660 252133 298854 252699
rect 1066 251045 1340 251611
rect 298660 251045 298854 251611
rect 1066 249957 1340 250523
rect 298660 249957 298854 250523
rect 1066 248869 1340 249435
rect 298660 248869 298854 249435
rect 1066 247781 1340 248347
rect 298660 247781 298854 248347
rect 1066 246693 1340 247259
rect 298660 246693 298854 247259
rect 1066 245605 1340 246171
rect 298660 245605 298854 246171
rect 1066 244517 1340 245083
rect 298660 244517 298854 245083
rect 1066 243429 1340 243995
rect 298660 243429 298854 243995
rect 1066 242341 1340 242907
rect 298660 242341 298854 242907
rect 1066 241253 1340 241819
rect 298660 241253 298854 241819
rect 1066 240165 1340 240731
rect 298660 240165 298854 240731
rect 1066 239077 1340 239643
rect 298660 239077 298854 239643
rect 1066 237989 1340 238555
rect 298660 237989 298854 238555
rect 1066 236901 1340 237467
rect 298660 236901 298854 237467
rect 1066 235813 1340 236379
rect 298660 235813 298854 236379
rect 1066 234725 1340 235291
rect 298660 234725 298854 235291
rect 1066 233637 1340 234203
rect 298660 233637 298854 234203
rect 1066 232549 1340 233115
rect 298660 232549 298854 233115
rect 1066 231461 1340 232027
rect 298660 231461 298854 232027
rect 1066 230373 1340 230939
rect 298660 230373 298854 230939
rect 1066 229285 1340 229851
rect 298660 229285 298854 229851
rect 1066 228197 1340 228763
rect 298660 228197 298854 228763
rect 1066 227109 1340 227675
rect 298660 227109 298854 227675
rect 1066 226021 1340 226587
rect 298660 226021 298854 226587
rect 1066 224933 1340 225499
rect 298660 224933 298854 225499
rect 1066 223845 1340 224411
rect 298660 223845 298854 224411
rect 1066 222757 1340 223323
rect 298660 222757 298854 223323
rect 1066 221669 1340 222235
rect 298660 221669 298854 222235
rect 1066 220581 1340 221147
rect 298660 220581 298854 221147
rect 1066 219493 1340 220059
rect 298660 219493 298854 220059
rect 1066 218405 1340 218971
rect 298660 218405 298854 218971
rect 1066 217317 1340 217883
rect 298660 217317 298854 217883
rect 1066 216229 1340 216795
rect 298660 216229 298854 216795
rect 1066 215141 1340 215707
rect 298660 215141 298854 215707
rect 1066 214053 1340 214619
rect 298660 214053 298854 214619
rect 1066 212965 1340 213531
rect 298660 212965 298854 213531
rect 1066 211877 1340 212443
rect 298660 211877 298854 212443
rect 1066 210789 1340 211355
rect 298660 210789 298854 211355
rect 1066 209701 1340 210267
rect 298660 209701 298854 210267
rect 1066 208613 1340 209179
rect 298660 208613 298854 209179
rect 1066 207525 1340 208091
rect 298660 207525 298854 208091
rect 1066 206437 1340 207003
rect 298660 206437 298854 207003
rect 1066 205349 1340 205915
rect 298660 205349 298854 205915
rect 1066 204261 1340 204827
rect 298660 204261 298854 204827
rect 1066 203173 1340 203739
rect 298660 203173 298854 203739
rect 1066 202085 1340 202651
rect 298660 202085 298854 202651
rect 1066 200997 1340 201563
rect 298660 200997 298854 201563
rect 1066 199909 1340 200475
rect 298660 199909 298854 200475
rect 1066 198821 1340 199387
rect 298660 198821 298854 199387
rect 1066 197733 1340 198299
rect 298660 197733 298854 198299
rect 1066 196645 1340 197211
rect 298660 196645 298854 197211
rect 1066 195557 1340 196123
rect 298660 195557 298854 196123
rect 1066 194469 1340 195035
rect 298660 194469 298854 195035
rect 1066 193381 1340 193947
rect 298660 193381 298854 193947
rect 1066 192293 1340 192859
rect 298660 192293 298854 192859
rect 1066 191205 1340 191771
rect 298660 191205 298854 191771
rect 1066 190117 1340 190683
rect 298660 190117 298854 190683
rect 1066 189029 1340 189595
rect 298660 189029 298854 189595
rect 1066 187941 1340 188507
rect 298660 187941 298854 188507
rect 1066 186853 1340 187419
rect 298660 186853 298854 187419
rect 1066 185765 1340 186331
rect 298660 185765 298854 186331
rect 1066 184677 1340 185243
rect 298660 184677 298854 185243
rect 1066 183589 1340 184155
rect 298660 183589 298854 184155
rect 1066 182501 1340 183067
rect 298660 182501 298854 183067
rect 1066 181413 1340 181979
rect 298660 181413 298854 181979
rect 1066 180325 1340 180891
rect 298660 180325 298854 180891
rect 1066 179237 1340 179803
rect 298660 179237 298854 179803
rect 1066 178149 1340 178715
rect 298660 178149 298854 178715
rect 1066 177061 1340 177627
rect 298660 177061 298854 177627
rect 1066 175973 1340 176539
rect 298660 175973 298854 176539
rect 1066 174885 1340 175451
rect 298660 174885 298854 175451
rect 1066 173797 1340 174363
rect 298660 173797 298854 174363
rect 1066 172709 1340 173275
rect 298660 172709 298854 173275
rect 1066 171621 1340 172187
rect 298660 171621 298854 172187
rect 1066 170533 1340 171099
rect 298660 170533 298854 171099
rect 1066 169445 1340 170011
rect 298660 169445 298854 170011
rect 1066 168357 1340 168923
rect 298660 168357 298854 168923
rect 1066 167269 1340 167835
rect 298660 167269 298854 167835
rect 1066 166181 1340 166747
rect 298660 166181 298854 166747
rect 1066 165093 1340 165659
rect 298660 165093 298854 165659
rect 1066 164005 1340 164571
rect 298660 164005 298854 164571
rect 1066 162917 1340 163483
rect 298660 162917 298854 163483
rect 1066 161829 1340 162395
rect 298660 161829 298854 162395
rect 1066 160741 1340 161307
rect 298660 160741 298854 161307
rect 1066 159653 1340 160219
rect 298660 159653 298854 160219
rect 1066 158565 1340 159131
rect 298660 158565 298854 159131
rect 1066 157477 1340 158043
rect 298660 157477 298854 158043
rect 1066 156389 1340 156955
rect 298660 156389 298854 156955
rect 1066 155301 1340 155867
rect 298660 155301 298854 155867
rect 1066 154213 1340 154779
rect 298660 154213 298854 154779
rect 1066 153125 1340 153691
rect 298660 153125 298854 153691
rect 1066 152037 1340 152603
rect 298660 152037 298854 152603
rect 1066 150949 1340 151515
rect 298660 150949 298854 151515
rect 1066 149861 1340 150427
rect 298660 149861 298854 150427
rect 1066 148773 1340 149339
rect 298660 148773 298854 149339
rect 1066 147685 1340 148251
rect 298660 147685 298854 148251
rect 1066 146597 1340 147163
rect 298660 146597 298854 147163
rect 1066 145509 1340 146075
rect 298660 145509 298854 146075
rect 1066 144421 1340 144987
rect 298660 144421 298854 144987
rect 1066 143333 1340 143899
rect 298660 143333 298854 143899
rect 1066 142245 1340 142811
rect 298660 142245 298854 142811
rect 1066 141157 1340 141723
rect 298660 141157 298854 141723
rect 1066 140069 1340 140635
rect 298660 140069 298854 140635
rect 1066 138981 1340 139547
rect 298660 138981 298854 139547
rect 1066 137893 1340 138459
rect 298660 137893 298854 138459
rect 1066 136805 1340 137371
rect 298660 136805 298854 137371
rect 1066 135717 1340 136283
rect 298660 135717 298854 136283
rect 1066 134629 1340 135195
rect 298660 134629 298854 135195
rect 1066 133541 1340 134107
rect 298660 133541 298854 134107
rect 1066 132453 1340 133019
rect 298660 132453 298854 133019
rect 1066 131365 1340 131931
rect 298660 131365 298854 131931
rect 1066 130277 1340 130843
rect 298660 130277 298854 130843
rect 1066 129189 1340 129755
rect 298660 129189 298854 129755
rect 1066 128101 1340 128667
rect 298660 128101 298854 128667
rect 1066 127013 1340 127579
rect 298660 127013 298854 127579
rect 1066 125925 1340 126491
rect 298660 125925 298854 126491
rect 1066 124837 1340 125403
rect 298660 124837 298854 125403
rect 1066 123749 1340 124315
rect 298660 123749 298854 124315
rect 1066 122661 1340 123227
rect 298660 122661 298854 123227
rect 1066 121573 1340 122139
rect 298660 121573 298854 122139
rect 1066 120485 1340 121051
rect 298660 120485 298854 121051
rect 1066 119397 1340 119963
rect 298660 119397 298854 119963
rect 1066 118309 1340 118875
rect 298660 118309 298854 118875
rect 1066 117221 1340 117787
rect 298660 117221 298854 117787
rect 1066 116133 1340 116699
rect 298660 116133 298854 116699
rect 1066 115045 1340 115611
rect 298660 115045 298854 115611
rect 1066 113957 1340 114523
rect 298660 113957 298854 114523
rect 1066 112869 1340 113435
rect 298660 112869 298854 113435
rect 1066 111781 1340 112347
rect 298660 111781 298854 112347
rect 1066 110693 1340 111259
rect 298660 110693 298854 111259
rect 1066 109605 1340 110171
rect 298660 109605 298854 110171
rect 1066 108517 1340 109083
rect 298660 108517 298854 109083
rect 1066 107429 1340 107995
rect 298660 107429 298854 107995
rect 1066 106341 1340 106907
rect 298660 106341 298854 106907
rect 1066 105253 1340 105819
rect 298660 105253 298854 105819
rect 1066 104165 1340 104731
rect 298660 104165 298854 104731
rect 1066 103077 1340 103643
rect 298660 103077 298854 103643
rect 1066 101989 1340 102555
rect 298660 101989 298854 102555
rect 1066 100901 1340 101467
rect 298660 100901 298854 101467
rect 1066 99813 1340 100379
rect 298660 99813 298854 100379
rect 1066 98725 1340 99291
rect 298660 98725 298854 99291
rect 1066 97637 1340 98203
rect 298660 97637 298854 98203
rect 1066 96549 1340 97115
rect 298660 96549 298854 97115
rect 1066 95461 1340 96027
rect 298660 95461 298854 96027
rect 1066 94373 1340 94939
rect 298660 94373 298854 94939
rect 1066 93285 1340 93851
rect 298660 93285 298854 93851
rect 1066 92197 1340 92763
rect 298660 92197 298854 92763
rect 1066 91109 1340 91675
rect 298660 91109 298854 91675
rect 1066 90021 1340 90587
rect 298660 90021 298854 90587
rect 1066 88933 1340 89499
rect 298660 88933 298854 89499
rect 1066 87845 1340 88411
rect 298660 87845 298854 88411
rect 1066 86757 1340 87323
rect 298660 86757 298854 87323
rect 1066 85669 1340 86235
rect 298660 85669 298854 86235
rect 1066 84581 1340 85147
rect 298660 84581 298854 85147
rect 1066 83493 1340 84059
rect 298660 83493 298854 84059
rect 1066 82405 1340 82971
rect 298660 82405 298854 82971
rect 1066 81317 1340 81883
rect 298660 81317 298854 81883
rect 1066 80229 1340 80795
rect 298660 80229 298854 80795
rect 1066 79141 1340 79707
rect 298660 79141 298854 79707
rect 1066 78053 1340 78619
rect 298660 78053 298854 78619
rect 1066 76965 1340 77531
rect 298660 76965 298854 77531
rect 1066 75877 1340 76443
rect 298660 75877 298854 76443
rect 1066 74789 1340 75355
rect 298660 74789 298854 75355
rect 1066 73701 1340 74267
rect 298660 73701 298854 74267
rect 1066 72613 1340 73179
rect 298660 72613 298854 73179
rect 1066 71525 1340 72091
rect 298660 71525 298854 72091
rect 1066 70437 1340 71003
rect 298660 70437 298854 71003
rect 1066 69349 1340 69915
rect 298660 69349 298854 69915
rect 1066 68261 1340 68827
rect 298660 68261 298854 68827
rect 1066 67173 1340 67739
rect 298660 67173 298854 67739
rect 1066 66085 1340 66651
rect 298660 66085 298854 66651
rect 1066 64997 1340 65563
rect 298660 64997 298854 65563
rect 1066 63909 1340 64475
rect 298660 63909 298854 64475
rect 1066 62821 1340 63387
rect 298660 62821 298854 63387
rect 1066 61733 1340 62299
rect 298660 61733 298854 62299
rect 1066 60645 1340 61211
rect 298660 60645 298854 61211
rect 1066 59557 1340 60123
rect 298660 59557 298854 60123
rect 1066 58469 1340 59035
rect 298660 58469 298854 59035
rect 1066 57381 1340 57947
rect 298660 57381 298854 57947
rect 1066 56293 1340 56859
rect 298660 56293 298854 56859
rect 1066 55205 1340 55771
rect 298660 55205 298854 55771
rect 1066 54117 1340 54683
rect 298660 54117 298854 54683
rect 1066 53029 1340 53595
rect 298660 53029 298854 53595
rect 1066 51941 1340 52507
rect 298660 51941 298854 52507
rect 1066 50853 1340 51419
rect 298660 50853 298854 51419
rect 1066 49765 1340 50331
rect 298660 49765 298854 50331
rect 1066 48677 1340 49243
rect 298660 48677 298854 49243
rect 1066 47589 1340 48155
rect 298660 47589 298854 48155
rect 1066 46501 1340 47067
rect 298660 46501 298854 47067
rect 1066 45413 1340 45979
rect 298660 45413 298854 45979
rect 1066 44325 1340 44891
rect 298660 44325 298854 44891
rect 1066 43237 1340 43803
rect 298660 43237 298854 43803
rect 1066 42149 1340 42715
rect 298660 42149 298854 42715
rect 1066 41061 1340 41627
rect 298660 41061 298854 41627
rect 1066 39973 1340 40539
rect 298660 39973 298854 40539
rect 1066 38885 1340 39451
rect 298660 38885 298854 39451
rect 1066 37797 1340 38363
rect 298660 37797 298854 38363
rect 1066 36709 1340 37275
rect 298660 36709 298854 37275
rect 1066 35621 1340 36187
rect 298660 35621 298854 36187
rect 1066 34533 1340 35099
rect 298660 34533 298854 35099
rect 1066 33445 1340 34011
rect 298660 33445 298854 34011
rect 1066 32357 1340 32923
rect 298660 32357 298854 32923
rect 1066 31269 1340 31835
rect 298660 31269 298854 31835
rect 1066 30181 1340 30747
rect 298660 30181 298854 30747
rect 1066 29093 1340 29659
rect 298660 29093 298854 29659
rect 1066 28005 1340 28571
rect 298660 28005 298854 28571
rect 1066 26917 1340 27483
rect 298660 26917 298854 27483
rect 1066 25829 1340 26395
rect 298660 25829 298854 26395
rect 1066 24741 1340 25307
rect 298660 24741 298854 25307
rect 1066 23653 1340 24219
rect 298660 23653 298854 24219
rect 1066 22565 1340 23131
rect 298660 22565 298854 23131
rect 1066 21477 1340 22043
rect 298660 21477 298854 22043
rect 1066 20389 1340 20955
rect 298660 20389 298854 20955
rect 1066 19301 1340 19867
rect 298660 19301 298854 19867
rect 1066 18213 1340 18779
rect 298660 18213 298854 18779
rect 1066 17125 1340 17691
rect 298660 17125 298854 17691
rect 1066 16037 1340 16603
rect 298660 16037 298854 16603
rect 1066 14949 1340 15515
rect 298660 14949 298854 15515
rect 1066 13861 1340 14427
rect 298660 13861 298854 14427
rect 1066 12773 1340 13339
rect 298660 12773 298854 13339
rect 1066 11685 1340 12251
rect 298660 11685 298854 12251
rect 1066 10597 1340 11163
rect 298660 10597 298854 11163
rect 1066 9509 1340 10075
rect 298660 9509 298854 10075
rect 1066 8421 1340 8987
rect 298660 8421 298854 8987
rect 1066 7333 1340 7899
rect 298660 7333 298854 7899
rect 1066 6245 1340 6811
rect 298660 6245 298854 6811
rect 1066 5157 1340 5723
rect 298660 5157 298854 5723
rect 1066 4069 1340 4635
rect 298660 4069 298854 4635
rect 1066 2981 1340 3547
rect 298660 2981 298854 3547
rect 1066 2138 1340 2459
rect 298660 2138 298854 2459
<< pwell >>
rect 1133 297551 1167 297585
rect 298753 297551 298787 297585
rect 1133 296463 1167 296497
rect 298753 296463 298787 296497
rect 1133 295375 1167 295409
rect 298753 295375 298787 295409
rect 1133 294287 1167 294321
rect 298753 294287 298787 294321
rect 1133 293199 1167 293233
rect 298753 293199 298787 293233
rect 1133 292111 1167 292145
rect 298753 292111 298787 292145
rect 1133 291023 1167 291057
rect 298753 291023 298787 291057
rect 1133 289935 1167 289969
rect 298753 289935 298787 289969
rect 1133 288847 1167 288881
rect 298753 288847 298787 288881
rect 1133 287759 1167 287793
rect 298753 287759 298787 287793
rect 1133 286671 1167 286705
rect 298753 286671 298787 286705
rect 1133 285583 1167 285617
rect 298753 285583 298787 285617
rect 1133 284495 1167 284529
rect 298753 284495 298787 284529
rect 1133 283407 1167 283441
rect 298753 283407 298787 283441
rect 1133 282319 1167 282353
rect 298753 282319 298787 282353
rect 1133 281231 1167 281265
rect 298753 281231 298787 281265
rect 1133 280143 1167 280177
rect 298753 280143 298787 280177
rect 1133 279055 1167 279089
rect 298753 279055 298787 279089
rect 1133 277967 1167 278001
rect 298753 277967 298787 278001
rect 1133 276879 1167 276913
rect 298753 276879 298787 276913
rect 1133 275791 1167 275825
rect 298753 275791 298787 275825
rect 1133 274703 1167 274737
rect 298753 274703 298787 274737
rect 1133 273615 1167 273649
rect 298753 273615 298787 273649
rect 1133 272527 1167 272561
rect 298753 272527 298787 272561
rect 1133 271439 1167 271473
rect 298753 271439 298787 271473
rect 1133 270351 1167 270385
rect 298753 270351 298787 270385
rect 1133 269263 1167 269297
rect 298753 269263 298787 269297
rect 1133 268175 1167 268209
rect 298753 268175 298787 268209
rect 1133 267087 1167 267121
rect 298753 267087 298787 267121
rect 1133 265999 1167 266033
rect 298753 265999 298787 266033
rect 1133 264911 1167 264945
rect 298753 264911 298787 264945
rect 1133 263823 1167 263857
rect 298753 263823 298787 263857
rect 1133 262735 1167 262769
rect 298753 262735 298787 262769
rect 1133 261647 1167 261681
rect 298753 261647 298787 261681
rect 1133 260559 1167 260593
rect 298753 260559 298787 260593
rect 1133 259471 1167 259505
rect 298753 259471 298787 259505
rect 1133 258383 1167 258417
rect 298753 258383 298787 258417
rect 1133 257295 1167 257329
rect 298753 257295 298787 257329
rect 1133 256207 1167 256241
rect 298753 256207 298787 256241
rect 1133 255119 1167 255153
rect 298753 255119 298787 255153
rect 1133 254031 1167 254065
rect 298753 254031 298787 254065
rect 1133 252943 1167 252977
rect 298753 252943 298787 252977
rect 1133 251855 1167 251889
rect 298753 251855 298787 251889
rect 1133 250767 1167 250801
rect 298753 250767 298787 250801
rect 1133 249679 1167 249713
rect 298753 249679 298787 249713
rect 1133 248591 1167 248625
rect 298753 248591 298787 248625
rect 1133 247503 1167 247537
rect 298753 247503 298787 247537
rect 1133 246415 1167 246449
rect 298753 246415 298787 246449
rect 1133 245327 1167 245361
rect 298753 245327 298787 245361
rect 1133 244239 1167 244273
rect 298753 244239 298787 244273
rect 1133 243151 1167 243185
rect 298753 243151 298787 243185
rect 1133 242063 1167 242097
rect 298753 242063 298787 242097
rect 1133 240975 1167 241009
rect 298753 240975 298787 241009
rect 1133 239887 1167 239921
rect 298753 239887 298787 239921
rect 1133 238799 1167 238833
rect 298753 238799 298787 238833
rect 1133 237711 1167 237745
rect 298753 237711 298787 237745
rect 1133 236623 1167 236657
rect 298753 236623 298787 236657
rect 1133 235535 1167 235569
rect 298753 235535 298787 235569
rect 1133 234447 1167 234481
rect 298753 234447 298787 234481
rect 1133 233359 1167 233393
rect 298753 233359 298787 233393
rect 1133 232271 1167 232305
rect 298753 232271 298787 232305
rect 1133 231183 1167 231217
rect 298753 231183 298787 231217
rect 1133 230095 1167 230129
rect 298753 230095 298787 230129
rect 1133 229007 1167 229041
rect 298753 229007 298787 229041
rect 1133 227919 1167 227953
rect 298753 227919 298787 227953
rect 1133 226831 1167 226865
rect 298753 226831 298787 226865
rect 1133 225743 1167 225777
rect 298753 225743 298787 225777
rect 1133 224655 1167 224689
rect 298753 224655 298787 224689
rect 1133 223567 1167 223601
rect 298753 223567 298787 223601
rect 1133 222479 1167 222513
rect 298753 222479 298787 222513
rect 1133 221391 1167 221425
rect 298753 221391 298787 221425
rect 1133 220303 1167 220337
rect 298753 220303 298787 220337
rect 1133 219215 1167 219249
rect 298753 219215 298787 219249
rect 1133 218127 1167 218161
rect 298753 218127 298787 218161
rect 1133 217039 1167 217073
rect 298753 217039 298787 217073
rect 1133 215951 1167 215985
rect 298753 215951 298787 215985
rect 1133 214863 1167 214897
rect 298753 214863 298787 214897
rect 1133 213775 1167 213809
rect 298753 213775 298787 213809
rect 1133 212687 1167 212721
rect 298753 212687 298787 212721
rect 1133 211599 1167 211633
rect 298753 211599 298787 211633
rect 1133 210511 1167 210545
rect 298753 210511 298787 210545
rect 1133 209423 1167 209457
rect 298753 209423 298787 209457
rect 1133 208335 1167 208369
rect 298753 208335 298787 208369
rect 1133 207247 1167 207281
rect 298753 207247 298787 207281
rect 1133 206159 1167 206193
rect 298753 206159 298787 206193
rect 1133 205071 1167 205105
rect 298753 205071 298787 205105
rect 1133 203983 1167 204017
rect 298753 203983 298787 204017
rect 1133 202895 1167 202929
rect 298753 202895 298787 202929
rect 1133 201807 1167 201841
rect 298753 201807 298787 201841
rect 1133 200719 1167 200753
rect 298753 200719 298787 200753
rect 1133 199631 1167 199665
rect 298753 199631 298787 199665
rect 1133 198543 1167 198577
rect 298753 198543 298787 198577
rect 1133 197455 1167 197489
rect 298753 197455 298787 197489
rect 1133 196367 1167 196401
rect 298753 196367 298787 196401
rect 1133 195279 1167 195313
rect 298753 195279 298787 195313
rect 1133 194191 1167 194225
rect 298753 194191 298787 194225
rect 1133 193103 1167 193137
rect 298753 193103 298787 193137
rect 1133 192015 1167 192049
rect 298753 192015 298787 192049
rect 1133 190927 1167 190961
rect 298753 190927 298787 190961
rect 1133 189839 1167 189873
rect 298753 189839 298787 189873
rect 1133 188751 1167 188785
rect 298753 188751 298787 188785
rect 1133 187663 1167 187697
rect 298753 187663 298787 187697
rect 1133 186575 1167 186609
rect 298753 186575 298787 186609
rect 1133 185487 1167 185521
rect 298753 185487 298787 185521
rect 1133 184399 1167 184433
rect 298753 184399 298787 184433
rect 1133 183311 1167 183345
rect 298753 183311 298787 183345
rect 1133 182223 1167 182257
rect 298753 182223 298787 182257
rect 1133 181135 1167 181169
rect 298753 181135 298787 181169
rect 1133 180047 1167 180081
rect 298753 180047 298787 180081
rect 1133 178959 1167 178993
rect 298753 178959 298787 178993
rect 1133 177871 1167 177905
rect 298753 177871 298787 177905
rect 1133 176783 1167 176817
rect 298753 176783 298787 176817
rect 1133 175695 1167 175729
rect 298753 175695 298787 175729
rect 1133 174607 1167 174641
rect 298753 174607 298787 174641
rect 1133 173519 1167 173553
rect 298753 173519 298787 173553
rect 1133 172431 1167 172465
rect 298753 172431 298787 172465
rect 1133 171343 1167 171377
rect 298753 171343 298787 171377
rect 1133 170255 1167 170289
rect 298753 170255 298787 170289
rect 1133 169167 1167 169201
rect 298753 169167 298787 169201
rect 1133 168079 1167 168113
rect 298753 168079 298787 168113
rect 1133 166991 1167 167025
rect 298753 166991 298787 167025
rect 1133 165903 1167 165937
rect 298753 165903 298787 165937
rect 1133 164815 1167 164849
rect 298753 164815 298787 164849
rect 1133 163727 1167 163761
rect 298753 163727 298787 163761
rect 1133 162639 1167 162673
rect 298753 162639 298787 162673
rect 1133 161551 1167 161585
rect 298753 161551 298787 161585
rect 1133 160463 1167 160497
rect 298753 160463 298787 160497
rect 1133 159375 1167 159409
rect 298753 159375 298787 159409
rect 1133 158287 1167 158321
rect 298753 158287 298787 158321
rect 1133 157199 1167 157233
rect 298753 157199 298787 157233
rect 1133 156111 1167 156145
rect 298753 156111 298787 156145
rect 1133 155023 1167 155057
rect 298753 155023 298787 155057
rect 1133 153935 1167 153969
rect 298753 153935 298787 153969
rect 1133 152847 1167 152881
rect 298753 152847 298787 152881
rect 1133 151759 1167 151793
rect 298753 151759 298787 151793
rect 1133 150671 1167 150705
rect 298753 150671 298787 150705
rect 1133 149583 1167 149617
rect 298753 149583 298787 149617
rect 1133 148495 1167 148529
rect 298753 148495 298787 148529
rect 1133 147407 1167 147441
rect 298753 147407 298787 147441
rect 1133 146319 1167 146353
rect 298753 146319 298787 146353
rect 1133 145231 1167 145265
rect 298753 145231 298787 145265
rect 1133 144143 1167 144177
rect 298753 144143 298787 144177
rect 1133 143055 1167 143089
rect 298753 143055 298787 143089
rect 1133 141967 1167 142001
rect 298753 141967 298787 142001
rect 1133 140879 1167 140913
rect 298753 140879 298787 140913
rect 1133 139791 1167 139825
rect 298753 139791 298787 139825
rect 1133 138703 1167 138737
rect 298753 138703 298787 138737
rect 1133 137615 1167 137649
rect 298753 137615 298787 137649
rect 1133 136527 1167 136561
rect 298753 136527 298787 136561
rect 1133 135439 1167 135473
rect 298753 135439 298787 135473
rect 1133 134351 1167 134385
rect 298753 134351 298787 134385
rect 1133 133263 1167 133297
rect 298753 133263 298787 133297
rect 1133 132175 1167 132209
rect 298753 132175 298787 132209
rect 1133 131087 1167 131121
rect 298753 131087 298787 131121
rect 1133 129999 1167 130033
rect 298753 129999 298787 130033
rect 1133 128911 1167 128945
rect 298753 128911 298787 128945
rect 1133 127823 1167 127857
rect 298753 127823 298787 127857
rect 1133 126735 1167 126769
rect 298753 126735 298787 126769
rect 1133 125647 1167 125681
rect 298753 125647 298787 125681
rect 1133 124559 1167 124593
rect 298753 124559 298787 124593
rect 1133 123471 1167 123505
rect 298753 123471 298787 123505
rect 1133 122383 1167 122417
rect 298753 122383 298787 122417
rect 1133 121295 1167 121329
rect 298753 121295 298787 121329
rect 1133 120207 1167 120241
rect 298753 120207 298787 120241
rect 1133 119119 1167 119153
rect 298753 119119 298787 119153
rect 1133 118031 1167 118065
rect 298753 118031 298787 118065
rect 1133 116943 1167 116977
rect 298753 116943 298787 116977
rect 1133 115855 1167 115889
rect 298753 115855 298787 115889
rect 1133 114767 1167 114801
rect 298753 114767 298787 114801
rect 1133 113679 1167 113713
rect 298753 113679 298787 113713
rect 1133 112591 1167 112625
rect 298753 112591 298787 112625
rect 1133 111503 1167 111537
rect 298753 111503 298787 111537
rect 1133 110415 1167 110449
rect 298753 110415 298787 110449
rect 1133 109327 1167 109361
rect 298753 109327 298787 109361
rect 1133 108239 1167 108273
rect 298753 108239 298787 108273
rect 1133 107151 1167 107185
rect 298753 107151 298787 107185
rect 1133 106063 1167 106097
rect 298753 106063 298787 106097
rect 1133 104975 1167 105009
rect 298753 104975 298787 105009
rect 1133 103887 1167 103921
rect 298753 103887 298787 103921
rect 1133 102799 1167 102833
rect 298753 102799 298787 102833
rect 1133 101711 1167 101745
rect 298753 101711 298787 101745
rect 1133 100623 1167 100657
rect 298753 100623 298787 100657
rect 1133 99535 1167 99569
rect 298753 99535 298787 99569
rect 1133 98447 1167 98481
rect 298753 98447 298787 98481
rect 1133 97359 1167 97393
rect 298753 97359 298787 97393
rect 1133 96271 1167 96305
rect 298753 96271 298787 96305
rect 1133 95183 1167 95217
rect 298753 95183 298787 95217
rect 1133 94095 1167 94129
rect 298753 94095 298787 94129
rect 1133 93007 1167 93041
rect 298753 93007 298787 93041
rect 1133 91919 1167 91953
rect 298753 91919 298787 91953
rect 1133 90831 1167 90865
rect 298753 90831 298787 90865
rect 1133 89743 1167 89777
rect 298753 89743 298787 89777
rect 1133 88655 1167 88689
rect 298753 88655 298787 88689
rect 1133 87567 1167 87601
rect 298753 87567 298787 87601
rect 1133 86479 1167 86513
rect 298753 86479 298787 86513
rect 1133 85391 1167 85425
rect 298753 85391 298787 85425
rect 1133 84303 1167 84337
rect 298753 84303 298787 84337
rect 1133 83215 1167 83249
rect 298753 83215 298787 83249
rect 1133 82127 1167 82161
rect 298753 82127 298787 82161
rect 1133 81039 1167 81073
rect 298753 81039 298787 81073
rect 1133 79951 1167 79985
rect 298753 79951 298787 79985
rect 1133 78863 1167 78897
rect 298753 78863 298787 78897
rect 1133 77775 1167 77809
rect 298753 77775 298787 77809
rect 1133 76687 1167 76721
rect 298753 76687 298787 76721
rect 1133 75599 1167 75633
rect 298753 75599 298787 75633
rect 1133 74511 1167 74545
rect 298753 74511 298787 74545
rect 1133 73423 1167 73457
rect 298753 73423 298787 73457
rect 1133 72335 1167 72369
rect 298753 72335 298787 72369
rect 1133 71247 1167 71281
rect 298753 71247 298787 71281
rect 1133 70159 1167 70193
rect 298753 70159 298787 70193
rect 1133 69071 1167 69105
rect 298753 69071 298787 69105
rect 1133 67983 1167 68017
rect 298753 67983 298787 68017
rect 1133 66895 1167 66929
rect 298753 66895 298787 66929
rect 1133 65807 1167 65841
rect 298753 65807 298787 65841
rect 1133 64719 1167 64753
rect 298753 64719 298787 64753
rect 1133 63631 1167 63665
rect 298753 63631 298787 63665
rect 1133 62543 1167 62577
rect 298753 62543 298787 62577
rect 1133 61455 1167 61489
rect 298753 61455 298787 61489
rect 1133 60367 1167 60401
rect 298753 60367 298787 60401
rect 1133 59279 1167 59313
rect 298753 59279 298787 59313
rect 1133 58191 1167 58225
rect 298753 58191 298787 58225
rect 1133 57103 1167 57137
rect 298753 57103 298787 57137
rect 1133 56015 1167 56049
rect 298753 56015 298787 56049
rect 1133 54927 1167 54961
rect 298753 54927 298787 54961
rect 1133 53839 1167 53873
rect 298753 53839 298787 53873
rect 1133 52751 1167 52785
rect 298753 52751 298787 52785
rect 1133 51663 1167 51697
rect 298753 51663 298787 51697
rect 1133 50575 1167 50609
rect 298753 50575 298787 50609
rect 1133 49487 1167 49521
rect 298753 49487 298787 49521
rect 1133 48399 1167 48433
rect 298753 48399 298787 48433
rect 1133 47311 1167 47345
rect 298753 47311 298787 47345
rect 1133 46223 1167 46257
rect 298753 46223 298787 46257
rect 1133 45135 1167 45169
rect 298753 45135 298787 45169
rect 1133 44047 1167 44081
rect 298753 44047 298787 44081
rect 1133 42959 1167 42993
rect 298753 42959 298787 42993
rect 1133 41871 1167 41905
rect 298753 41871 298787 41905
rect 1133 40783 1167 40817
rect 298753 40783 298787 40817
rect 1133 39695 1167 39729
rect 298753 39695 298787 39729
rect 1133 38607 1167 38641
rect 298753 38607 298787 38641
rect 1133 37519 1167 37553
rect 298753 37519 298787 37553
rect 1133 36431 1167 36465
rect 298753 36431 298787 36465
rect 1133 35343 1167 35377
rect 298753 35343 298787 35377
rect 1133 34255 1167 34289
rect 298753 34255 298787 34289
rect 1133 33167 1167 33201
rect 298753 33167 298787 33201
rect 1133 32079 1167 32113
rect 298753 32079 298787 32113
rect 1133 30991 1167 31025
rect 298753 30991 298787 31025
rect 1133 29903 1167 29937
rect 298753 29903 298787 29937
rect 1133 28815 1167 28849
rect 298753 28815 298787 28849
rect 1133 27727 1167 27761
rect 298753 27727 298787 27761
rect 1133 26639 1167 26673
rect 298753 26639 298787 26673
rect 1133 25551 1167 25585
rect 298753 25551 298787 25585
rect 1133 24463 1167 24497
rect 298753 24463 298787 24497
rect 1133 23375 1167 23409
rect 298753 23375 298787 23409
rect 1133 22287 1167 22321
rect 298753 22287 298787 22321
rect 1133 21199 1167 21233
rect 298753 21199 298787 21233
rect 1133 20111 1167 20145
rect 298753 20111 298787 20145
rect 1133 19023 1167 19057
rect 298753 19023 298787 19057
rect 1133 17935 1167 17969
rect 298753 17935 298787 17969
rect 1133 16847 1167 16881
rect 298753 16847 298787 16881
rect 1133 15759 1167 15793
rect 298753 15759 298787 15793
rect 1133 14671 1167 14705
rect 298753 14671 298787 14705
rect 1133 13583 1167 13617
rect 298753 13583 298787 13617
rect 1133 12495 1167 12529
rect 298753 12495 298787 12529
rect 1133 11407 1167 11441
rect 298753 11407 298787 11441
rect 1133 10319 1167 10353
rect 298753 10319 298787 10353
rect 1133 9231 1167 9265
rect 298753 9231 298787 9265
rect 1133 8143 1167 8177
rect 298753 8143 298787 8177
rect 1133 7055 1167 7089
rect 298753 7055 298787 7089
rect 1133 5967 1167 6001
rect 298753 5967 298787 6001
rect 1133 4879 1167 4913
rect 298753 4879 298787 4913
rect 1133 3791 1167 3825
rect 298753 3791 298787 3825
rect 1133 2703 1167 2737
rect 298753 2703 298787 2737
<< locali >>
rect 1104 297551 1133 297585
rect 1167 297551 1225 297585
rect 1259 297551 1317 297585
rect 1121 297401 1340 297551
rect 1121 297293 1225 297401
rect 1259 297259 1340 297367
rect 1121 297041 1340 297259
rect 1104 297007 1133 297041
rect 1167 297007 1225 297041
rect 1259 297007 1317 297041
rect 1121 296789 1340 297007
rect 1121 296647 1225 296755
rect 1259 296681 1340 296789
rect 1121 296497 1340 296647
rect 1104 296463 1133 296497
rect 1167 296463 1225 296497
rect 1259 296463 1317 296497
rect 1121 296313 1340 296463
rect 1121 296205 1225 296313
rect 1259 296171 1340 296279
rect 1121 295953 1340 296171
rect 1104 295919 1133 295953
rect 1167 295919 1225 295953
rect 1259 295919 1317 295953
rect 1121 295701 1340 295919
rect 1121 295559 1225 295667
rect 1259 295593 1340 295701
rect 1121 295409 1340 295559
rect 1104 295375 1133 295409
rect 1167 295375 1225 295409
rect 1259 295375 1317 295409
rect 1121 295225 1340 295375
rect 1121 295117 1225 295225
rect 1259 295083 1340 295191
rect 1121 294865 1340 295083
rect 1104 294831 1133 294865
rect 1167 294831 1225 294865
rect 1259 294831 1317 294865
rect 1121 294613 1340 294831
rect 1121 294471 1225 294579
rect 1259 294505 1340 294613
rect 1121 294321 1340 294471
rect 1104 294287 1133 294321
rect 1167 294287 1225 294321
rect 1259 294287 1317 294321
rect 1121 294137 1340 294287
rect 1121 294029 1225 294137
rect 1259 293995 1340 294103
rect 1121 293777 1340 293995
rect 1104 293743 1133 293777
rect 1167 293743 1225 293777
rect 1259 293743 1317 293777
rect 1121 293525 1340 293743
rect 1121 293383 1225 293491
rect 1259 293417 1340 293525
rect 1121 293233 1340 293383
rect 1104 293199 1133 293233
rect 1167 293199 1225 293233
rect 1259 293199 1317 293233
rect 1121 293049 1340 293199
rect 1121 292941 1225 293049
rect 1259 292907 1340 293015
rect 1121 292689 1340 292907
rect 1104 292655 1133 292689
rect 1167 292655 1225 292689
rect 1259 292655 1317 292689
rect 1121 292437 1340 292655
rect 1121 292295 1225 292403
rect 1259 292329 1340 292437
rect 1121 292145 1340 292295
rect 1104 292111 1133 292145
rect 1167 292111 1225 292145
rect 1259 292111 1317 292145
rect 1121 291961 1340 292111
rect 1121 291853 1225 291961
rect 1259 291819 1340 291927
rect 1121 291601 1340 291819
rect 1104 291567 1133 291601
rect 1167 291567 1225 291601
rect 1259 291567 1317 291601
rect 1121 291349 1340 291567
rect 1121 291207 1225 291315
rect 1259 291241 1340 291349
rect 1121 291057 1340 291207
rect 1104 291023 1133 291057
rect 1167 291023 1225 291057
rect 1259 291023 1317 291057
rect 1121 290873 1340 291023
rect 1121 290765 1225 290873
rect 1259 290731 1340 290839
rect 1121 290513 1340 290731
rect 1104 290479 1133 290513
rect 1167 290479 1225 290513
rect 1259 290479 1317 290513
rect 1121 290261 1340 290479
rect 1121 290119 1225 290227
rect 1259 290153 1340 290261
rect 1121 289969 1340 290119
rect 1104 289935 1133 289969
rect 1167 289935 1225 289969
rect 1259 289935 1317 289969
rect 1121 289785 1340 289935
rect 1121 289677 1225 289785
rect 1259 289643 1340 289751
rect 1121 289425 1340 289643
rect 1104 289391 1133 289425
rect 1167 289391 1225 289425
rect 1259 289391 1317 289425
rect 1121 289173 1340 289391
rect 1121 289031 1225 289139
rect 1259 289065 1340 289173
rect 1121 288881 1340 289031
rect 1104 288847 1133 288881
rect 1167 288847 1225 288881
rect 1259 288847 1317 288881
rect 1121 288697 1340 288847
rect 1121 288589 1225 288697
rect 1259 288555 1340 288663
rect 1121 288337 1340 288555
rect 1104 288303 1133 288337
rect 1167 288303 1225 288337
rect 1259 288303 1317 288337
rect 1121 288085 1340 288303
rect 1121 287943 1225 288051
rect 1259 287977 1340 288085
rect 1121 287793 1340 287943
rect 1104 287759 1133 287793
rect 1167 287759 1225 287793
rect 1259 287759 1317 287793
rect 1121 287609 1340 287759
rect 1121 287501 1225 287609
rect 1259 287467 1340 287575
rect 1121 287249 1340 287467
rect 1104 287215 1133 287249
rect 1167 287215 1225 287249
rect 1259 287215 1317 287249
rect 1121 286997 1340 287215
rect 1121 286855 1225 286963
rect 1259 286889 1340 286997
rect 1121 286705 1340 286855
rect 1104 286671 1133 286705
rect 1167 286671 1225 286705
rect 1259 286671 1317 286705
rect 1121 286521 1340 286671
rect 1121 286413 1225 286521
rect 1259 286379 1340 286487
rect 1121 286161 1340 286379
rect 1104 286127 1133 286161
rect 1167 286127 1225 286161
rect 1259 286127 1317 286161
rect 1121 285909 1340 286127
rect 1121 285767 1225 285875
rect 1259 285801 1340 285909
rect 1121 285617 1340 285767
rect 1104 285583 1133 285617
rect 1167 285583 1225 285617
rect 1259 285583 1317 285617
rect 1121 285433 1340 285583
rect 1121 285325 1225 285433
rect 1259 285291 1340 285399
rect 1121 285073 1340 285291
rect 1104 285039 1133 285073
rect 1167 285039 1225 285073
rect 1259 285039 1317 285073
rect 1121 284821 1340 285039
rect 1121 284679 1225 284787
rect 1259 284713 1340 284821
rect 1121 284529 1340 284679
rect 1104 284495 1133 284529
rect 1167 284495 1225 284529
rect 1259 284495 1317 284529
rect 1121 284345 1340 284495
rect 1121 284237 1225 284345
rect 1259 284203 1340 284311
rect 1121 283985 1340 284203
rect 1104 283951 1133 283985
rect 1167 283951 1225 283985
rect 1259 283951 1317 283985
rect 1121 283733 1340 283951
rect 1121 283591 1225 283699
rect 1259 283625 1340 283733
rect 1121 283441 1340 283591
rect 1104 283407 1133 283441
rect 1167 283407 1225 283441
rect 1259 283407 1317 283441
rect 1121 283257 1340 283407
rect 1121 283149 1225 283257
rect 1259 283115 1340 283223
rect 1121 282897 1340 283115
rect 1104 282863 1133 282897
rect 1167 282863 1225 282897
rect 1259 282863 1317 282897
rect 1121 282645 1340 282863
rect 1121 282503 1225 282611
rect 1259 282537 1340 282645
rect 1121 282353 1340 282503
rect 1104 282319 1133 282353
rect 1167 282319 1225 282353
rect 1259 282319 1317 282353
rect 1121 282169 1340 282319
rect 1121 282061 1225 282169
rect 1259 282027 1340 282135
rect 1121 281809 1340 282027
rect 1104 281775 1133 281809
rect 1167 281775 1225 281809
rect 1259 281775 1317 281809
rect 1121 281557 1340 281775
rect 1121 281415 1225 281523
rect 1259 281449 1340 281557
rect 1121 281265 1340 281415
rect 1104 281231 1133 281265
rect 1167 281231 1225 281265
rect 1259 281231 1317 281265
rect 1121 281081 1340 281231
rect 1121 280973 1225 281081
rect 1259 280939 1340 281047
rect 1121 280721 1340 280939
rect 1104 280687 1133 280721
rect 1167 280687 1225 280721
rect 1259 280687 1317 280721
rect 1121 280469 1340 280687
rect 1121 280327 1225 280435
rect 1259 280361 1340 280469
rect 1121 280177 1340 280327
rect 1104 280143 1133 280177
rect 1167 280143 1225 280177
rect 1259 280143 1317 280177
rect 1121 279993 1340 280143
rect 1121 279885 1225 279993
rect 1259 279851 1340 279959
rect 1121 279633 1340 279851
rect 1104 279599 1133 279633
rect 1167 279599 1225 279633
rect 1259 279599 1317 279633
rect 1121 279381 1340 279599
rect 1121 279239 1225 279347
rect 1259 279273 1340 279381
rect 1121 279089 1340 279239
rect 1104 279055 1133 279089
rect 1167 279055 1225 279089
rect 1259 279055 1317 279089
rect 1121 278905 1340 279055
rect 1121 278797 1225 278905
rect 1259 278763 1340 278871
rect 1121 278545 1340 278763
rect 1104 278511 1133 278545
rect 1167 278511 1225 278545
rect 1259 278511 1317 278545
rect 1121 278293 1340 278511
rect 1121 278151 1225 278259
rect 1259 278185 1340 278293
rect 1121 278001 1340 278151
rect 1104 277967 1133 278001
rect 1167 277967 1225 278001
rect 1259 277967 1317 278001
rect 1121 277817 1340 277967
rect 1121 277709 1225 277817
rect 1259 277675 1340 277783
rect 1121 277457 1340 277675
rect 1104 277423 1133 277457
rect 1167 277423 1225 277457
rect 1259 277423 1317 277457
rect 1121 277205 1340 277423
rect 1121 277063 1225 277171
rect 1259 277097 1340 277205
rect 1121 276913 1340 277063
rect 1104 276879 1133 276913
rect 1167 276879 1225 276913
rect 1259 276879 1317 276913
rect 1121 276729 1340 276879
rect 1121 276621 1225 276729
rect 1259 276587 1340 276695
rect 1121 276369 1340 276587
rect 1104 276335 1133 276369
rect 1167 276335 1225 276369
rect 1259 276335 1317 276369
rect 1121 276117 1340 276335
rect 1121 275975 1225 276083
rect 1259 276009 1340 276117
rect 1121 275825 1340 275975
rect 1104 275791 1133 275825
rect 1167 275791 1225 275825
rect 1259 275791 1317 275825
rect 1121 275641 1340 275791
rect 1121 275533 1225 275641
rect 1259 275499 1340 275607
rect 1121 275281 1340 275499
rect 1104 275247 1133 275281
rect 1167 275247 1225 275281
rect 1259 275247 1317 275281
rect 1121 275029 1340 275247
rect 1121 274887 1225 274995
rect 1259 274921 1340 275029
rect 1121 274737 1340 274887
rect 1104 274703 1133 274737
rect 1167 274703 1225 274737
rect 1259 274703 1317 274737
rect 1121 274553 1340 274703
rect 1121 274445 1225 274553
rect 1259 274411 1340 274519
rect 1121 274193 1340 274411
rect 1104 274159 1133 274193
rect 1167 274159 1225 274193
rect 1259 274159 1317 274193
rect 1121 273941 1340 274159
rect 1121 273799 1225 273907
rect 1259 273833 1340 273941
rect 1121 273649 1340 273799
rect 1104 273615 1133 273649
rect 1167 273615 1225 273649
rect 1259 273615 1317 273649
rect 1121 273465 1340 273615
rect 1121 273357 1225 273465
rect 1259 273323 1340 273431
rect 1121 273105 1340 273323
rect 1104 273071 1133 273105
rect 1167 273071 1225 273105
rect 1259 273071 1317 273105
rect 1121 272853 1340 273071
rect 1121 272711 1225 272819
rect 1259 272745 1340 272853
rect 1121 272561 1340 272711
rect 1104 272527 1133 272561
rect 1167 272527 1225 272561
rect 1259 272527 1317 272561
rect 1121 272377 1340 272527
rect 1121 272269 1225 272377
rect 1259 272235 1340 272343
rect 1121 272017 1340 272235
rect 1104 271983 1133 272017
rect 1167 271983 1225 272017
rect 1259 271983 1317 272017
rect 1121 271765 1340 271983
rect 1121 271623 1225 271731
rect 1259 271657 1340 271765
rect 1121 271473 1340 271623
rect 1104 271439 1133 271473
rect 1167 271439 1225 271473
rect 1259 271439 1317 271473
rect 1121 271289 1340 271439
rect 1121 271181 1225 271289
rect 1259 271147 1340 271255
rect 1121 270929 1340 271147
rect 1104 270895 1133 270929
rect 1167 270895 1225 270929
rect 1259 270895 1317 270929
rect 1121 270677 1340 270895
rect 1121 270535 1225 270643
rect 1259 270569 1340 270677
rect 1121 270385 1340 270535
rect 1104 270351 1133 270385
rect 1167 270351 1225 270385
rect 1259 270351 1317 270385
rect 1121 270201 1340 270351
rect 1121 270093 1225 270201
rect 1259 270059 1340 270167
rect 1121 269841 1340 270059
rect 1104 269807 1133 269841
rect 1167 269807 1225 269841
rect 1259 269807 1317 269841
rect 1121 269589 1340 269807
rect 1121 269447 1225 269555
rect 1259 269481 1340 269589
rect 1121 269297 1340 269447
rect 1104 269263 1133 269297
rect 1167 269263 1225 269297
rect 1259 269263 1317 269297
rect 1121 269113 1340 269263
rect 1121 269005 1225 269113
rect 1259 268971 1340 269079
rect 1121 268753 1340 268971
rect 1104 268719 1133 268753
rect 1167 268719 1225 268753
rect 1259 268719 1317 268753
rect 1121 268501 1340 268719
rect 1121 268359 1225 268467
rect 1259 268393 1340 268501
rect 1121 268209 1340 268359
rect 1104 268175 1133 268209
rect 1167 268175 1225 268209
rect 1259 268175 1317 268209
rect 1121 268025 1340 268175
rect 1121 267917 1225 268025
rect 1259 267883 1340 267991
rect 1121 267665 1340 267883
rect 1104 267631 1133 267665
rect 1167 267631 1225 267665
rect 1259 267631 1317 267665
rect 1121 267413 1340 267631
rect 1121 267271 1225 267379
rect 1259 267305 1340 267413
rect 1121 267121 1340 267271
rect 1104 267087 1133 267121
rect 1167 267087 1225 267121
rect 1259 267087 1317 267121
rect 1121 266937 1340 267087
rect 1121 266829 1225 266937
rect 1259 266795 1340 266903
rect 1121 266577 1340 266795
rect 1104 266543 1133 266577
rect 1167 266543 1225 266577
rect 1259 266543 1317 266577
rect 1121 266325 1340 266543
rect 1121 266183 1225 266291
rect 1259 266217 1340 266325
rect 1121 266033 1340 266183
rect 1104 265999 1133 266033
rect 1167 265999 1225 266033
rect 1259 265999 1317 266033
rect 1121 265849 1340 265999
rect 1121 265741 1225 265849
rect 1259 265707 1340 265815
rect 1121 265489 1340 265707
rect 1104 265455 1133 265489
rect 1167 265455 1225 265489
rect 1259 265455 1317 265489
rect 1121 265237 1340 265455
rect 1121 265095 1225 265203
rect 1259 265129 1340 265237
rect 1121 264945 1340 265095
rect 1104 264911 1133 264945
rect 1167 264911 1225 264945
rect 1259 264911 1317 264945
rect 1121 264761 1340 264911
rect 1121 264653 1225 264761
rect 1259 264619 1340 264727
rect 1121 264401 1340 264619
rect 1104 264367 1133 264401
rect 1167 264367 1225 264401
rect 1259 264367 1317 264401
rect 1121 264149 1340 264367
rect 1121 264007 1225 264115
rect 1259 264041 1340 264149
rect 1121 263857 1340 264007
rect 1104 263823 1133 263857
rect 1167 263823 1225 263857
rect 1259 263823 1317 263857
rect 1121 263673 1340 263823
rect 1121 263565 1225 263673
rect 1259 263531 1340 263639
rect 1121 263313 1340 263531
rect 1104 263279 1133 263313
rect 1167 263279 1225 263313
rect 1259 263279 1317 263313
rect 1121 263061 1340 263279
rect 1121 262919 1225 263027
rect 1259 262953 1340 263061
rect 1121 262769 1340 262919
rect 1104 262735 1133 262769
rect 1167 262735 1225 262769
rect 1259 262735 1317 262769
rect 1121 262585 1340 262735
rect 1121 262477 1225 262585
rect 1259 262443 1340 262551
rect 1121 262225 1340 262443
rect 1104 262191 1133 262225
rect 1167 262191 1225 262225
rect 1259 262191 1317 262225
rect 1121 261973 1340 262191
rect 1121 261831 1225 261939
rect 1259 261865 1340 261973
rect 1121 261681 1340 261831
rect 1104 261647 1133 261681
rect 1167 261647 1225 261681
rect 1259 261647 1317 261681
rect 1121 261497 1340 261647
rect 1121 261389 1225 261497
rect 1259 261355 1340 261463
rect 1121 261137 1340 261355
rect 1104 261103 1133 261137
rect 1167 261103 1225 261137
rect 1259 261103 1317 261137
rect 1121 260885 1340 261103
rect 1121 260743 1225 260851
rect 1259 260777 1340 260885
rect 1121 260593 1340 260743
rect 1104 260559 1133 260593
rect 1167 260559 1225 260593
rect 1259 260559 1317 260593
rect 1121 260409 1340 260559
rect 1121 260301 1225 260409
rect 1259 260267 1340 260375
rect 1121 260049 1340 260267
rect 1104 260015 1133 260049
rect 1167 260015 1225 260049
rect 1259 260015 1317 260049
rect 1121 259797 1340 260015
rect 1121 259655 1225 259763
rect 1259 259689 1340 259797
rect 1121 259505 1340 259655
rect 1104 259471 1133 259505
rect 1167 259471 1225 259505
rect 1259 259471 1317 259505
rect 1121 259321 1340 259471
rect 1121 259213 1225 259321
rect 1259 259179 1340 259287
rect 1121 258961 1340 259179
rect 1104 258927 1133 258961
rect 1167 258927 1225 258961
rect 1259 258927 1317 258961
rect 1121 258709 1340 258927
rect 1121 258567 1225 258675
rect 1259 258601 1340 258709
rect 1121 258417 1340 258567
rect 1104 258383 1133 258417
rect 1167 258383 1225 258417
rect 1259 258383 1317 258417
rect 1121 258233 1340 258383
rect 1121 258125 1225 258233
rect 1259 258091 1340 258199
rect 1121 257873 1340 258091
rect 1104 257839 1133 257873
rect 1167 257839 1225 257873
rect 1259 257839 1317 257873
rect 1121 257621 1340 257839
rect 1121 257479 1225 257587
rect 1259 257513 1340 257621
rect 1121 257329 1340 257479
rect 1104 257295 1133 257329
rect 1167 257295 1225 257329
rect 1259 257295 1317 257329
rect 1121 257145 1340 257295
rect 1121 257037 1225 257145
rect 1259 257003 1340 257111
rect 1121 256785 1340 257003
rect 1104 256751 1133 256785
rect 1167 256751 1225 256785
rect 1259 256751 1317 256785
rect 1121 256533 1340 256751
rect 1121 256391 1225 256499
rect 1259 256425 1340 256533
rect 1121 256241 1340 256391
rect 1104 256207 1133 256241
rect 1167 256207 1225 256241
rect 1259 256207 1317 256241
rect 1121 256057 1340 256207
rect 1121 255949 1225 256057
rect 1259 255915 1340 256023
rect 1121 255697 1340 255915
rect 1104 255663 1133 255697
rect 1167 255663 1225 255697
rect 1259 255663 1317 255697
rect 1121 255445 1340 255663
rect 1121 255303 1225 255411
rect 1259 255337 1340 255445
rect 1121 255153 1340 255303
rect 1104 255119 1133 255153
rect 1167 255119 1225 255153
rect 1259 255119 1317 255153
rect 1121 254969 1340 255119
rect 1121 254861 1225 254969
rect 1259 254827 1340 254935
rect 1121 254609 1340 254827
rect 1104 254575 1133 254609
rect 1167 254575 1225 254609
rect 1259 254575 1317 254609
rect 1121 254357 1340 254575
rect 1121 254215 1225 254323
rect 1259 254249 1340 254357
rect 1121 254065 1340 254215
rect 1104 254031 1133 254065
rect 1167 254031 1225 254065
rect 1259 254031 1317 254065
rect 1121 253881 1340 254031
rect 1121 253773 1225 253881
rect 1259 253739 1340 253847
rect 1121 253521 1340 253739
rect 1104 253487 1133 253521
rect 1167 253487 1225 253521
rect 1259 253487 1317 253521
rect 1121 253269 1340 253487
rect 1121 253127 1225 253235
rect 1259 253161 1340 253269
rect 1121 252977 1340 253127
rect 1104 252943 1133 252977
rect 1167 252943 1225 252977
rect 1259 252943 1317 252977
rect 1121 252793 1340 252943
rect 1121 252685 1225 252793
rect 1259 252651 1340 252759
rect 1121 252433 1340 252651
rect 1104 252399 1133 252433
rect 1167 252399 1225 252433
rect 1259 252399 1317 252433
rect 1121 252181 1340 252399
rect 1121 252039 1225 252147
rect 1259 252073 1340 252181
rect 1121 251889 1340 252039
rect 1104 251855 1133 251889
rect 1167 251855 1225 251889
rect 1259 251855 1317 251889
rect 1121 251705 1340 251855
rect 1121 251597 1225 251705
rect 1259 251563 1340 251671
rect 1121 251345 1340 251563
rect 1104 251311 1133 251345
rect 1167 251311 1225 251345
rect 1259 251311 1317 251345
rect 1121 251093 1340 251311
rect 1121 250951 1225 251059
rect 1259 250985 1340 251093
rect 1121 250801 1340 250951
rect 1104 250767 1133 250801
rect 1167 250767 1225 250801
rect 1259 250767 1317 250801
rect 1121 250617 1340 250767
rect 1121 250509 1225 250617
rect 1259 250475 1340 250583
rect 1121 250257 1340 250475
rect 1104 250223 1133 250257
rect 1167 250223 1225 250257
rect 1259 250223 1317 250257
rect 1121 250005 1340 250223
rect 1121 249863 1225 249971
rect 1259 249897 1340 250005
rect 1121 249713 1340 249863
rect 1104 249679 1133 249713
rect 1167 249679 1225 249713
rect 1259 249679 1317 249713
rect 1121 249529 1340 249679
rect 1121 249421 1225 249529
rect 1259 249387 1340 249495
rect 1121 249169 1340 249387
rect 1104 249135 1133 249169
rect 1167 249135 1225 249169
rect 1259 249135 1317 249169
rect 1121 248917 1340 249135
rect 1121 248775 1225 248883
rect 1259 248809 1340 248917
rect 1121 248625 1340 248775
rect 1104 248591 1133 248625
rect 1167 248591 1225 248625
rect 1259 248591 1317 248625
rect 1121 248441 1340 248591
rect 1121 248333 1225 248441
rect 1259 248299 1340 248407
rect 1121 248081 1340 248299
rect 1104 248047 1133 248081
rect 1167 248047 1225 248081
rect 1259 248047 1317 248081
rect 1121 247829 1340 248047
rect 1121 247687 1225 247795
rect 1259 247721 1340 247829
rect 1121 247537 1340 247687
rect 1104 247503 1133 247537
rect 1167 247503 1225 247537
rect 1259 247503 1317 247537
rect 1121 247353 1340 247503
rect 1121 247245 1225 247353
rect 1259 247211 1340 247319
rect 1121 246993 1340 247211
rect 1104 246959 1133 246993
rect 1167 246959 1225 246993
rect 1259 246959 1317 246993
rect 1121 246741 1340 246959
rect 1121 246599 1225 246707
rect 1259 246633 1340 246741
rect 1121 246449 1340 246599
rect 1104 246415 1133 246449
rect 1167 246415 1225 246449
rect 1259 246415 1317 246449
rect 1121 246265 1340 246415
rect 1121 246157 1225 246265
rect 1259 246123 1340 246231
rect 1121 245905 1340 246123
rect 1104 245871 1133 245905
rect 1167 245871 1225 245905
rect 1259 245871 1317 245905
rect 1121 245653 1340 245871
rect 1121 245511 1225 245619
rect 1259 245545 1340 245653
rect 1121 245361 1340 245511
rect 1104 245327 1133 245361
rect 1167 245327 1225 245361
rect 1259 245327 1317 245361
rect 1121 245177 1340 245327
rect 1121 245069 1225 245177
rect 1259 245035 1340 245143
rect 1121 244817 1340 245035
rect 1104 244783 1133 244817
rect 1167 244783 1225 244817
rect 1259 244783 1317 244817
rect 1121 244565 1340 244783
rect 1121 244423 1225 244531
rect 1259 244457 1340 244565
rect 1121 244273 1340 244423
rect 1104 244239 1133 244273
rect 1167 244239 1225 244273
rect 1259 244239 1317 244273
rect 1121 244089 1340 244239
rect 1121 243981 1225 244089
rect 1259 243947 1340 244055
rect 1121 243729 1340 243947
rect 1104 243695 1133 243729
rect 1167 243695 1225 243729
rect 1259 243695 1317 243729
rect 1121 243477 1340 243695
rect 1121 243335 1225 243443
rect 1259 243369 1340 243477
rect 1121 243185 1340 243335
rect 1104 243151 1133 243185
rect 1167 243151 1225 243185
rect 1259 243151 1317 243185
rect 1121 243001 1340 243151
rect 1121 242893 1225 243001
rect 1259 242859 1340 242967
rect 1121 242641 1340 242859
rect 1104 242607 1133 242641
rect 1167 242607 1225 242641
rect 1259 242607 1317 242641
rect 1121 242389 1340 242607
rect 1121 242247 1225 242355
rect 1259 242281 1340 242389
rect 1121 242097 1340 242247
rect 1104 242063 1133 242097
rect 1167 242063 1225 242097
rect 1259 242063 1317 242097
rect 1121 241913 1340 242063
rect 1121 241805 1225 241913
rect 1259 241771 1340 241879
rect 1121 241553 1340 241771
rect 1104 241519 1133 241553
rect 1167 241519 1225 241553
rect 1259 241519 1317 241553
rect 1121 241301 1340 241519
rect 1121 241159 1225 241267
rect 1259 241193 1340 241301
rect 1121 241009 1340 241159
rect 1104 240975 1133 241009
rect 1167 240975 1225 241009
rect 1259 240975 1317 241009
rect 1121 240825 1340 240975
rect 1121 240717 1225 240825
rect 1259 240683 1340 240791
rect 1121 240465 1340 240683
rect 1104 240431 1133 240465
rect 1167 240431 1225 240465
rect 1259 240431 1317 240465
rect 1121 240213 1340 240431
rect 1121 240071 1225 240179
rect 1259 240105 1340 240213
rect 1121 239921 1340 240071
rect 1104 239887 1133 239921
rect 1167 239887 1225 239921
rect 1259 239887 1317 239921
rect 1121 239737 1340 239887
rect 1121 239629 1225 239737
rect 1259 239595 1340 239703
rect 1121 239377 1340 239595
rect 1104 239343 1133 239377
rect 1167 239343 1225 239377
rect 1259 239343 1317 239377
rect 1121 239125 1340 239343
rect 1121 238983 1225 239091
rect 1259 239017 1340 239125
rect 1121 238833 1340 238983
rect 1104 238799 1133 238833
rect 1167 238799 1225 238833
rect 1259 238799 1317 238833
rect 1121 238649 1340 238799
rect 1121 238541 1225 238649
rect 1259 238507 1340 238615
rect 1121 238289 1340 238507
rect 1104 238255 1133 238289
rect 1167 238255 1225 238289
rect 1259 238255 1317 238289
rect 1121 238037 1340 238255
rect 1121 237895 1225 238003
rect 1259 237929 1340 238037
rect 1121 237745 1340 237895
rect 1104 237711 1133 237745
rect 1167 237711 1225 237745
rect 1259 237711 1317 237745
rect 1121 237561 1340 237711
rect 1121 237453 1225 237561
rect 1259 237419 1340 237527
rect 1121 237201 1340 237419
rect 1104 237167 1133 237201
rect 1167 237167 1225 237201
rect 1259 237167 1317 237201
rect 1121 236949 1340 237167
rect 1121 236807 1225 236915
rect 1259 236841 1340 236949
rect 1121 236657 1340 236807
rect 1104 236623 1133 236657
rect 1167 236623 1225 236657
rect 1259 236623 1317 236657
rect 1121 236473 1340 236623
rect 1121 236365 1225 236473
rect 1259 236331 1340 236439
rect 1121 236113 1340 236331
rect 1104 236079 1133 236113
rect 1167 236079 1225 236113
rect 1259 236079 1317 236113
rect 1121 235861 1340 236079
rect 1121 235719 1225 235827
rect 1259 235753 1340 235861
rect 1121 235569 1340 235719
rect 1104 235535 1133 235569
rect 1167 235535 1225 235569
rect 1259 235535 1317 235569
rect 1121 235385 1340 235535
rect 1121 235277 1225 235385
rect 1259 235243 1340 235351
rect 1121 235025 1340 235243
rect 1104 234991 1133 235025
rect 1167 234991 1225 235025
rect 1259 234991 1317 235025
rect 1121 234773 1340 234991
rect 1121 234631 1225 234739
rect 1259 234665 1340 234773
rect 1121 234481 1340 234631
rect 1104 234447 1133 234481
rect 1167 234447 1225 234481
rect 1259 234447 1317 234481
rect 1121 234297 1340 234447
rect 1121 234189 1225 234297
rect 1259 234155 1340 234263
rect 1121 233937 1340 234155
rect 1104 233903 1133 233937
rect 1167 233903 1225 233937
rect 1259 233903 1317 233937
rect 1121 233685 1340 233903
rect 1121 233543 1225 233651
rect 1259 233577 1340 233685
rect 1121 233393 1340 233543
rect 1104 233359 1133 233393
rect 1167 233359 1225 233393
rect 1259 233359 1317 233393
rect 1121 233209 1340 233359
rect 1121 233101 1225 233209
rect 1259 233067 1340 233175
rect 1121 232849 1340 233067
rect 1104 232815 1133 232849
rect 1167 232815 1225 232849
rect 1259 232815 1317 232849
rect 1121 232597 1340 232815
rect 1121 232455 1225 232563
rect 1259 232489 1340 232597
rect 1121 232305 1340 232455
rect 1104 232271 1133 232305
rect 1167 232271 1225 232305
rect 1259 232271 1317 232305
rect 1121 232121 1340 232271
rect 1121 232013 1225 232121
rect 1259 231979 1340 232087
rect 1121 231761 1340 231979
rect 1104 231727 1133 231761
rect 1167 231727 1225 231761
rect 1259 231727 1317 231761
rect 1121 231509 1340 231727
rect 1121 231367 1225 231475
rect 1259 231401 1340 231509
rect 1121 231217 1340 231367
rect 1104 231183 1133 231217
rect 1167 231183 1225 231217
rect 1259 231183 1317 231217
rect 1121 231033 1340 231183
rect 1121 230925 1225 231033
rect 1259 230891 1340 230999
rect 1121 230673 1340 230891
rect 1104 230639 1133 230673
rect 1167 230639 1225 230673
rect 1259 230639 1317 230673
rect 1121 230421 1340 230639
rect 1121 230279 1225 230387
rect 1259 230313 1340 230421
rect 1121 230129 1340 230279
rect 1104 230095 1133 230129
rect 1167 230095 1225 230129
rect 1259 230095 1317 230129
rect 1121 229945 1340 230095
rect 1121 229837 1225 229945
rect 1259 229803 1340 229911
rect 1121 229585 1340 229803
rect 1104 229551 1133 229585
rect 1167 229551 1225 229585
rect 1259 229551 1317 229585
rect 1121 229333 1340 229551
rect 1121 229191 1225 229299
rect 1259 229225 1340 229333
rect 1121 229041 1340 229191
rect 1104 229007 1133 229041
rect 1167 229007 1225 229041
rect 1259 229007 1317 229041
rect 1121 228857 1340 229007
rect 1121 228749 1225 228857
rect 1259 228715 1340 228823
rect 1121 228497 1340 228715
rect 1104 228463 1133 228497
rect 1167 228463 1225 228497
rect 1259 228463 1317 228497
rect 1121 228245 1340 228463
rect 1121 228103 1225 228211
rect 1259 228137 1340 228245
rect 1121 227953 1340 228103
rect 1104 227919 1133 227953
rect 1167 227919 1225 227953
rect 1259 227919 1317 227953
rect 1121 227769 1340 227919
rect 1121 227661 1225 227769
rect 1259 227627 1340 227735
rect 1121 227409 1340 227627
rect 1104 227375 1133 227409
rect 1167 227375 1225 227409
rect 1259 227375 1317 227409
rect 1121 227157 1340 227375
rect 1121 227015 1225 227123
rect 1259 227049 1340 227157
rect 1121 226865 1340 227015
rect 1104 226831 1133 226865
rect 1167 226831 1225 226865
rect 1259 226831 1317 226865
rect 1121 226681 1340 226831
rect 1121 226573 1225 226681
rect 1259 226539 1340 226647
rect 1121 226321 1340 226539
rect 1104 226287 1133 226321
rect 1167 226287 1225 226321
rect 1259 226287 1317 226321
rect 1121 226069 1340 226287
rect 1121 225927 1225 226035
rect 1259 225961 1340 226069
rect 1121 225777 1340 225927
rect 1104 225743 1133 225777
rect 1167 225743 1225 225777
rect 1259 225743 1317 225777
rect 1121 225593 1340 225743
rect 1121 225485 1225 225593
rect 1259 225451 1340 225559
rect 1121 225233 1340 225451
rect 1104 225199 1133 225233
rect 1167 225199 1225 225233
rect 1259 225199 1317 225233
rect 1121 224981 1340 225199
rect 1121 224839 1225 224947
rect 1259 224873 1340 224981
rect 1121 224689 1340 224839
rect 1104 224655 1133 224689
rect 1167 224655 1225 224689
rect 1259 224655 1317 224689
rect 1121 224505 1340 224655
rect 1121 224397 1225 224505
rect 1259 224363 1340 224471
rect 1121 224145 1340 224363
rect 1104 224111 1133 224145
rect 1167 224111 1225 224145
rect 1259 224111 1317 224145
rect 1121 223893 1340 224111
rect 1121 223751 1225 223859
rect 1259 223785 1340 223893
rect 1121 223601 1340 223751
rect 1104 223567 1133 223601
rect 1167 223567 1225 223601
rect 1259 223567 1317 223601
rect 1121 223417 1340 223567
rect 1121 223309 1225 223417
rect 1259 223275 1340 223383
rect 1121 223057 1340 223275
rect 1104 223023 1133 223057
rect 1167 223023 1225 223057
rect 1259 223023 1317 223057
rect 1121 222805 1340 223023
rect 1121 222663 1225 222771
rect 1259 222697 1340 222805
rect 1121 222513 1340 222663
rect 1104 222479 1133 222513
rect 1167 222479 1225 222513
rect 1259 222479 1317 222513
rect 1121 222329 1340 222479
rect 1121 222221 1225 222329
rect 1259 222187 1340 222295
rect 1121 221969 1340 222187
rect 1104 221935 1133 221969
rect 1167 221935 1225 221969
rect 1259 221935 1317 221969
rect 1121 221717 1340 221935
rect 1121 221575 1225 221683
rect 1259 221609 1340 221717
rect 1121 221425 1340 221575
rect 1104 221391 1133 221425
rect 1167 221391 1225 221425
rect 1259 221391 1317 221425
rect 1121 221241 1340 221391
rect 1121 221133 1225 221241
rect 1259 221099 1340 221207
rect 1121 220881 1340 221099
rect 1104 220847 1133 220881
rect 1167 220847 1225 220881
rect 1259 220847 1317 220881
rect 1121 220629 1340 220847
rect 1121 220487 1225 220595
rect 1259 220521 1340 220629
rect 1121 220337 1340 220487
rect 1104 220303 1133 220337
rect 1167 220303 1225 220337
rect 1259 220303 1317 220337
rect 1121 220153 1340 220303
rect 1121 220045 1225 220153
rect 1259 220011 1340 220119
rect 1121 219793 1340 220011
rect 1104 219759 1133 219793
rect 1167 219759 1225 219793
rect 1259 219759 1317 219793
rect 1121 219541 1340 219759
rect 1121 219399 1225 219507
rect 1259 219433 1340 219541
rect 1121 219249 1340 219399
rect 1104 219215 1133 219249
rect 1167 219215 1225 219249
rect 1259 219215 1317 219249
rect 1121 219065 1340 219215
rect 1121 218957 1225 219065
rect 1259 218923 1340 219031
rect 1121 218705 1340 218923
rect 1104 218671 1133 218705
rect 1167 218671 1225 218705
rect 1259 218671 1317 218705
rect 1121 218453 1340 218671
rect 1121 218311 1225 218419
rect 1259 218345 1340 218453
rect 1121 218161 1340 218311
rect 1104 218127 1133 218161
rect 1167 218127 1225 218161
rect 1259 218127 1317 218161
rect 1121 217977 1340 218127
rect 1121 217869 1225 217977
rect 1259 217835 1340 217943
rect 1121 217617 1340 217835
rect 1104 217583 1133 217617
rect 1167 217583 1225 217617
rect 1259 217583 1317 217617
rect 1121 217365 1340 217583
rect 1121 217223 1225 217331
rect 1259 217257 1340 217365
rect 1121 217073 1340 217223
rect 1104 217039 1133 217073
rect 1167 217039 1225 217073
rect 1259 217039 1317 217073
rect 1121 216889 1340 217039
rect 1121 216781 1225 216889
rect 1259 216747 1340 216855
rect 1121 216529 1340 216747
rect 1104 216495 1133 216529
rect 1167 216495 1225 216529
rect 1259 216495 1317 216529
rect 1121 216277 1340 216495
rect 1121 216135 1225 216243
rect 1259 216169 1340 216277
rect 1121 215985 1340 216135
rect 1104 215951 1133 215985
rect 1167 215951 1225 215985
rect 1259 215951 1317 215985
rect 1121 215801 1340 215951
rect 1121 215693 1225 215801
rect 1259 215659 1340 215767
rect 1121 215441 1340 215659
rect 1104 215407 1133 215441
rect 1167 215407 1225 215441
rect 1259 215407 1317 215441
rect 1121 215189 1340 215407
rect 1121 215047 1225 215155
rect 1259 215081 1340 215189
rect 1121 214897 1340 215047
rect 1104 214863 1133 214897
rect 1167 214863 1225 214897
rect 1259 214863 1317 214897
rect 1121 214713 1340 214863
rect 1121 214605 1225 214713
rect 1259 214571 1340 214679
rect 1121 214353 1340 214571
rect 1104 214319 1133 214353
rect 1167 214319 1225 214353
rect 1259 214319 1317 214353
rect 1121 214101 1340 214319
rect 1121 213959 1225 214067
rect 1259 213993 1340 214101
rect 1121 213809 1340 213959
rect 1104 213775 1133 213809
rect 1167 213775 1225 213809
rect 1259 213775 1317 213809
rect 1121 213625 1340 213775
rect 1121 213517 1225 213625
rect 1259 213483 1340 213591
rect 1121 213265 1340 213483
rect 1104 213231 1133 213265
rect 1167 213231 1225 213265
rect 1259 213231 1317 213265
rect 1121 213013 1340 213231
rect 1121 212871 1225 212979
rect 1259 212905 1340 213013
rect 1121 212721 1340 212871
rect 1104 212687 1133 212721
rect 1167 212687 1225 212721
rect 1259 212687 1317 212721
rect 1121 212537 1340 212687
rect 1121 212429 1225 212537
rect 1259 212395 1340 212503
rect 1121 212177 1340 212395
rect 1104 212143 1133 212177
rect 1167 212143 1225 212177
rect 1259 212143 1317 212177
rect 1121 211925 1340 212143
rect 1121 211783 1225 211891
rect 1259 211817 1340 211925
rect 1121 211633 1340 211783
rect 1104 211599 1133 211633
rect 1167 211599 1225 211633
rect 1259 211599 1317 211633
rect 1121 211449 1340 211599
rect 1121 211341 1225 211449
rect 1259 211307 1340 211415
rect 1121 211089 1340 211307
rect 1104 211055 1133 211089
rect 1167 211055 1225 211089
rect 1259 211055 1317 211089
rect 1121 210837 1340 211055
rect 1121 210695 1225 210803
rect 1259 210729 1340 210837
rect 1121 210545 1340 210695
rect 1104 210511 1133 210545
rect 1167 210511 1225 210545
rect 1259 210511 1317 210545
rect 1121 210361 1340 210511
rect 1121 210253 1225 210361
rect 1259 210219 1340 210327
rect 1121 210001 1340 210219
rect 1104 209967 1133 210001
rect 1167 209967 1225 210001
rect 1259 209967 1317 210001
rect 1121 209749 1340 209967
rect 1121 209607 1225 209715
rect 1259 209641 1340 209749
rect 1121 209457 1340 209607
rect 1104 209423 1133 209457
rect 1167 209423 1225 209457
rect 1259 209423 1317 209457
rect 1121 209273 1340 209423
rect 1121 209165 1225 209273
rect 1259 209131 1340 209239
rect 1121 208913 1340 209131
rect 1104 208879 1133 208913
rect 1167 208879 1225 208913
rect 1259 208879 1317 208913
rect 1121 208661 1340 208879
rect 1121 208519 1225 208627
rect 1259 208553 1340 208661
rect 1121 208369 1340 208519
rect 1104 208335 1133 208369
rect 1167 208335 1225 208369
rect 1259 208335 1317 208369
rect 1121 208185 1340 208335
rect 1121 208077 1225 208185
rect 1259 208043 1340 208151
rect 1121 207825 1340 208043
rect 1104 207791 1133 207825
rect 1167 207791 1225 207825
rect 1259 207791 1317 207825
rect 1121 207573 1340 207791
rect 1121 207431 1225 207539
rect 1259 207465 1340 207573
rect 1121 207281 1340 207431
rect 1104 207247 1133 207281
rect 1167 207247 1225 207281
rect 1259 207247 1317 207281
rect 1121 207097 1340 207247
rect 1121 206989 1225 207097
rect 1259 206955 1340 207063
rect 1121 206737 1340 206955
rect 1104 206703 1133 206737
rect 1167 206703 1225 206737
rect 1259 206703 1317 206737
rect 1121 206485 1340 206703
rect 1121 206343 1225 206451
rect 1259 206377 1340 206485
rect 1121 206193 1340 206343
rect 1104 206159 1133 206193
rect 1167 206159 1225 206193
rect 1259 206159 1317 206193
rect 1121 206009 1340 206159
rect 1121 205901 1225 206009
rect 1259 205867 1340 205975
rect 1121 205649 1340 205867
rect 1104 205615 1133 205649
rect 1167 205615 1225 205649
rect 1259 205615 1317 205649
rect 1121 205397 1340 205615
rect 1121 205255 1225 205363
rect 1259 205289 1340 205397
rect 1121 205105 1340 205255
rect 1104 205071 1133 205105
rect 1167 205071 1225 205105
rect 1259 205071 1317 205105
rect 1121 204921 1340 205071
rect 1121 204813 1225 204921
rect 1259 204779 1340 204887
rect 1121 204561 1340 204779
rect 1104 204527 1133 204561
rect 1167 204527 1225 204561
rect 1259 204527 1317 204561
rect 1121 204309 1340 204527
rect 1121 204167 1225 204275
rect 1259 204201 1340 204309
rect 1121 204017 1340 204167
rect 1104 203983 1133 204017
rect 1167 203983 1225 204017
rect 1259 203983 1317 204017
rect 1121 203833 1340 203983
rect 1121 203725 1225 203833
rect 1259 203691 1340 203799
rect 1121 203473 1340 203691
rect 1104 203439 1133 203473
rect 1167 203439 1225 203473
rect 1259 203439 1317 203473
rect 1121 203221 1340 203439
rect 1121 203079 1225 203187
rect 1259 203113 1340 203221
rect 1121 202929 1340 203079
rect 1104 202895 1133 202929
rect 1167 202895 1225 202929
rect 1259 202895 1317 202929
rect 1121 202745 1340 202895
rect 1121 202637 1225 202745
rect 1259 202603 1340 202711
rect 1121 202385 1340 202603
rect 1104 202351 1133 202385
rect 1167 202351 1225 202385
rect 1259 202351 1317 202385
rect 1121 202133 1340 202351
rect 1121 201991 1225 202099
rect 1259 202025 1340 202133
rect 1121 201841 1340 201991
rect 1104 201807 1133 201841
rect 1167 201807 1225 201841
rect 1259 201807 1317 201841
rect 1121 201657 1340 201807
rect 1121 201549 1225 201657
rect 1259 201515 1340 201623
rect 1121 201297 1340 201515
rect 1104 201263 1133 201297
rect 1167 201263 1225 201297
rect 1259 201263 1317 201297
rect 1121 201045 1340 201263
rect 1121 200903 1225 201011
rect 1259 200937 1340 201045
rect 1121 200753 1340 200903
rect 1104 200719 1133 200753
rect 1167 200719 1225 200753
rect 1259 200719 1317 200753
rect 1121 200569 1340 200719
rect 1121 200461 1225 200569
rect 1259 200427 1340 200535
rect 1121 200209 1340 200427
rect 1104 200175 1133 200209
rect 1167 200175 1225 200209
rect 1259 200175 1317 200209
rect 1121 199957 1340 200175
rect 1121 199815 1225 199923
rect 1259 199849 1340 199957
rect 1121 199665 1340 199815
rect 1104 199631 1133 199665
rect 1167 199631 1225 199665
rect 1259 199631 1317 199665
rect 1121 199481 1340 199631
rect 1121 199373 1225 199481
rect 1259 199339 1340 199447
rect 1121 199121 1340 199339
rect 1104 199087 1133 199121
rect 1167 199087 1225 199121
rect 1259 199087 1317 199121
rect 1121 198869 1340 199087
rect 1121 198727 1225 198835
rect 1259 198761 1340 198869
rect 1121 198577 1340 198727
rect 1104 198543 1133 198577
rect 1167 198543 1225 198577
rect 1259 198543 1317 198577
rect 1121 198393 1340 198543
rect 1121 198285 1225 198393
rect 1259 198251 1340 198359
rect 1121 198033 1340 198251
rect 1104 197999 1133 198033
rect 1167 197999 1225 198033
rect 1259 197999 1317 198033
rect 1121 197781 1340 197999
rect 1121 197639 1225 197747
rect 1259 197673 1340 197781
rect 1121 197489 1340 197639
rect 1104 197455 1133 197489
rect 1167 197455 1225 197489
rect 1259 197455 1317 197489
rect 1121 197305 1340 197455
rect 1121 197197 1225 197305
rect 1259 197163 1340 197271
rect 1121 196945 1340 197163
rect 1104 196911 1133 196945
rect 1167 196911 1225 196945
rect 1259 196911 1317 196945
rect 1121 196693 1340 196911
rect 1121 196551 1225 196659
rect 1259 196585 1340 196693
rect 1121 196401 1340 196551
rect 1104 196367 1133 196401
rect 1167 196367 1225 196401
rect 1259 196367 1317 196401
rect 1121 196217 1340 196367
rect 1121 196109 1225 196217
rect 1259 196075 1340 196183
rect 1121 195857 1340 196075
rect 1104 195823 1133 195857
rect 1167 195823 1225 195857
rect 1259 195823 1317 195857
rect 1121 195605 1340 195823
rect 1121 195463 1225 195571
rect 1259 195497 1340 195605
rect 1121 195313 1340 195463
rect 1104 195279 1133 195313
rect 1167 195279 1225 195313
rect 1259 195279 1317 195313
rect 1121 195129 1340 195279
rect 1121 195021 1225 195129
rect 1259 194987 1340 195095
rect 1121 194769 1340 194987
rect 1104 194735 1133 194769
rect 1167 194735 1225 194769
rect 1259 194735 1317 194769
rect 1121 194517 1340 194735
rect 1121 194375 1225 194483
rect 1259 194409 1340 194517
rect 1121 194225 1340 194375
rect 1104 194191 1133 194225
rect 1167 194191 1225 194225
rect 1259 194191 1317 194225
rect 1121 194041 1340 194191
rect 1121 193933 1225 194041
rect 1259 193899 1340 194007
rect 1121 193681 1340 193899
rect 1104 193647 1133 193681
rect 1167 193647 1225 193681
rect 1259 193647 1317 193681
rect 1121 193429 1340 193647
rect 1121 193287 1225 193395
rect 1259 193321 1340 193429
rect 1121 193137 1340 193287
rect 1104 193103 1133 193137
rect 1167 193103 1225 193137
rect 1259 193103 1317 193137
rect 1121 192953 1340 193103
rect 1121 192845 1225 192953
rect 1259 192811 1340 192919
rect 1121 192593 1340 192811
rect 1104 192559 1133 192593
rect 1167 192559 1225 192593
rect 1259 192559 1317 192593
rect 1121 192341 1340 192559
rect 1121 192199 1225 192307
rect 1259 192233 1340 192341
rect 1121 192049 1340 192199
rect 1104 192015 1133 192049
rect 1167 192015 1225 192049
rect 1259 192015 1317 192049
rect 1121 191865 1340 192015
rect 1121 191757 1225 191865
rect 1259 191723 1340 191831
rect 1121 191505 1340 191723
rect 1104 191471 1133 191505
rect 1167 191471 1225 191505
rect 1259 191471 1317 191505
rect 1121 191253 1340 191471
rect 1121 191111 1225 191219
rect 1259 191145 1340 191253
rect 1121 190961 1340 191111
rect 1104 190927 1133 190961
rect 1167 190927 1225 190961
rect 1259 190927 1317 190961
rect 1121 190777 1340 190927
rect 1121 190669 1225 190777
rect 1259 190635 1340 190743
rect 1121 190417 1340 190635
rect 1104 190383 1133 190417
rect 1167 190383 1225 190417
rect 1259 190383 1317 190417
rect 1121 190165 1340 190383
rect 1121 190023 1225 190131
rect 1259 190057 1340 190165
rect 1121 189873 1340 190023
rect 1104 189839 1133 189873
rect 1167 189839 1225 189873
rect 1259 189839 1317 189873
rect 1121 189689 1340 189839
rect 1121 189581 1225 189689
rect 1259 189547 1340 189655
rect 1121 189329 1340 189547
rect 1104 189295 1133 189329
rect 1167 189295 1225 189329
rect 1259 189295 1317 189329
rect 1121 189077 1340 189295
rect 1121 188935 1225 189043
rect 1259 188969 1340 189077
rect 1121 188785 1340 188935
rect 1104 188751 1133 188785
rect 1167 188751 1225 188785
rect 1259 188751 1317 188785
rect 1121 188601 1340 188751
rect 1121 188493 1225 188601
rect 1259 188459 1340 188567
rect 1121 188241 1340 188459
rect 1104 188207 1133 188241
rect 1167 188207 1225 188241
rect 1259 188207 1317 188241
rect 1121 187989 1340 188207
rect 1121 187847 1225 187955
rect 1259 187881 1340 187989
rect 1121 187697 1340 187847
rect 1104 187663 1133 187697
rect 1167 187663 1225 187697
rect 1259 187663 1317 187697
rect 1121 187513 1340 187663
rect 1121 187405 1225 187513
rect 1259 187371 1340 187479
rect 1121 187153 1340 187371
rect 1104 187119 1133 187153
rect 1167 187119 1225 187153
rect 1259 187119 1317 187153
rect 1121 186901 1340 187119
rect 1121 186759 1225 186867
rect 1259 186793 1340 186901
rect 1121 186609 1340 186759
rect 1104 186575 1133 186609
rect 1167 186575 1225 186609
rect 1259 186575 1317 186609
rect 1121 186425 1340 186575
rect 1121 186317 1225 186425
rect 1259 186283 1340 186391
rect 1121 186065 1340 186283
rect 1104 186031 1133 186065
rect 1167 186031 1225 186065
rect 1259 186031 1317 186065
rect 1121 185813 1340 186031
rect 1121 185671 1225 185779
rect 1259 185705 1340 185813
rect 1121 185521 1340 185671
rect 1104 185487 1133 185521
rect 1167 185487 1225 185521
rect 1259 185487 1317 185521
rect 1121 185337 1340 185487
rect 1121 185229 1225 185337
rect 1259 185195 1340 185303
rect 1121 184977 1340 185195
rect 1104 184943 1133 184977
rect 1167 184943 1225 184977
rect 1259 184943 1317 184977
rect 1121 184725 1340 184943
rect 1121 184583 1225 184691
rect 1259 184617 1340 184725
rect 1121 184433 1340 184583
rect 1104 184399 1133 184433
rect 1167 184399 1225 184433
rect 1259 184399 1317 184433
rect 1121 184249 1340 184399
rect 1121 184141 1225 184249
rect 1259 184107 1340 184215
rect 1121 183889 1340 184107
rect 1104 183855 1133 183889
rect 1167 183855 1225 183889
rect 1259 183855 1317 183889
rect 1121 183637 1340 183855
rect 1121 183495 1225 183603
rect 1259 183529 1340 183637
rect 1121 183345 1340 183495
rect 1104 183311 1133 183345
rect 1167 183311 1225 183345
rect 1259 183311 1317 183345
rect 1121 183161 1340 183311
rect 1121 183053 1225 183161
rect 1259 183019 1340 183127
rect 1121 182801 1340 183019
rect 1104 182767 1133 182801
rect 1167 182767 1225 182801
rect 1259 182767 1317 182801
rect 1121 182549 1340 182767
rect 1121 182407 1225 182515
rect 1259 182441 1340 182549
rect 1121 182257 1340 182407
rect 1104 182223 1133 182257
rect 1167 182223 1225 182257
rect 1259 182223 1317 182257
rect 1121 182073 1340 182223
rect 1121 181965 1225 182073
rect 1259 181931 1340 182039
rect 1121 181713 1340 181931
rect 1104 181679 1133 181713
rect 1167 181679 1225 181713
rect 1259 181679 1317 181713
rect 1121 181461 1340 181679
rect 1121 181319 1225 181427
rect 1259 181353 1340 181461
rect 1121 181169 1340 181319
rect 1104 181135 1133 181169
rect 1167 181135 1225 181169
rect 1259 181135 1317 181169
rect 1121 180985 1340 181135
rect 1121 180877 1225 180985
rect 1259 180843 1340 180951
rect 1121 180625 1340 180843
rect 1104 180591 1133 180625
rect 1167 180591 1225 180625
rect 1259 180591 1317 180625
rect 1121 180373 1340 180591
rect 1121 180231 1225 180339
rect 1259 180265 1340 180373
rect 1121 180081 1340 180231
rect 1104 180047 1133 180081
rect 1167 180047 1225 180081
rect 1259 180047 1317 180081
rect 1121 179897 1340 180047
rect 1121 179789 1225 179897
rect 1259 179755 1340 179863
rect 1121 179537 1340 179755
rect 1104 179503 1133 179537
rect 1167 179503 1225 179537
rect 1259 179503 1317 179537
rect 1121 179285 1340 179503
rect 1121 179143 1225 179251
rect 1259 179177 1340 179285
rect 1121 178993 1340 179143
rect 1104 178959 1133 178993
rect 1167 178959 1225 178993
rect 1259 178959 1317 178993
rect 1121 178809 1340 178959
rect 1121 178701 1225 178809
rect 1259 178667 1340 178775
rect 1121 178449 1340 178667
rect 1104 178415 1133 178449
rect 1167 178415 1225 178449
rect 1259 178415 1317 178449
rect 1121 178197 1340 178415
rect 1121 178055 1225 178163
rect 1259 178089 1340 178197
rect 1121 177905 1340 178055
rect 1104 177871 1133 177905
rect 1167 177871 1225 177905
rect 1259 177871 1317 177905
rect 1121 177721 1340 177871
rect 1121 177613 1225 177721
rect 1259 177579 1340 177687
rect 1121 177361 1340 177579
rect 1104 177327 1133 177361
rect 1167 177327 1225 177361
rect 1259 177327 1317 177361
rect 1121 177109 1340 177327
rect 1121 176967 1225 177075
rect 1259 177001 1340 177109
rect 1121 176817 1340 176967
rect 1104 176783 1133 176817
rect 1167 176783 1225 176817
rect 1259 176783 1317 176817
rect 1121 176633 1340 176783
rect 1121 176525 1225 176633
rect 1259 176491 1340 176599
rect 1121 176273 1340 176491
rect 1104 176239 1133 176273
rect 1167 176239 1225 176273
rect 1259 176239 1317 176273
rect 1121 176021 1340 176239
rect 1121 175879 1225 175987
rect 1259 175913 1340 176021
rect 1121 175729 1340 175879
rect 1104 175695 1133 175729
rect 1167 175695 1225 175729
rect 1259 175695 1317 175729
rect 1121 175545 1340 175695
rect 1121 175437 1225 175545
rect 1259 175403 1340 175511
rect 1121 175185 1340 175403
rect 1104 175151 1133 175185
rect 1167 175151 1225 175185
rect 1259 175151 1317 175185
rect 1121 174933 1340 175151
rect 1121 174791 1225 174899
rect 1259 174825 1340 174933
rect 1121 174641 1340 174791
rect 1104 174607 1133 174641
rect 1167 174607 1225 174641
rect 1259 174607 1317 174641
rect 1121 174457 1340 174607
rect 1121 174349 1225 174457
rect 1259 174315 1340 174423
rect 1121 174097 1340 174315
rect 1104 174063 1133 174097
rect 1167 174063 1225 174097
rect 1259 174063 1317 174097
rect 1121 173845 1340 174063
rect 1121 173703 1225 173811
rect 1259 173737 1340 173845
rect 1121 173553 1340 173703
rect 1104 173519 1133 173553
rect 1167 173519 1225 173553
rect 1259 173519 1317 173553
rect 1121 173369 1340 173519
rect 1121 173261 1225 173369
rect 1259 173227 1340 173335
rect 1121 173009 1340 173227
rect 1104 172975 1133 173009
rect 1167 172975 1225 173009
rect 1259 172975 1317 173009
rect 1121 172757 1340 172975
rect 1121 172615 1225 172723
rect 1259 172649 1340 172757
rect 1121 172465 1340 172615
rect 1104 172431 1133 172465
rect 1167 172431 1225 172465
rect 1259 172431 1317 172465
rect 1121 172281 1340 172431
rect 1121 172173 1225 172281
rect 1259 172139 1340 172247
rect 1121 171921 1340 172139
rect 1104 171887 1133 171921
rect 1167 171887 1225 171921
rect 1259 171887 1317 171921
rect 1121 171669 1340 171887
rect 1121 171527 1225 171635
rect 1259 171561 1340 171669
rect 1121 171377 1340 171527
rect 1104 171343 1133 171377
rect 1167 171343 1225 171377
rect 1259 171343 1317 171377
rect 1121 171193 1340 171343
rect 1121 171085 1225 171193
rect 1259 171051 1340 171159
rect 1121 170833 1340 171051
rect 1104 170799 1133 170833
rect 1167 170799 1225 170833
rect 1259 170799 1317 170833
rect 1121 170581 1340 170799
rect 1121 170439 1225 170547
rect 1259 170473 1340 170581
rect 1121 170289 1340 170439
rect 1104 170255 1133 170289
rect 1167 170255 1225 170289
rect 1259 170255 1317 170289
rect 1121 170105 1340 170255
rect 1121 169997 1225 170105
rect 1259 169963 1340 170071
rect 1121 169745 1340 169963
rect 1104 169711 1133 169745
rect 1167 169711 1225 169745
rect 1259 169711 1317 169745
rect 1121 169493 1340 169711
rect 1121 169351 1225 169459
rect 1259 169385 1340 169493
rect 1121 169201 1340 169351
rect 1104 169167 1133 169201
rect 1167 169167 1225 169201
rect 1259 169167 1317 169201
rect 1121 169017 1340 169167
rect 1121 168909 1225 169017
rect 1259 168875 1340 168983
rect 1121 168657 1340 168875
rect 1104 168623 1133 168657
rect 1167 168623 1225 168657
rect 1259 168623 1317 168657
rect 1121 168405 1340 168623
rect 1121 168263 1225 168371
rect 1259 168297 1340 168405
rect 1121 168113 1340 168263
rect 1104 168079 1133 168113
rect 1167 168079 1225 168113
rect 1259 168079 1317 168113
rect 1121 167929 1340 168079
rect 1121 167821 1225 167929
rect 1259 167787 1340 167895
rect 1121 167569 1340 167787
rect 1104 167535 1133 167569
rect 1167 167535 1225 167569
rect 1259 167535 1317 167569
rect 1121 167317 1340 167535
rect 1121 167175 1225 167283
rect 1259 167209 1340 167317
rect 1121 167025 1340 167175
rect 1104 166991 1133 167025
rect 1167 166991 1225 167025
rect 1259 166991 1317 167025
rect 1121 166841 1340 166991
rect 1121 166733 1225 166841
rect 1259 166699 1340 166807
rect 1121 166481 1340 166699
rect 1104 166447 1133 166481
rect 1167 166447 1225 166481
rect 1259 166447 1317 166481
rect 1121 166229 1340 166447
rect 1121 166087 1225 166195
rect 1259 166121 1340 166229
rect 1121 165937 1340 166087
rect 1104 165903 1133 165937
rect 1167 165903 1225 165937
rect 1259 165903 1317 165937
rect 1121 165753 1340 165903
rect 1121 165645 1225 165753
rect 1259 165611 1340 165719
rect 1121 165393 1340 165611
rect 1104 165359 1133 165393
rect 1167 165359 1225 165393
rect 1259 165359 1317 165393
rect 1121 165141 1340 165359
rect 1121 164999 1225 165107
rect 1259 165033 1340 165141
rect 1121 164849 1340 164999
rect 1104 164815 1133 164849
rect 1167 164815 1225 164849
rect 1259 164815 1317 164849
rect 1121 164665 1340 164815
rect 1121 164557 1225 164665
rect 1259 164523 1340 164631
rect 1121 164305 1340 164523
rect 1104 164271 1133 164305
rect 1167 164271 1225 164305
rect 1259 164271 1317 164305
rect 1121 164053 1340 164271
rect 1121 163911 1225 164019
rect 1259 163945 1340 164053
rect 1121 163761 1340 163911
rect 1104 163727 1133 163761
rect 1167 163727 1225 163761
rect 1259 163727 1317 163761
rect 1121 163577 1340 163727
rect 1121 163469 1225 163577
rect 1259 163435 1340 163543
rect 1121 163217 1340 163435
rect 1104 163183 1133 163217
rect 1167 163183 1225 163217
rect 1259 163183 1317 163217
rect 1121 162965 1340 163183
rect 1121 162823 1225 162931
rect 1259 162857 1340 162965
rect 1121 162673 1340 162823
rect 1104 162639 1133 162673
rect 1167 162639 1225 162673
rect 1259 162639 1317 162673
rect 1121 162489 1340 162639
rect 1121 162381 1225 162489
rect 1259 162347 1340 162455
rect 1121 162129 1340 162347
rect 1104 162095 1133 162129
rect 1167 162095 1225 162129
rect 1259 162095 1317 162129
rect 1121 161877 1340 162095
rect 1121 161735 1225 161843
rect 1259 161769 1340 161877
rect 1121 161585 1340 161735
rect 1104 161551 1133 161585
rect 1167 161551 1225 161585
rect 1259 161551 1317 161585
rect 1121 161401 1340 161551
rect 1121 161293 1225 161401
rect 1259 161259 1340 161367
rect 1121 161041 1340 161259
rect 1104 161007 1133 161041
rect 1167 161007 1225 161041
rect 1259 161007 1317 161041
rect 1121 160789 1340 161007
rect 1121 160647 1225 160755
rect 1259 160681 1340 160789
rect 1121 160497 1340 160647
rect 1104 160463 1133 160497
rect 1167 160463 1225 160497
rect 1259 160463 1317 160497
rect 1121 160313 1340 160463
rect 1121 160205 1225 160313
rect 1259 160171 1340 160279
rect 1121 159953 1340 160171
rect 1104 159919 1133 159953
rect 1167 159919 1225 159953
rect 1259 159919 1317 159953
rect 1121 159701 1340 159919
rect 1121 159559 1225 159667
rect 1259 159593 1340 159701
rect 1121 159409 1340 159559
rect 1104 159375 1133 159409
rect 1167 159375 1225 159409
rect 1259 159375 1317 159409
rect 1121 159225 1340 159375
rect 1121 159117 1225 159225
rect 1259 159083 1340 159191
rect 1121 158865 1340 159083
rect 1104 158831 1133 158865
rect 1167 158831 1225 158865
rect 1259 158831 1317 158865
rect 1121 158613 1340 158831
rect 1121 158471 1225 158579
rect 1259 158505 1340 158613
rect 1121 158321 1340 158471
rect 1104 158287 1133 158321
rect 1167 158287 1225 158321
rect 1259 158287 1317 158321
rect 1121 158137 1340 158287
rect 1121 158029 1225 158137
rect 1259 157995 1340 158103
rect 1121 157777 1340 157995
rect 1104 157743 1133 157777
rect 1167 157743 1225 157777
rect 1259 157743 1317 157777
rect 1121 157525 1340 157743
rect 1121 157383 1225 157491
rect 1259 157417 1340 157525
rect 1121 157233 1340 157383
rect 1104 157199 1133 157233
rect 1167 157199 1225 157233
rect 1259 157199 1317 157233
rect 1121 157049 1340 157199
rect 1121 156941 1225 157049
rect 1259 156907 1340 157015
rect 1121 156689 1340 156907
rect 1104 156655 1133 156689
rect 1167 156655 1225 156689
rect 1259 156655 1317 156689
rect 1121 156437 1340 156655
rect 1121 156295 1225 156403
rect 1259 156329 1340 156437
rect 1121 156145 1340 156295
rect 1104 156111 1133 156145
rect 1167 156111 1225 156145
rect 1259 156111 1317 156145
rect 1121 155961 1340 156111
rect 1121 155853 1225 155961
rect 1259 155819 1340 155927
rect 1121 155601 1340 155819
rect 1104 155567 1133 155601
rect 1167 155567 1225 155601
rect 1259 155567 1317 155601
rect 1121 155349 1340 155567
rect 1121 155207 1225 155315
rect 1259 155241 1340 155349
rect 1121 155057 1340 155207
rect 1104 155023 1133 155057
rect 1167 155023 1225 155057
rect 1259 155023 1317 155057
rect 1121 154873 1340 155023
rect 1121 154765 1225 154873
rect 1259 154731 1340 154839
rect 1121 154513 1340 154731
rect 1104 154479 1133 154513
rect 1167 154479 1225 154513
rect 1259 154479 1317 154513
rect 1121 154261 1340 154479
rect 1121 154119 1225 154227
rect 1259 154153 1340 154261
rect 1121 153969 1340 154119
rect 1104 153935 1133 153969
rect 1167 153935 1225 153969
rect 1259 153935 1317 153969
rect 1121 153785 1340 153935
rect 1121 153677 1225 153785
rect 1259 153643 1340 153751
rect 1121 153425 1340 153643
rect 1104 153391 1133 153425
rect 1167 153391 1225 153425
rect 1259 153391 1317 153425
rect 1121 153173 1340 153391
rect 1121 153031 1225 153139
rect 1259 153065 1340 153173
rect 1121 152881 1340 153031
rect 1104 152847 1133 152881
rect 1167 152847 1225 152881
rect 1259 152847 1317 152881
rect 1121 152697 1340 152847
rect 1121 152589 1225 152697
rect 1259 152555 1340 152663
rect 1121 152337 1340 152555
rect 1104 152303 1133 152337
rect 1167 152303 1225 152337
rect 1259 152303 1317 152337
rect 1121 152085 1340 152303
rect 1121 151943 1225 152051
rect 1259 151977 1340 152085
rect 1121 151793 1340 151943
rect 1104 151759 1133 151793
rect 1167 151759 1225 151793
rect 1259 151759 1317 151793
rect 1121 151609 1340 151759
rect 1121 151501 1225 151609
rect 1259 151467 1340 151575
rect 1121 151249 1340 151467
rect 1104 151215 1133 151249
rect 1167 151215 1225 151249
rect 1259 151215 1317 151249
rect 1121 150997 1340 151215
rect 1121 150855 1225 150963
rect 1259 150889 1340 150997
rect 1121 150705 1340 150855
rect 1104 150671 1133 150705
rect 1167 150671 1225 150705
rect 1259 150671 1317 150705
rect 1121 150521 1340 150671
rect 1121 150413 1225 150521
rect 1259 150379 1340 150487
rect 1121 150161 1340 150379
rect 1104 150127 1133 150161
rect 1167 150127 1225 150161
rect 1259 150127 1317 150161
rect 1121 149909 1340 150127
rect 1121 149767 1225 149875
rect 1259 149801 1340 149909
rect 1121 149617 1340 149767
rect 1104 149583 1133 149617
rect 1167 149583 1225 149617
rect 1259 149583 1317 149617
rect 1121 149433 1340 149583
rect 1121 149325 1225 149433
rect 1259 149291 1340 149399
rect 1121 149073 1340 149291
rect 1104 149039 1133 149073
rect 1167 149039 1225 149073
rect 1259 149039 1317 149073
rect 1121 148821 1340 149039
rect 1121 148679 1225 148787
rect 1259 148713 1340 148821
rect 1121 148529 1340 148679
rect 1104 148495 1133 148529
rect 1167 148495 1225 148529
rect 1259 148495 1317 148529
rect 1121 148345 1340 148495
rect 1121 148237 1225 148345
rect 1259 148203 1340 148311
rect 1121 147985 1340 148203
rect 1104 147951 1133 147985
rect 1167 147951 1225 147985
rect 1259 147951 1317 147985
rect 1121 147733 1340 147951
rect 1121 147591 1225 147699
rect 1259 147625 1340 147733
rect 1121 147441 1340 147591
rect 1104 147407 1133 147441
rect 1167 147407 1225 147441
rect 1259 147407 1317 147441
rect 1121 147257 1340 147407
rect 1121 147149 1225 147257
rect 1259 147115 1340 147223
rect 1121 146897 1340 147115
rect 1104 146863 1133 146897
rect 1167 146863 1225 146897
rect 1259 146863 1317 146897
rect 1121 146645 1340 146863
rect 1121 146503 1225 146611
rect 1259 146537 1340 146645
rect 1121 146353 1340 146503
rect 1104 146319 1133 146353
rect 1167 146319 1225 146353
rect 1259 146319 1317 146353
rect 1121 146169 1340 146319
rect 1121 146061 1225 146169
rect 1259 146027 1340 146135
rect 1121 145809 1340 146027
rect 1104 145775 1133 145809
rect 1167 145775 1225 145809
rect 1259 145775 1317 145809
rect 1121 145557 1340 145775
rect 1121 145415 1225 145523
rect 1259 145449 1340 145557
rect 1121 145265 1340 145415
rect 1104 145231 1133 145265
rect 1167 145231 1225 145265
rect 1259 145231 1317 145265
rect 1121 145081 1340 145231
rect 1121 144973 1225 145081
rect 1259 144939 1340 145047
rect 1121 144721 1340 144939
rect 1104 144687 1133 144721
rect 1167 144687 1225 144721
rect 1259 144687 1317 144721
rect 1121 144469 1340 144687
rect 1121 144327 1225 144435
rect 1259 144361 1340 144469
rect 1121 144177 1340 144327
rect 1104 144143 1133 144177
rect 1167 144143 1225 144177
rect 1259 144143 1317 144177
rect 1121 143993 1340 144143
rect 1121 143885 1225 143993
rect 1259 143851 1340 143959
rect 1121 143633 1340 143851
rect 1104 143599 1133 143633
rect 1167 143599 1225 143633
rect 1259 143599 1317 143633
rect 1121 143381 1340 143599
rect 1121 143239 1225 143347
rect 1259 143273 1340 143381
rect 1121 143089 1340 143239
rect 1104 143055 1133 143089
rect 1167 143055 1225 143089
rect 1259 143055 1317 143089
rect 1121 142905 1340 143055
rect 1121 142797 1225 142905
rect 1259 142763 1340 142871
rect 1121 142545 1340 142763
rect 1104 142511 1133 142545
rect 1167 142511 1225 142545
rect 1259 142511 1317 142545
rect 1121 142293 1340 142511
rect 1121 142151 1225 142259
rect 1259 142185 1340 142293
rect 1121 142001 1340 142151
rect 1104 141967 1133 142001
rect 1167 141967 1225 142001
rect 1259 141967 1317 142001
rect 1121 141817 1340 141967
rect 1121 141709 1225 141817
rect 1259 141675 1340 141783
rect 1121 141457 1340 141675
rect 1104 141423 1133 141457
rect 1167 141423 1225 141457
rect 1259 141423 1317 141457
rect 1121 141205 1340 141423
rect 1121 141063 1225 141171
rect 1259 141097 1340 141205
rect 1121 140913 1340 141063
rect 1104 140879 1133 140913
rect 1167 140879 1225 140913
rect 1259 140879 1317 140913
rect 1121 140729 1340 140879
rect 1121 140621 1225 140729
rect 1259 140587 1340 140695
rect 1121 140369 1340 140587
rect 1104 140335 1133 140369
rect 1167 140335 1225 140369
rect 1259 140335 1317 140369
rect 1121 140117 1340 140335
rect 1121 139975 1225 140083
rect 1259 140009 1340 140117
rect 1121 139825 1340 139975
rect 1104 139791 1133 139825
rect 1167 139791 1225 139825
rect 1259 139791 1317 139825
rect 1121 139641 1340 139791
rect 1121 139533 1225 139641
rect 1259 139499 1340 139607
rect 1121 139281 1340 139499
rect 1104 139247 1133 139281
rect 1167 139247 1225 139281
rect 1259 139247 1317 139281
rect 1121 139029 1340 139247
rect 1121 138887 1225 138995
rect 1259 138921 1340 139029
rect 1121 138737 1340 138887
rect 1104 138703 1133 138737
rect 1167 138703 1225 138737
rect 1259 138703 1317 138737
rect 1121 138553 1340 138703
rect 1121 138445 1225 138553
rect 1259 138411 1340 138519
rect 1121 138193 1340 138411
rect 1104 138159 1133 138193
rect 1167 138159 1225 138193
rect 1259 138159 1317 138193
rect 1121 137941 1340 138159
rect 1121 137799 1225 137907
rect 1259 137833 1340 137941
rect 1121 137649 1340 137799
rect 1104 137615 1133 137649
rect 1167 137615 1225 137649
rect 1259 137615 1317 137649
rect 1121 137465 1340 137615
rect 1121 137357 1225 137465
rect 1259 137323 1340 137431
rect 1121 137105 1340 137323
rect 1104 137071 1133 137105
rect 1167 137071 1225 137105
rect 1259 137071 1317 137105
rect 1121 136853 1340 137071
rect 1121 136711 1225 136819
rect 1259 136745 1340 136853
rect 1121 136561 1340 136711
rect 1104 136527 1133 136561
rect 1167 136527 1225 136561
rect 1259 136527 1317 136561
rect 1121 136377 1340 136527
rect 1121 136269 1225 136377
rect 1259 136235 1340 136343
rect 1121 136017 1340 136235
rect 1104 135983 1133 136017
rect 1167 135983 1225 136017
rect 1259 135983 1317 136017
rect 1121 135765 1340 135983
rect 1121 135623 1225 135731
rect 1259 135657 1340 135765
rect 1121 135473 1340 135623
rect 1104 135439 1133 135473
rect 1167 135439 1225 135473
rect 1259 135439 1317 135473
rect 1121 135289 1340 135439
rect 1121 135181 1225 135289
rect 1259 135147 1340 135255
rect 1121 134929 1340 135147
rect 1104 134895 1133 134929
rect 1167 134895 1225 134929
rect 1259 134895 1317 134929
rect 1121 134677 1340 134895
rect 1121 134535 1225 134643
rect 1259 134569 1340 134677
rect 1121 134385 1340 134535
rect 1104 134351 1133 134385
rect 1167 134351 1225 134385
rect 1259 134351 1317 134385
rect 1121 134201 1340 134351
rect 1121 134093 1225 134201
rect 1259 134059 1340 134167
rect 1121 133841 1340 134059
rect 1104 133807 1133 133841
rect 1167 133807 1225 133841
rect 1259 133807 1317 133841
rect 1121 133589 1340 133807
rect 1121 133447 1225 133555
rect 1259 133481 1340 133589
rect 1121 133297 1340 133447
rect 1104 133263 1133 133297
rect 1167 133263 1225 133297
rect 1259 133263 1317 133297
rect 1121 133113 1340 133263
rect 1121 133005 1225 133113
rect 1259 132971 1340 133079
rect 1121 132753 1340 132971
rect 1104 132719 1133 132753
rect 1167 132719 1225 132753
rect 1259 132719 1317 132753
rect 1121 132501 1340 132719
rect 1121 132359 1225 132467
rect 1259 132393 1340 132501
rect 1121 132209 1340 132359
rect 1104 132175 1133 132209
rect 1167 132175 1225 132209
rect 1259 132175 1317 132209
rect 1121 132025 1340 132175
rect 1121 131917 1225 132025
rect 1259 131883 1340 131991
rect 1121 131665 1340 131883
rect 1104 131631 1133 131665
rect 1167 131631 1225 131665
rect 1259 131631 1317 131665
rect 1121 131413 1340 131631
rect 1121 131271 1225 131379
rect 1259 131305 1340 131413
rect 1121 131121 1340 131271
rect 1104 131087 1133 131121
rect 1167 131087 1225 131121
rect 1259 131087 1317 131121
rect 1121 130937 1340 131087
rect 1121 130829 1225 130937
rect 1259 130795 1340 130903
rect 1121 130577 1340 130795
rect 1104 130543 1133 130577
rect 1167 130543 1225 130577
rect 1259 130543 1317 130577
rect 1121 130325 1340 130543
rect 1121 130183 1225 130291
rect 1259 130217 1340 130325
rect 1121 130033 1340 130183
rect 1104 129999 1133 130033
rect 1167 129999 1225 130033
rect 1259 129999 1317 130033
rect 1121 129849 1340 129999
rect 1121 129741 1225 129849
rect 1259 129707 1340 129815
rect 1121 129489 1340 129707
rect 1104 129455 1133 129489
rect 1167 129455 1225 129489
rect 1259 129455 1317 129489
rect 1121 129237 1340 129455
rect 1121 129095 1225 129203
rect 1259 129129 1340 129237
rect 1121 128945 1340 129095
rect 1104 128911 1133 128945
rect 1167 128911 1225 128945
rect 1259 128911 1317 128945
rect 1121 128761 1340 128911
rect 1121 128653 1225 128761
rect 1259 128619 1340 128727
rect 1121 128401 1340 128619
rect 1104 128367 1133 128401
rect 1167 128367 1225 128401
rect 1259 128367 1317 128401
rect 1121 128149 1340 128367
rect 1121 128007 1225 128115
rect 1259 128041 1340 128149
rect 1121 127857 1340 128007
rect 1104 127823 1133 127857
rect 1167 127823 1225 127857
rect 1259 127823 1317 127857
rect 1121 127673 1340 127823
rect 1121 127565 1225 127673
rect 1259 127531 1340 127639
rect 1121 127313 1340 127531
rect 1104 127279 1133 127313
rect 1167 127279 1225 127313
rect 1259 127279 1317 127313
rect 1121 127061 1340 127279
rect 1121 126919 1225 127027
rect 1259 126953 1340 127061
rect 1121 126769 1340 126919
rect 1104 126735 1133 126769
rect 1167 126735 1225 126769
rect 1259 126735 1317 126769
rect 1121 126585 1340 126735
rect 1121 126477 1225 126585
rect 1259 126443 1340 126551
rect 1121 126225 1340 126443
rect 1104 126191 1133 126225
rect 1167 126191 1225 126225
rect 1259 126191 1317 126225
rect 1121 125973 1340 126191
rect 1121 125831 1225 125939
rect 1259 125865 1340 125973
rect 1121 125681 1340 125831
rect 1104 125647 1133 125681
rect 1167 125647 1225 125681
rect 1259 125647 1317 125681
rect 1121 125497 1340 125647
rect 1121 125389 1225 125497
rect 1259 125355 1340 125463
rect 1121 125137 1340 125355
rect 1104 125103 1133 125137
rect 1167 125103 1225 125137
rect 1259 125103 1317 125137
rect 1121 124885 1340 125103
rect 1121 124743 1225 124851
rect 1259 124777 1340 124885
rect 1121 124593 1340 124743
rect 1104 124559 1133 124593
rect 1167 124559 1225 124593
rect 1259 124559 1317 124593
rect 1121 124409 1340 124559
rect 1121 124301 1225 124409
rect 1259 124267 1340 124375
rect 1121 124049 1340 124267
rect 1104 124015 1133 124049
rect 1167 124015 1225 124049
rect 1259 124015 1317 124049
rect 1121 123797 1340 124015
rect 1121 123655 1225 123763
rect 1259 123689 1340 123797
rect 1121 123505 1340 123655
rect 1104 123471 1133 123505
rect 1167 123471 1225 123505
rect 1259 123471 1317 123505
rect 1121 123321 1340 123471
rect 1121 123213 1225 123321
rect 1259 123179 1340 123287
rect 1121 122961 1340 123179
rect 1104 122927 1133 122961
rect 1167 122927 1225 122961
rect 1259 122927 1317 122961
rect 1121 122709 1340 122927
rect 1121 122567 1225 122675
rect 1259 122601 1340 122709
rect 1121 122417 1340 122567
rect 1104 122383 1133 122417
rect 1167 122383 1225 122417
rect 1259 122383 1317 122417
rect 1121 122233 1340 122383
rect 1121 122125 1225 122233
rect 1259 122091 1340 122199
rect 1121 121873 1340 122091
rect 1104 121839 1133 121873
rect 1167 121839 1225 121873
rect 1259 121839 1317 121873
rect 1121 121621 1340 121839
rect 1121 121479 1225 121587
rect 1259 121513 1340 121621
rect 1121 121329 1340 121479
rect 1104 121295 1133 121329
rect 1167 121295 1225 121329
rect 1259 121295 1317 121329
rect 1121 121145 1340 121295
rect 1121 121037 1225 121145
rect 1259 121003 1340 121111
rect 1121 120785 1340 121003
rect 1104 120751 1133 120785
rect 1167 120751 1225 120785
rect 1259 120751 1317 120785
rect 1121 120533 1340 120751
rect 1121 120391 1225 120499
rect 1259 120425 1340 120533
rect 1121 120241 1340 120391
rect 1104 120207 1133 120241
rect 1167 120207 1225 120241
rect 1259 120207 1317 120241
rect 1121 120057 1340 120207
rect 1121 119949 1225 120057
rect 1259 119915 1340 120023
rect 1121 119697 1340 119915
rect 1104 119663 1133 119697
rect 1167 119663 1225 119697
rect 1259 119663 1317 119697
rect 1121 119445 1340 119663
rect 1121 119303 1225 119411
rect 1259 119337 1340 119445
rect 1121 119153 1340 119303
rect 1104 119119 1133 119153
rect 1167 119119 1225 119153
rect 1259 119119 1317 119153
rect 1121 118969 1340 119119
rect 1121 118861 1225 118969
rect 1259 118827 1340 118935
rect 1121 118609 1340 118827
rect 1104 118575 1133 118609
rect 1167 118575 1225 118609
rect 1259 118575 1317 118609
rect 1121 118357 1340 118575
rect 1121 118215 1225 118323
rect 1259 118249 1340 118357
rect 1121 118065 1340 118215
rect 1104 118031 1133 118065
rect 1167 118031 1225 118065
rect 1259 118031 1317 118065
rect 1121 117881 1340 118031
rect 1121 117773 1225 117881
rect 1259 117739 1340 117847
rect 1121 117521 1340 117739
rect 1104 117487 1133 117521
rect 1167 117487 1225 117521
rect 1259 117487 1317 117521
rect 1121 117269 1340 117487
rect 1121 117127 1225 117235
rect 1259 117161 1340 117269
rect 1121 116977 1340 117127
rect 1104 116943 1133 116977
rect 1167 116943 1225 116977
rect 1259 116943 1317 116977
rect 1121 116793 1340 116943
rect 1121 116685 1225 116793
rect 1259 116651 1340 116759
rect 1121 116433 1340 116651
rect 1104 116399 1133 116433
rect 1167 116399 1225 116433
rect 1259 116399 1317 116433
rect 1121 116181 1340 116399
rect 1121 116039 1225 116147
rect 1259 116073 1340 116181
rect 1121 115889 1340 116039
rect 1104 115855 1133 115889
rect 1167 115855 1225 115889
rect 1259 115855 1317 115889
rect 1121 115705 1340 115855
rect 1121 115597 1225 115705
rect 1259 115563 1340 115671
rect 1121 115345 1340 115563
rect 1104 115311 1133 115345
rect 1167 115311 1225 115345
rect 1259 115311 1317 115345
rect 1121 115093 1340 115311
rect 1121 114951 1225 115059
rect 1259 114985 1340 115093
rect 1121 114801 1340 114951
rect 1104 114767 1133 114801
rect 1167 114767 1225 114801
rect 1259 114767 1317 114801
rect 1121 114617 1340 114767
rect 1121 114509 1225 114617
rect 1259 114475 1340 114583
rect 1121 114257 1340 114475
rect 1104 114223 1133 114257
rect 1167 114223 1225 114257
rect 1259 114223 1317 114257
rect 1121 114005 1340 114223
rect 1121 113863 1225 113971
rect 1259 113897 1340 114005
rect 1121 113713 1340 113863
rect 1104 113679 1133 113713
rect 1167 113679 1225 113713
rect 1259 113679 1317 113713
rect 1121 113529 1340 113679
rect 1121 113421 1225 113529
rect 1259 113387 1340 113495
rect 1121 113169 1340 113387
rect 1104 113135 1133 113169
rect 1167 113135 1225 113169
rect 1259 113135 1317 113169
rect 1121 112917 1340 113135
rect 1121 112775 1225 112883
rect 1259 112809 1340 112917
rect 1121 112625 1340 112775
rect 1104 112591 1133 112625
rect 1167 112591 1225 112625
rect 1259 112591 1317 112625
rect 1121 112441 1340 112591
rect 1121 112333 1225 112441
rect 1259 112299 1340 112407
rect 1121 112081 1340 112299
rect 1104 112047 1133 112081
rect 1167 112047 1225 112081
rect 1259 112047 1317 112081
rect 1121 111829 1340 112047
rect 1121 111687 1225 111795
rect 1259 111721 1340 111829
rect 1121 111537 1340 111687
rect 1104 111503 1133 111537
rect 1167 111503 1225 111537
rect 1259 111503 1317 111537
rect 1121 111353 1340 111503
rect 1121 111245 1225 111353
rect 1259 111211 1340 111319
rect 1121 110993 1340 111211
rect 1104 110959 1133 110993
rect 1167 110959 1225 110993
rect 1259 110959 1317 110993
rect 1121 110741 1340 110959
rect 1121 110599 1225 110707
rect 1259 110633 1340 110741
rect 1121 110449 1340 110599
rect 1104 110415 1133 110449
rect 1167 110415 1225 110449
rect 1259 110415 1317 110449
rect 1121 110265 1340 110415
rect 1121 110157 1225 110265
rect 1259 110123 1340 110231
rect 1121 109905 1340 110123
rect 1104 109871 1133 109905
rect 1167 109871 1225 109905
rect 1259 109871 1317 109905
rect 1121 109653 1340 109871
rect 1121 109511 1225 109619
rect 1259 109545 1340 109653
rect 1121 109361 1340 109511
rect 1104 109327 1133 109361
rect 1167 109327 1225 109361
rect 1259 109327 1317 109361
rect 1121 109177 1340 109327
rect 1121 109069 1225 109177
rect 1259 109035 1340 109143
rect 1121 108817 1340 109035
rect 1104 108783 1133 108817
rect 1167 108783 1225 108817
rect 1259 108783 1317 108817
rect 1121 108565 1340 108783
rect 1121 108423 1225 108531
rect 1259 108457 1340 108565
rect 1121 108273 1340 108423
rect 1104 108239 1133 108273
rect 1167 108239 1225 108273
rect 1259 108239 1317 108273
rect 1121 108089 1340 108239
rect 1121 107981 1225 108089
rect 1259 107947 1340 108055
rect 1121 107729 1340 107947
rect 1104 107695 1133 107729
rect 1167 107695 1225 107729
rect 1259 107695 1317 107729
rect 1121 107477 1340 107695
rect 1121 107335 1225 107443
rect 1259 107369 1340 107477
rect 1121 107185 1340 107335
rect 1104 107151 1133 107185
rect 1167 107151 1225 107185
rect 1259 107151 1317 107185
rect 1121 107001 1340 107151
rect 1121 106893 1225 107001
rect 1259 106859 1340 106967
rect 1121 106641 1340 106859
rect 1104 106607 1133 106641
rect 1167 106607 1225 106641
rect 1259 106607 1317 106641
rect 1121 106389 1340 106607
rect 1121 106247 1225 106355
rect 1259 106281 1340 106389
rect 1121 106097 1340 106247
rect 1104 106063 1133 106097
rect 1167 106063 1225 106097
rect 1259 106063 1317 106097
rect 1121 105913 1340 106063
rect 1121 105805 1225 105913
rect 1259 105771 1340 105879
rect 1121 105553 1340 105771
rect 1104 105519 1133 105553
rect 1167 105519 1225 105553
rect 1259 105519 1317 105553
rect 1121 105301 1340 105519
rect 1121 105159 1225 105267
rect 1259 105193 1340 105301
rect 1121 105009 1340 105159
rect 1104 104975 1133 105009
rect 1167 104975 1225 105009
rect 1259 104975 1317 105009
rect 1121 104825 1340 104975
rect 1121 104717 1225 104825
rect 1259 104683 1340 104791
rect 1121 104465 1340 104683
rect 1104 104431 1133 104465
rect 1167 104431 1225 104465
rect 1259 104431 1317 104465
rect 1121 104213 1340 104431
rect 1121 104071 1225 104179
rect 1259 104105 1340 104213
rect 1121 103921 1340 104071
rect 1104 103887 1133 103921
rect 1167 103887 1225 103921
rect 1259 103887 1317 103921
rect 1121 103737 1340 103887
rect 1121 103629 1225 103737
rect 1259 103595 1340 103703
rect 1121 103377 1340 103595
rect 1104 103343 1133 103377
rect 1167 103343 1225 103377
rect 1259 103343 1317 103377
rect 1121 103125 1340 103343
rect 1121 102983 1225 103091
rect 1259 103017 1340 103125
rect 1121 102833 1340 102983
rect 1104 102799 1133 102833
rect 1167 102799 1225 102833
rect 1259 102799 1317 102833
rect 1121 102649 1340 102799
rect 1121 102541 1225 102649
rect 1259 102507 1340 102615
rect 1121 102289 1340 102507
rect 1104 102255 1133 102289
rect 1167 102255 1225 102289
rect 1259 102255 1317 102289
rect 1121 102037 1340 102255
rect 1121 101895 1225 102003
rect 1259 101929 1340 102037
rect 1121 101745 1340 101895
rect 1104 101711 1133 101745
rect 1167 101711 1225 101745
rect 1259 101711 1317 101745
rect 1121 101561 1340 101711
rect 1121 101453 1225 101561
rect 1259 101419 1340 101527
rect 1121 101201 1340 101419
rect 1104 101167 1133 101201
rect 1167 101167 1225 101201
rect 1259 101167 1317 101201
rect 1121 100949 1340 101167
rect 1121 100807 1225 100915
rect 1259 100841 1340 100949
rect 1121 100657 1340 100807
rect 1104 100623 1133 100657
rect 1167 100623 1225 100657
rect 1259 100623 1317 100657
rect 1121 100473 1340 100623
rect 1121 100365 1225 100473
rect 1259 100331 1340 100439
rect 1121 100113 1340 100331
rect 1104 100079 1133 100113
rect 1167 100079 1225 100113
rect 1259 100079 1317 100113
rect 1121 99861 1340 100079
rect 1121 99719 1225 99827
rect 1259 99753 1340 99861
rect 1121 99569 1340 99719
rect 1104 99535 1133 99569
rect 1167 99535 1225 99569
rect 1259 99535 1317 99569
rect 1121 99385 1340 99535
rect 1121 99277 1225 99385
rect 1259 99243 1340 99351
rect 1121 99025 1340 99243
rect 1104 98991 1133 99025
rect 1167 98991 1225 99025
rect 1259 98991 1317 99025
rect 1121 98773 1340 98991
rect 1121 98631 1225 98739
rect 1259 98665 1340 98773
rect 1121 98481 1340 98631
rect 1104 98447 1133 98481
rect 1167 98447 1225 98481
rect 1259 98447 1317 98481
rect 1121 98297 1340 98447
rect 1121 98189 1225 98297
rect 1259 98155 1340 98263
rect 1121 97937 1340 98155
rect 1104 97903 1133 97937
rect 1167 97903 1225 97937
rect 1259 97903 1317 97937
rect 1121 97685 1340 97903
rect 1121 97543 1225 97651
rect 1259 97577 1340 97685
rect 1121 97393 1340 97543
rect 1104 97359 1133 97393
rect 1167 97359 1225 97393
rect 1259 97359 1317 97393
rect 1121 97209 1340 97359
rect 1121 97101 1225 97209
rect 1259 97067 1340 97175
rect 1121 96849 1340 97067
rect 1104 96815 1133 96849
rect 1167 96815 1225 96849
rect 1259 96815 1317 96849
rect 1121 96597 1340 96815
rect 1121 96455 1225 96563
rect 1259 96489 1340 96597
rect 1121 96305 1340 96455
rect 1104 96271 1133 96305
rect 1167 96271 1225 96305
rect 1259 96271 1317 96305
rect 1121 96121 1340 96271
rect 1121 96013 1225 96121
rect 1259 95979 1340 96087
rect 1121 95761 1340 95979
rect 1104 95727 1133 95761
rect 1167 95727 1225 95761
rect 1259 95727 1317 95761
rect 1121 95509 1340 95727
rect 1121 95367 1225 95475
rect 1259 95401 1340 95509
rect 1121 95217 1340 95367
rect 1104 95183 1133 95217
rect 1167 95183 1225 95217
rect 1259 95183 1317 95217
rect 1121 95033 1340 95183
rect 1121 94925 1225 95033
rect 1259 94891 1340 94999
rect 1121 94673 1340 94891
rect 1104 94639 1133 94673
rect 1167 94639 1225 94673
rect 1259 94639 1317 94673
rect 1121 94421 1340 94639
rect 1121 94279 1225 94387
rect 1259 94313 1340 94421
rect 1121 94129 1340 94279
rect 1104 94095 1133 94129
rect 1167 94095 1225 94129
rect 1259 94095 1317 94129
rect 1121 93945 1340 94095
rect 1121 93837 1225 93945
rect 1259 93803 1340 93911
rect 1121 93585 1340 93803
rect 1104 93551 1133 93585
rect 1167 93551 1225 93585
rect 1259 93551 1317 93585
rect 1121 93333 1340 93551
rect 1121 93191 1225 93299
rect 1259 93225 1340 93333
rect 1121 93041 1340 93191
rect 1104 93007 1133 93041
rect 1167 93007 1225 93041
rect 1259 93007 1317 93041
rect 1121 92857 1340 93007
rect 1121 92749 1225 92857
rect 1259 92715 1340 92823
rect 1121 92497 1340 92715
rect 1104 92463 1133 92497
rect 1167 92463 1225 92497
rect 1259 92463 1317 92497
rect 1121 92245 1340 92463
rect 1121 92103 1225 92211
rect 1259 92137 1340 92245
rect 1121 91953 1340 92103
rect 1104 91919 1133 91953
rect 1167 91919 1225 91953
rect 1259 91919 1317 91953
rect 1121 91769 1340 91919
rect 1121 91661 1225 91769
rect 1259 91627 1340 91735
rect 1121 91409 1340 91627
rect 1104 91375 1133 91409
rect 1167 91375 1225 91409
rect 1259 91375 1317 91409
rect 1121 91157 1340 91375
rect 1121 91015 1225 91123
rect 1259 91049 1340 91157
rect 1121 90865 1340 91015
rect 1104 90831 1133 90865
rect 1167 90831 1225 90865
rect 1259 90831 1317 90865
rect 1121 90681 1340 90831
rect 1121 90573 1225 90681
rect 1259 90539 1340 90647
rect 1121 90321 1340 90539
rect 1104 90287 1133 90321
rect 1167 90287 1225 90321
rect 1259 90287 1317 90321
rect 1121 90069 1340 90287
rect 1121 89927 1225 90035
rect 1259 89961 1340 90069
rect 1121 89777 1340 89927
rect 1104 89743 1133 89777
rect 1167 89743 1225 89777
rect 1259 89743 1317 89777
rect 1121 89593 1340 89743
rect 1121 89485 1225 89593
rect 1259 89451 1340 89559
rect 1121 89233 1340 89451
rect 1104 89199 1133 89233
rect 1167 89199 1225 89233
rect 1259 89199 1317 89233
rect 1121 88981 1340 89199
rect 1121 88839 1225 88947
rect 1259 88873 1340 88981
rect 1121 88689 1340 88839
rect 1104 88655 1133 88689
rect 1167 88655 1225 88689
rect 1259 88655 1317 88689
rect 1121 88505 1340 88655
rect 1121 88397 1225 88505
rect 1259 88363 1340 88471
rect 1121 88145 1340 88363
rect 1104 88111 1133 88145
rect 1167 88111 1225 88145
rect 1259 88111 1317 88145
rect 1121 87893 1340 88111
rect 1121 87751 1225 87859
rect 1259 87785 1340 87893
rect 1121 87601 1340 87751
rect 1104 87567 1133 87601
rect 1167 87567 1225 87601
rect 1259 87567 1317 87601
rect 1121 87417 1340 87567
rect 1121 87309 1225 87417
rect 1259 87275 1340 87383
rect 1121 87057 1340 87275
rect 1104 87023 1133 87057
rect 1167 87023 1225 87057
rect 1259 87023 1317 87057
rect 1121 86805 1340 87023
rect 1121 86663 1225 86771
rect 1259 86697 1340 86805
rect 1121 86513 1340 86663
rect 1104 86479 1133 86513
rect 1167 86479 1225 86513
rect 1259 86479 1317 86513
rect 1121 86329 1340 86479
rect 1121 86221 1225 86329
rect 1259 86187 1340 86295
rect 1121 85969 1340 86187
rect 1104 85935 1133 85969
rect 1167 85935 1225 85969
rect 1259 85935 1317 85969
rect 1121 85717 1340 85935
rect 1121 85575 1225 85683
rect 1259 85609 1340 85717
rect 1121 85425 1340 85575
rect 1104 85391 1133 85425
rect 1167 85391 1225 85425
rect 1259 85391 1317 85425
rect 1121 85241 1340 85391
rect 1121 85133 1225 85241
rect 1259 85099 1340 85207
rect 1121 84881 1340 85099
rect 1104 84847 1133 84881
rect 1167 84847 1225 84881
rect 1259 84847 1317 84881
rect 1121 84629 1340 84847
rect 1121 84487 1225 84595
rect 1259 84521 1340 84629
rect 1121 84337 1340 84487
rect 1104 84303 1133 84337
rect 1167 84303 1225 84337
rect 1259 84303 1317 84337
rect 1121 84153 1340 84303
rect 1121 84045 1225 84153
rect 1259 84011 1340 84119
rect 1121 83793 1340 84011
rect 1104 83759 1133 83793
rect 1167 83759 1225 83793
rect 1259 83759 1317 83793
rect 1121 83541 1340 83759
rect 1121 83399 1225 83507
rect 1259 83433 1340 83541
rect 1121 83249 1340 83399
rect 1104 83215 1133 83249
rect 1167 83215 1225 83249
rect 1259 83215 1317 83249
rect 1121 83065 1340 83215
rect 1121 82957 1225 83065
rect 1259 82923 1340 83031
rect 1121 82705 1340 82923
rect 1104 82671 1133 82705
rect 1167 82671 1225 82705
rect 1259 82671 1317 82705
rect 1121 82453 1340 82671
rect 1121 82311 1225 82419
rect 1259 82345 1340 82453
rect 1121 82161 1340 82311
rect 1104 82127 1133 82161
rect 1167 82127 1225 82161
rect 1259 82127 1317 82161
rect 1121 81977 1340 82127
rect 1121 81869 1225 81977
rect 1259 81835 1340 81943
rect 1121 81617 1340 81835
rect 1104 81583 1133 81617
rect 1167 81583 1225 81617
rect 1259 81583 1317 81617
rect 1121 81365 1340 81583
rect 1121 81223 1225 81331
rect 1259 81257 1340 81365
rect 1121 81073 1340 81223
rect 1104 81039 1133 81073
rect 1167 81039 1225 81073
rect 1259 81039 1317 81073
rect 1121 80889 1340 81039
rect 1121 80781 1225 80889
rect 1259 80747 1340 80855
rect 1121 80529 1340 80747
rect 1104 80495 1133 80529
rect 1167 80495 1225 80529
rect 1259 80495 1317 80529
rect 1121 80277 1340 80495
rect 1121 80135 1225 80243
rect 1259 80169 1340 80277
rect 1121 79985 1340 80135
rect 1104 79951 1133 79985
rect 1167 79951 1225 79985
rect 1259 79951 1317 79985
rect 1121 79801 1340 79951
rect 1121 79693 1225 79801
rect 1259 79659 1340 79767
rect 1121 79441 1340 79659
rect 1104 79407 1133 79441
rect 1167 79407 1225 79441
rect 1259 79407 1317 79441
rect 1121 79189 1340 79407
rect 1121 79047 1225 79155
rect 1259 79081 1340 79189
rect 1121 78897 1340 79047
rect 1104 78863 1133 78897
rect 1167 78863 1225 78897
rect 1259 78863 1317 78897
rect 1121 78713 1340 78863
rect 1121 78605 1225 78713
rect 1259 78571 1340 78679
rect 1121 78353 1340 78571
rect 1104 78319 1133 78353
rect 1167 78319 1225 78353
rect 1259 78319 1317 78353
rect 1121 78101 1340 78319
rect 1121 77959 1225 78067
rect 1259 77993 1340 78101
rect 1121 77809 1340 77959
rect 1104 77775 1133 77809
rect 1167 77775 1225 77809
rect 1259 77775 1317 77809
rect 1121 77625 1340 77775
rect 1121 77517 1225 77625
rect 1259 77483 1340 77591
rect 1121 77265 1340 77483
rect 1104 77231 1133 77265
rect 1167 77231 1225 77265
rect 1259 77231 1317 77265
rect 1121 77013 1340 77231
rect 1121 76871 1225 76979
rect 1259 76905 1340 77013
rect 1121 76721 1340 76871
rect 1104 76687 1133 76721
rect 1167 76687 1225 76721
rect 1259 76687 1317 76721
rect 1121 76537 1340 76687
rect 1121 76429 1225 76537
rect 1259 76395 1340 76503
rect 1121 76177 1340 76395
rect 1104 76143 1133 76177
rect 1167 76143 1225 76177
rect 1259 76143 1317 76177
rect 1121 75925 1340 76143
rect 1121 75783 1225 75891
rect 1259 75817 1340 75925
rect 1121 75633 1340 75783
rect 1104 75599 1133 75633
rect 1167 75599 1225 75633
rect 1259 75599 1317 75633
rect 1121 75449 1340 75599
rect 1121 75341 1225 75449
rect 1259 75307 1340 75415
rect 1121 75089 1340 75307
rect 1104 75055 1133 75089
rect 1167 75055 1225 75089
rect 1259 75055 1317 75089
rect 1121 74837 1340 75055
rect 1121 74695 1225 74803
rect 1259 74729 1340 74837
rect 1121 74545 1340 74695
rect 1104 74511 1133 74545
rect 1167 74511 1225 74545
rect 1259 74511 1317 74545
rect 1121 74361 1340 74511
rect 1121 74253 1225 74361
rect 1259 74219 1340 74327
rect 1121 74001 1340 74219
rect 1104 73967 1133 74001
rect 1167 73967 1225 74001
rect 1259 73967 1317 74001
rect 1121 73749 1340 73967
rect 1121 73607 1225 73715
rect 1259 73641 1340 73749
rect 1121 73457 1340 73607
rect 1104 73423 1133 73457
rect 1167 73423 1225 73457
rect 1259 73423 1317 73457
rect 1121 73273 1340 73423
rect 1121 73165 1225 73273
rect 1259 73131 1340 73239
rect 1121 72913 1340 73131
rect 1104 72879 1133 72913
rect 1167 72879 1225 72913
rect 1259 72879 1317 72913
rect 1121 72661 1340 72879
rect 1121 72519 1225 72627
rect 1259 72553 1340 72661
rect 1121 72369 1340 72519
rect 1104 72335 1133 72369
rect 1167 72335 1225 72369
rect 1259 72335 1317 72369
rect 1121 72185 1340 72335
rect 1121 72077 1225 72185
rect 1259 72043 1340 72151
rect 1121 71825 1340 72043
rect 1104 71791 1133 71825
rect 1167 71791 1225 71825
rect 1259 71791 1317 71825
rect 1121 71573 1340 71791
rect 1121 71431 1225 71539
rect 1259 71465 1340 71573
rect 1121 71281 1340 71431
rect 1104 71247 1133 71281
rect 1167 71247 1225 71281
rect 1259 71247 1317 71281
rect 1121 71097 1340 71247
rect 1121 70989 1225 71097
rect 1259 70955 1340 71063
rect 1121 70737 1340 70955
rect 1104 70703 1133 70737
rect 1167 70703 1225 70737
rect 1259 70703 1317 70737
rect 1121 70485 1340 70703
rect 1121 70343 1225 70451
rect 1259 70377 1340 70485
rect 1121 70193 1340 70343
rect 1104 70159 1133 70193
rect 1167 70159 1225 70193
rect 1259 70159 1317 70193
rect 1121 70009 1340 70159
rect 1121 69901 1225 70009
rect 1259 69867 1340 69975
rect 1121 69649 1340 69867
rect 1104 69615 1133 69649
rect 1167 69615 1225 69649
rect 1259 69615 1317 69649
rect 1121 69397 1340 69615
rect 1121 69255 1225 69363
rect 1259 69289 1340 69397
rect 1121 69105 1340 69255
rect 1104 69071 1133 69105
rect 1167 69071 1225 69105
rect 1259 69071 1317 69105
rect 1121 68921 1340 69071
rect 1121 68813 1225 68921
rect 1259 68779 1340 68887
rect 1121 68561 1340 68779
rect 1104 68527 1133 68561
rect 1167 68527 1225 68561
rect 1259 68527 1317 68561
rect 1121 68309 1340 68527
rect 1121 68167 1225 68275
rect 1259 68201 1340 68309
rect 1121 68017 1340 68167
rect 1104 67983 1133 68017
rect 1167 67983 1225 68017
rect 1259 67983 1317 68017
rect 1121 67833 1340 67983
rect 1121 67725 1225 67833
rect 1259 67691 1340 67799
rect 1121 67473 1340 67691
rect 1104 67439 1133 67473
rect 1167 67439 1225 67473
rect 1259 67439 1317 67473
rect 1121 67221 1340 67439
rect 1121 67079 1225 67187
rect 1259 67113 1340 67221
rect 1121 66929 1340 67079
rect 1104 66895 1133 66929
rect 1167 66895 1225 66929
rect 1259 66895 1317 66929
rect 1121 66745 1340 66895
rect 1121 66637 1225 66745
rect 1259 66603 1340 66711
rect 1121 66385 1340 66603
rect 1104 66351 1133 66385
rect 1167 66351 1225 66385
rect 1259 66351 1317 66385
rect 1121 66133 1340 66351
rect 1121 65991 1225 66099
rect 1259 66025 1340 66133
rect 1121 65841 1340 65991
rect 1104 65807 1133 65841
rect 1167 65807 1225 65841
rect 1259 65807 1317 65841
rect 1121 65657 1340 65807
rect 1121 65549 1225 65657
rect 1259 65515 1340 65623
rect 1121 65297 1340 65515
rect 1104 65263 1133 65297
rect 1167 65263 1225 65297
rect 1259 65263 1317 65297
rect 1121 65045 1340 65263
rect 1121 64903 1225 65011
rect 1259 64937 1340 65045
rect 1121 64753 1340 64903
rect 1104 64719 1133 64753
rect 1167 64719 1225 64753
rect 1259 64719 1317 64753
rect 1121 64569 1340 64719
rect 1121 64461 1225 64569
rect 1259 64427 1340 64535
rect 1121 64209 1340 64427
rect 1104 64175 1133 64209
rect 1167 64175 1225 64209
rect 1259 64175 1317 64209
rect 1121 63957 1340 64175
rect 1121 63815 1225 63923
rect 1259 63849 1340 63957
rect 1121 63665 1340 63815
rect 1104 63631 1133 63665
rect 1167 63631 1225 63665
rect 1259 63631 1317 63665
rect 1121 63481 1340 63631
rect 1121 63373 1225 63481
rect 1259 63339 1340 63447
rect 1121 63121 1340 63339
rect 1104 63087 1133 63121
rect 1167 63087 1225 63121
rect 1259 63087 1317 63121
rect 1121 62869 1340 63087
rect 1121 62727 1225 62835
rect 1259 62761 1340 62869
rect 1121 62577 1340 62727
rect 1104 62543 1133 62577
rect 1167 62543 1225 62577
rect 1259 62543 1317 62577
rect 1121 62393 1340 62543
rect 1121 62285 1225 62393
rect 1259 62251 1340 62359
rect 1121 62033 1340 62251
rect 1104 61999 1133 62033
rect 1167 61999 1225 62033
rect 1259 61999 1317 62033
rect 1121 61781 1340 61999
rect 1121 61639 1225 61747
rect 1259 61673 1340 61781
rect 1121 61489 1340 61639
rect 1104 61455 1133 61489
rect 1167 61455 1225 61489
rect 1259 61455 1317 61489
rect 1121 61305 1340 61455
rect 1121 61197 1225 61305
rect 1259 61163 1340 61271
rect 1121 60945 1340 61163
rect 1104 60911 1133 60945
rect 1167 60911 1225 60945
rect 1259 60911 1317 60945
rect 1121 60693 1340 60911
rect 1121 60551 1225 60659
rect 1259 60585 1340 60693
rect 1121 60401 1340 60551
rect 1104 60367 1133 60401
rect 1167 60367 1225 60401
rect 1259 60367 1317 60401
rect 1121 60217 1340 60367
rect 1121 60109 1225 60217
rect 1259 60075 1340 60183
rect 1121 59857 1340 60075
rect 1104 59823 1133 59857
rect 1167 59823 1225 59857
rect 1259 59823 1317 59857
rect 1121 59605 1340 59823
rect 1121 59463 1225 59571
rect 1259 59497 1340 59605
rect 1121 59313 1340 59463
rect 1104 59279 1133 59313
rect 1167 59279 1225 59313
rect 1259 59279 1317 59313
rect 1121 59129 1340 59279
rect 1121 59021 1225 59129
rect 1259 58987 1340 59095
rect 1121 58769 1340 58987
rect 1104 58735 1133 58769
rect 1167 58735 1225 58769
rect 1259 58735 1317 58769
rect 1121 58517 1340 58735
rect 1121 58375 1225 58483
rect 1259 58409 1340 58517
rect 1121 58225 1340 58375
rect 1104 58191 1133 58225
rect 1167 58191 1225 58225
rect 1259 58191 1317 58225
rect 1121 58041 1340 58191
rect 1121 57933 1225 58041
rect 1259 57899 1340 58007
rect 1121 57681 1340 57899
rect 1104 57647 1133 57681
rect 1167 57647 1225 57681
rect 1259 57647 1317 57681
rect 1121 57429 1340 57647
rect 1121 57287 1225 57395
rect 1259 57321 1340 57429
rect 1121 57137 1340 57287
rect 1104 57103 1133 57137
rect 1167 57103 1225 57137
rect 1259 57103 1317 57137
rect 1121 56953 1340 57103
rect 1121 56845 1225 56953
rect 1259 56811 1340 56919
rect 1121 56593 1340 56811
rect 1104 56559 1133 56593
rect 1167 56559 1225 56593
rect 1259 56559 1317 56593
rect 1121 56341 1340 56559
rect 1121 56199 1225 56307
rect 1259 56233 1340 56341
rect 1121 56049 1340 56199
rect 1104 56015 1133 56049
rect 1167 56015 1225 56049
rect 1259 56015 1317 56049
rect 1121 55865 1340 56015
rect 1121 55757 1225 55865
rect 1259 55723 1340 55831
rect 1121 55505 1340 55723
rect 1104 55471 1133 55505
rect 1167 55471 1225 55505
rect 1259 55471 1317 55505
rect 1121 55253 1340 55471
rect 1121 55111 1225 55219
rect 1259 55145 1340 55253
rect 1121 54961 1340 55111
rect 1104 54927 1133 54961
rect 1167 54927 1225 54961
rect 1259 54927 1317 54961
rect 1121 54777 1340 54927
rect 1121 54669 1225 54777
rect 1259 54635 1340 54743
rect 1121 54417 1340 54635
rect 1104 54383 1133 54417
rect 1167 54383 1225 54417
rect 1259 54383 1317 54417
rect 1121 54165 1340 54383
rect 1121 54023 1225 54131
rect 1259 54057 1340 54165
rect 1121 53873 1340 54023
rect 1104 53839 1133 53873
rect 1167 53839 1225 53873
rect 1259 53839 1317 53873
rect 1121 53689 1340 53839
rect 1121 53581 1225 53689
rect 1259 53547 1340 53655
rect 1121 53329 1340 53547
rect 1104 53295 1133 53329
rect 1167 53295 1225 53329
rect 1259 53295 1317 53329
rect 1121 53077 1340 53295
rect 1121 52935 1225 53043
rect 1259 52969 1340 53077
rect 1121 52785 1340 52935
rect 1104 52751 1133 52785
rect 1167 52751 1225 52785
rect 1259 52751 1317 52785
rect 1121 52601 1340 52751
rect 1121 52493 1225 52601
rect 1259 52459 1340 52567
rect 1121 52241 1340 52459
rect 1104 52207 1133 52241
rect 1167 52207 1225 52241
rect 1259 52207 1317 52241
rect 1121 51989 1340 52207
rect 1121 51847 1225 51955
rect 1259 51881 1340 51989
rect 1121 51697 1340 51847
rect 1104 51663 1133 51697
rect 1167 51663 1225 51697
rect 1259 51663 1317 51697
rect 1121 51513 1340 51663
rect 1121 51405 1225 51513
rect 1259 51371 1340 51479
rect 1121 51153 1340 51371
rect 1104 51119 1133 51153
rect 1167 51119 1225 51153
rect 1259 51119 1317 51153
rect 1121 50901 1340 51119
rect 1121 50759 1225 50867
rect 1259 50793 1340 50901
rect 1121 50609 1340 50759
rect 1104 50575 1133 50609
rect 1167 50575 1225 50609
rect 1259 50575 1317 50609
rect 1121 50425 1340 50575
rect 1121 50317 1225 50425
rect 1259 50283 1340 50391
rect 1121 50065 1340 50283
rect 1104 50031 1133 50065
rect 1167 50031 1225 50065
rect 1259 50031 1317 50065
rect 1121 49813 1340 50031
rect 1121 49671 1225 49779
rect 1259 49705 1340 49813
rect 1121 49521 1340 49671
rect 1104 49487 1133 49521
rect 1167 49487 1225 49521
rect 1259 49487 1317 49521
rect 1121 49337 1340 49487
rect 1121 49229 1225 49337
rect 1259 49195 1340 49303
rect 1121 48977 1340 49195
rect 1104 48943 1133 48977
rect 1167 48943 1225 48977
rect 1259 48943 1317 48977
rect 1121 48725 1340 48943
rect 1121 48583 1225 48691
rect 1259 48617 1340 48725
rect 1121 48433 1340 48583
rect 1104 48399 1133 48433
rect 1167 48399 1225 48433
rect 1259 48399 1317 48433
rect 1121 48249 1340 48399
rect 1121 48141 1225 48249
rect 1259 48107 1340 48215
rect 1121 47889 1340 48107
rect 1104 47855 1133 47889
rect 1167 47855 1225 47889
rect 1259 47855 1317 47889
rect 1121 47637 1340 47855
rect 1121 47495 1225 47603
rect 1259 47529 1340 47637
rect 1121 47345 1340 47495
rect 1104 47311 1133 47345
rect 1167 47311 1225 47345
rect 1259 47311 1317 47345
rect 1121 47161 1340 47311
rect 1121 47053 1225 47161
rect 1259 47019 1340 47127
rect 1121 46801 1340 47019
rect 1104 46767 1133 46801
rect 1167 46767 1225 46801
rect 1259 46767 1317 46801
rect 1121 46549 1340 46767
rect 1121 46407 1225 46515
rect 1259 46441 1340 46549
rect 1121 46257 1340 46407
rect 1104 46223 1133 46257
rect 1167 46223 1225 46257
rect 1259 46223 1317 46257
rect 1121 46073 1340 46223
rect 1121 45965 1225 46073
rect 1259 45931 1340 46039
rect 1121 45713 1340 45931
rect 1104 45679 1133 45713
rect 1167 45679 1225 45713
rect 1259 45679 1317 45713
rect 1121 45461 1340 45679
rect 1121 45319 1225 45427
rect 1259 45353 1340 45461
rect 1121 45169 1340 45319
rect 1104 45135 1133 45169
rect 1167 45135 1225 45169
rect 1259 45135 1317 45169
rect 1121 44985 1340 45135
rect 1121 44877 1225 44985
rect 1259 44843 1340 44951
rect 1121 44625 1340 44843
rect 1104 44591 1133 44625
rect 1167 44591 1225 44625
rect 1259 44591 1317 44625
rect 1121 44373 1340 44591
rect 1121 44231 1225 44339
rect 1259 44265 1340 44373
rect 1121 44081 1340 44231
rect 1104 44047 1133 44081
rect 1167 44047 1225 44081
rect 1259 44047 1317 44081
rect 1121 43897 1340 44047
rect 1121 43789 1225 43897
rect 1259 43755 1340 43863
rect 1121 43537 1340 43755
rect 1104 43503 1133 43537
rect 1167 43503 1225 43537
rect 1259 43503 1317 43537
rect 1121 43285 1340 43503
rect 1121 43143 1225 43251
rect 1259 43177 1340 43285
rect 1121 42993 1340 43143
rect 1104 42959 1133 42993
rect 1167 42959 1225 42993
rect 1259 42959 1317 42993
rect 1121 42809 1340 42959
rect 1121 42701 1225 42809
rect 1259 42667 1340 42775
rect 1121 42449 1340 42667
rect 1104 42415 1133 42449
rect 1167 42415 1225 42449
rect 1259 42415 1317 42449
rect 1121 42197 1340 42415
rect 1121 42055 1225 42163
rect 1259 42089 1340 42197
rect 1121 41905 1340 42055
rect 1104 41871 1133 41905
rect 1167 41871 1225 41905
rect 1259 41871 1317 41905
rect 1121 41721 1340 41871
rect 1121 41613 1225 41721
rect 1259 41579 1340 41687
rect 1121 41361 1340 41579
rect 1104 41327 1133 41361
rect 1167 41327 1225 41361
rect 1259 41327 1317 41361
rect 1121 41109 1340 41327
rect 1121 40967 1225 41075
rect 1259 41001 1340 41109
rect 1121 40817 1340 40967
rect 1104 40783 1133 40817
rect 1167 40783 1225 40817
rect 1259 40783 1317 40817
rect 1121 40633 1340 40783
rect 1121 40525 1225 40633
rect 1259 40491 1340 40599
rect 1121 40273 1340 40491
rect 1104 40239 1133 40273
rect 1167 40239 1225 40273
rect 1259 40239 1317 40273
rect 1121 40021 1340 40239
rect 1121 39879 1225 39987
rect 1259 39913 1340 40021
rect 1121 39729 1340 39879
rect 1104 39695 1133 39729
rect 1167 39695 1225 39729
rect 1259 39695 1317 39729
rect 1121 39545 1340 39695
rect 1121 39437 1225 39545
rect 1259 39403 1340 39511
rect 1121 39185 1340 39403
rect 1104 39151 1133 39185
rect 1167 39151 1225 39185
rect 1259 39151 1317 39185
rect 1121 38933 1340 39151
rect 1121 38791 1225 38899
rect 1259 38825 1340 38933
rect 1121 38641 1340 38791
rect 1104 38607 1133 38641
rect 1167 38607 1225 38641
rect 1259 38607 1317 38641
rect 1121 38457 1340 38607
rect 1121 38349 1225 38457
rect 1259 38315 1340 38423
rect 1121 38097 1340 38315
rect 1104 38063 1133 38097
rect 1167 38063 1225 38097
rect 1259 38063 1317 38097
rect 1121 37845 1340 38063
rect 1121 37703 1225 37811
rect 1259 37737 1340 37845
rect 1121 37553 1340 37703
rect 1104 37519 1133 37553
rect 1167 37519 1225 37553
rect 1259 37519 1317 37553
rect 1121 37369 1340 37519
rect 1121 37261 1225 37369
rect 1259 37227 1340 37335
rect 1121 37009 1340 37227
rect 1104 36975 1133 37009
rect 1167 36975 1225 37009
rect 1259 36975 1317 37009
rect 1121 36757 1340 36975
rect 1121 36615 1225 36723
rect 1259 36649 1340 36757
rect 1121 36465 1340 36615
rect 1104 36431 1133 36465
rect 1167 36431 1225 36465
rect 1259 36431 1317 36465
rect 1121 36281 1340 36431
rect 1121 36173 1225 36281
rect 1259 36139 1340 36247
rect 1121 35921 1340 36139
rect 1104 35887 1133 35921
rect 1167 35887 1225 35921
rect 1259 35887 1317 35921
rect 1121 35669 1340 35887
rect 1121 35527 1225 35635
rect 1259 35561 1340 35669
rect 1121 35377 1340 35527
rect 1104 35343 1133 35377
rect 1167 35343 1225 35377
rect 1259 35343 1317 35377
rect 1121 35193 1340 35343
rect 1121 35085 1225 35193
rect 1259 35051 1340 35159
rect 1121 34833 1340 35051
rect 1104 34799 1133 34833
rect 1167 34799 1225 34833
rect 1259 34799 1317 34833
rect 1121 34581 1340 34799
rect 1121 34439 1225 34547
rect 1259 34473 1340 34581
rect 1121 34289 1340 34439
rect 1104 34255 1133 34289
rect 1167 34255 1225 34289
rect 1259 34255 1317 34289
rect 1121 34105 1340 34255
rect 1121 33997 1225 34105
rect 1259 33963 1340 34071
rect 1121 33745 1340 33963
rect 1104 33711 1133 33745
rect 1167 33711 1225 33745
rect 1259 33711 1317 33745
rect 1121 33493 1340 33711
rect 1121 33351 1225 33459
rect 1259 33385 1340 33493
rect 1121 33201 1340 33351
rect 1104 33167 1133 33201
rect 1167 33167 1225 33201
rect 1259 33167 1317 33201
rect 1121 33017 1340 33167
rect 1121 32909 1225 33017
rect 1259 32875 1340 32983
rect 1121 32657 1340 32875
rect 1104 32623 1133 32657
rect 1167 32623 1225 32657
rect 1259 32623 1317 32657
rect 1121 32405 1340 32623
rect 1121 32263 1225 32371
rect 1259 32297 1340 32405
rect 1121 32113 1340 32263
rect 1104 32079 1133 32113
rect 1167 32079 1225 32113
rect 1259 32079 1317 32113
rect 1121 31929 1340 32079
rect 1121 31821 1225 31929
rect 1259 31787 1340 31895
rect 1121 31569 1340 31787
rect 1104 31535 1133 31569
rect 1167 31535 1225 31569
rect 1259 31535 1317 31569
rect 1121 31317 1340 31535
rect 1121 31175 1225 31283
rect 1259 31209 1340 31317
rect 1121 31025 1340 31175
rect 1104 30991 1133 31025
rect 1167 30991 1225 31025
rect 1259 30991 1317 31025
rect 1121 30841 1340 30991
rect 1121 30733 1225 30841
rect 1259 30699 1340 30807
rect 1121 30481 1340 30699
rect 1104 30447 1133 30481
rect 1167 30447 1225 30481
rect 1259 30447 1317 30481
rect 1121 30229 1340 30447
rect 1121 30087 1225 30195
rect 1259 30121 1340 30229
rect 1121 29937 1340 30087
rect 1104 29903 1133 29937
rect 1167 29903 1225 29937
rect 1259 29903 1317 29937
rect 1121 29753 1340 29903
rect 1121 29645 1225 29753
rect 1259 29611 1340 29719
rect 1121 29393 1340 29611
rect 1104 29359 1133 29393
rect 1167 29359 1225 29393
rect 1259 29359 1317 29393
rect 1121 29141 1340 29359
rect 1121 28999 1225 29107
rect 1259 29033 1340 29141
rect 1121 28849 1340 28999
rect 1104 28815 1133 28849
rect 1167 28815 1225 28849
rect 1259 28815 1317 28849
rect 1121 28665 1340 28815
rect 1121 28557 1225 28665
rect 1259 28523 1340 28631
rect 1121 28305 1340 28523
rect 1104 28271 1133 28305
rect 1167 28271 1225 28305
rect 1259 28271 1317 28305
rect 1121 28053 1340 28271
rect 1121 27911 1225 28019
rect 1259 27945 1340 28053
rect 1121 27761 1340 27911
rect 1104 27727 1133 27761
rect 1167 27727 1225 27761
rect 1259 27727 1317 27761
rect 1121 27577 1340 27727
rect 1121 27469 1225 27577
rect 1259 27435 1340 27543
rect 1121 27217 1340 27435
rect 1104 27183 1133 27217
rect 1167 27183 1225 27217
rect 1259 27183 1317 27217
rect 1121 26965 1340 27183
rect 1121 26823 1225 26931
rect 1259 26857 1340 26965
rect 1121 26673 1340 26823
rect 1104 26639 1133 26673
rect 1167 26639 1225 26673
rect 1259 26639 1317 26673
rect 1121 26489 1340 26639
rect 1121 26381 1225 26489
rect 1259 26347 1340 26455
rect 1121 26129 1340 26347
rect 1104 26095 1133 26129
rect 1167 26095 1225 26129
rect 1259 26095 1317 26129
rect 1121 25877 1340 26095
rect 1121 25735 1225 25843
rect 1259 25769 1340 25877
rect 1121 25585 1340 25735
rect 1104 25551 1133 25585
rect 1167 25551 1225 25585
rect 1259 25551 1317 25585
rect 1121 25401 1340 25551
rect 1121 25293 1225 25401
rect 1259 25259 1340 25367
rect 1121 25041 1340 25259
rect 1104 25007 1133 25041
rect 1167 25007 1225 25041
rect 1259 25007 1317 25041
rect 1121 24789 1340 25007
rect 1121 24647 1225 24755
rect 1259 24681 1340 24789
rect 1121 24497 1340 24647
rect 1104 24463 1133 24497
rect 1167 24463 1225 24497
rect 1259 24463 1317 24497
rect 1121 24313 1340 24463
rect 1121 24205 1225 24313
rect 1259 24171 1340 24279
rect 1121 23953 1340 24171
rect 1104 23919 1133 23953
rect 1167 23919 1225 23953
rect 1259 23919 1317 23953
rect 1121 23701 1340 23919
rect 1121 23559 1225 23667
rect 1259 23593 1340 23701
rect 1121 23409 1340 23559
rect 1104 23375 1133 23409
rect 1167 23375 1225 23409
rect 1259 23375 1317 23409
rect 1121 23225 1340 23375
rect 1121 23117 1225 23225
rect 1259 23083 1340 23191
rect 1121 22865 1340 23083
rect 1104 22831 1133 22865
rect 1167 22831 1225 22865
rect 1259 22831 1317 22865
rect 1121 22613 1340 22831
rect 1121 22471 1225 22579
rect 1259 22505 1340 22613
rect 1121 22321 1340 22471
rect 1104 22287 1133 22321
rect 1167 22287 1225 22321
rect 1259 22287 1317 22321
rect 1121 22137 1340 22287
rect 1121 22029 1225 22137
rect 1259 21995 1340 22103
rect 1121 21777 1340 21995
rect 1104 21743 1133 21777
rect 1167 21743 1225 21777
rect 1259 21743 1317 21777
rect 1121 21525 1340 21743
rect 1121 21383 1225 21491
rect 1259 21417 1340 21525
rect 1121 21233 1340 21383
rect 1104 21199 1133 21233
rect 1167 21199 1225 21233
rect 1259 21199 1317 21233
rect 1121 21049 1340 21199
rect 1121 20941 1225 21049
rect 1259 20907 1340 21015
rect 1121 20689 1340 20907
rect 1104 20655 1133 20689
rect 1167 20655 1225 20689
rect 1259 20655 1317 20689
rect 1121 20437 1340 20655
rect 1121 20295 1225 20403
rect 1259 20329 1340 20437
rect 1121 20145 1340 20295
rect 1104 20111 1133 20145
rect 1167 20111 1225 20145
rect 1259 20111 1317 20145
rect 1121 19961 1340 20111
rect 1121 19853 1225 19961
rect 1259 19819 1340 19927
rect 1121 19601 1340 19819
rect 1104 19567 1133 19601
rect 1167 19567 1225 19601
rect 1259 19567 1317 19601
rect 1121 19349 1340 19567
rect 1121 19207 1225 19315
rect 1259 19241 1340 19349
rect 1121 19057 1340 19207
rect 1104 19023 1133 19057
rect 1167 19023 1225 19057
rect 1259 19023 1317 19057
rect 1121 18873 1340 19023
rect 1121 18765 1225 18873
rect 1259 18731 1340 18839
rect 1121 18513 1340 18731
rect 1104 18479 1133 18513
rect 1167 18479 1225 18513
rect 1259 18479 1317 18513
rect 1121 18261 1340 18479
rect 1121 18119 1225 18227
rect 1259 18153 1340 18261
rect 1121 17969 1340 18119
rect 1104 17935 1133 17969
rect 1167 17935 1225 17969
rect 1259 17935 1317 17969
rect 1121 17785 1340 17935
rect 1121 17677 1225 17785
rect 1259 17643 1340 17751
rect 1121 17425 1340 17643
rect 1104 17391 1133 17425
rect 1167 17391 1225 17425
rect 1259 17391 1317 17425
rect 1121 17173 1340 17391
rect 1121 17031 1225 17139
rect 1259 17065 1340 17173
rect 1121 16881 1340 17031
rect 1104 16847 1133 16881
rect 1167 16847 1225 16881
rect 1259 16847 1317 16881
rect 1121 16697 1340 16847
rect 1121 16589 1225 16697
rect 1259 16555 1340 16663
rect 1121 16337 1340 16555
rect 1104 16303 1133 16337
rect 1167 16303 1225 16337
rect 1259 16303 1317 16337
rect 1121 16085 1340 16303
rect 1121 15943 1225 16051
rect 1259 15977 1340 16085
rect 1121 15793 1340 15943
rect 1104 15759 1133 15793
rect 1167 15759 1225 15793
rect 1259 15759 1317 15793
rect 1121 15609 1340 15759
rect 1121 15501 1225 15609
rect 1259 15467 1340 15575
rect 1121 15249 1340 15467
rect 1104 15215 1133 15249
rect 1167 15215 1225 15249
rect 1259 15215 1317 15249
rect 1121 14997 1340 15215
rect 1121 14855 1225 14963
rect 1259 14889 1340 14997
rect 1121 14705 1340 14855
rect 1104 14671 1133 14705
rect 1167 14671 1225 14705
rect 1259 14671 1317 14705
rect 1121 14521 1340 14671
rect 1121 14413 1225 14521
rect 1259 14379 1340 14487
rect 1121 14161 1340 14379
rect 1104 14127 1133 14161
rect 1167 14127 1225 14161
rect 1259 14127 1317 14161
rect 1121 13909 1340 14127
rect 1121 13767 1225 13875
rect 1259 13801 1340 13909
rect 1121 13617 1340 13767
rect 1104 13583 1133 13617
rect 1167 13583 1225 13617
rect 1259 13583 1317 13617
rect 1121 13433 1340 13583
rect 1121 13325 1225 13433
rect 1259 13291 1340 13399
rect 1121 13073 1340 13291
rect 1104 13039 1133 13073
rect 1167 13039 1225 13073
rect 1259 13039 1317 13073
rect 1121 12821 1340 13039
rect 1121 12679 1225 12787
rect 1259 12713 1340 12821
rect 1121 12529 1340 12679
rect 1104 12495 1133 12529
rect 1167 12495 1225 12529
rect 1259 12495 1317 12529
rect 1121 12345 1340 12495
rect 1121 12237 1225 12345
rect 1259 12203 1340 12311
rect 1121 11985 1340 12203
rect 1104 11951 1133 11985
rect 1167 11951 1225 11985
rect 1259 11951 1317 11985
rect 1121 11733 1340 11951
rect 1121 11591 1225 11699
rect 1259 11625 1340 11733
rect 1121 11441 1340 11591
rect 1104 11407 1133 11441
rect 1167 11407 1225 11441
rect 1259 11407 1317 11441
rect 1121 11257 1340 11407
rect 1121 11149 1225 11257
rect 1259 11115 1340 11223
rect 1121 10897 1340 11115
rect 1104 10863 1133 10897
rect 1167 10863 1225 10897
rect 1259 10863 1317 10897
rect 1121 10645 1340 10863
rect 1121 10503 1225 10611
rect 1259 10537 1340 10645
rect 1121 10353 1340 10503
rect 1104 10319 1133 10353
rect 1167 10319 1225 10353
rect 1259 10319 1317 10353
rect 1121 10169 1340 10319
rect 1121 10061 1225 10169
rect 1259 10027 1340 10135
rect 1121 9809 1340 10027
rect 1104 9775 1133 9809
rect 1167 9775 1225 9809
rect 1259 9775 1317 9809
rect 1121 9557 1340 9775
rect 1121 9415 1225 9523
rect 1259 9449 1340 9557
rect 1121 9265 1340 9415
rect 1104 9231 1133 9265
rect 1167 9231 1225 9265
rect 1259 9231 1317 9265
rect 1121 9081 1340 9231
rect 1121 8973 1225 9081
rect 1259 8939 1340 9047
rect 1121 8721 1340 8939
rect 1104 8687 1133 8721
rect 1167 8687 1225 8721
rect 1259 8687 1317 8721
rect 1121 8469 1340 8687
rect 1121 8327 1225 8435
rect 1259 8361 1340 8469
rect 1121 8177 1340 8327
rect 1104 8143 1133 8177
rect 1167 8143 1225 8177
rect 1259 8143 1317 8177
rect 1121 7993 1340 8143
rect 1121 7885 1225 7993
rect 1259 7851 1340 7959
rect 1121 7633 1340 7851
rect 1104 7599 1133 7633
rect 1167 7599 1225 7633
rect 1259 7599 1317 7633
rect 1121 7381 1340 7599
rect 1121 7239 1225 7347
rect 1259 7273 1340 7381
rect 1121 7089 1340 7239
rect 1104 7055 1133 7089
rect 1167 7055 1225 7089
rect 1259 7055 1317 7089
rect 1121 6905 1340 7055
rect 1121 6797 1225 6905
rect 1259 6763 1340 6871
rect 1121 6545 1340 6763
rect 1104 6511 1133 6545
rect 1167 6511 1225 6545
rect 1259 6511 1317 6545
rect 1121 6293 1340 6511
rect 1121 6151 1225 6259
rect 1259 6185 1340 6293
rect 1121 6001 1340 6151
rect 1104 5967 1133 6001
rect 1167 5967 1225 6001
rect 1259 5967 1317 6001
rect 1121 5817 1340 5967
rect 1121 5709 1225 5817
rect 1259 5675 1340 5783
rect 1121 5457 1340 5675
rect 1104 5423 1133 5457
rect 1167 5423 1225 5457
rect 1259 5423 1317 5457
rect 1121 5205 1340 5423
rect 1121 5063 1225 5171
rect 1259 5097 1340 5205
rect 1121 4913 1340 5063
rect 1104 4879 1133 4913
rect 1167 4879 1225 4913
rect 1259 4879 1317 4913
rect 1121 4729 1340 4879
rect 1121 4621 1225 4729
rect 1259 4587 1340 4695
rect 1121 4369 1340 4587
rect 1104 4335 1133 4369
rect 1167 4335 1225 4369
rect 1259 4335 1317 4369
rect 1121 4117 1340 4335
rect 1121 3975 1225 4083
rect 1259 4009 1340 4117
rect 1121 3825 1340 3975
rect 1104 3791 1133 3825
rect 1167 3791 1225 3825
rect 1259 3791 1317 3825
rect 1121 3641 1340 3791
rect 1121 3533 1225 3641
rect 1259 3499 1340 3607
rect 1121 3281 1340 3499
rect 1104 3247 1133 3281
rect 1167 3247 1225 3281
rect 1259 3247 1317 3281
rect 1121 3029 1340 3247
rect 1121 2887 1225 2995
rect 1259 2921 1340 3029
rect 1121 2737 1340 2887
rect 1104 2703 1133 2737
rect 1167 2703 1225 2737
rect 1259 2703 1317 2737
rect 1121 2553 1340 2703
rect 1121 2445 1225 2553
rect 1259 2411 1340 2519
rect 1121 2193 1340 2411
rect 1104 2159 1133 2193
rect 1167 2159 1225 2193
rect 1259 2159 1317 2193
rect 298660 297551 298661 297585
rect 298695 297551 298753 297585
rect 298787 297551 298816 297585
rect 298660 297401 298799 297551
rect 298660 297259 298661 297367
rect 298695 297293 298799 297401
rect 298660 297041 298799 297259
rect 298660 297007 298661 297041
rect 298695 297007 298753 297041
rect 298787 297007 298816 297041
rect 298660 296789 298799 297007
rect 298660 296681 298661 296789
rect 298695 296647 298799 296755
rect 298660 296497 298799 296647
rect 298660 296463 298661 296497
rect 298695 296463 298753 296497
rect 298787 296463 298816 296497
rect 298660 296313 298799 296463
rect 298660 296171 298661 296279
rect 298695 296205 298799 296313
rect 298660 295953 298799 296171
rect 298660 295919 298661 295953
rect 298695 295919 298753 295953
rect 298787 295919 298816 295953
rect 298660 295701 298799 295919
rect 298660 295593 298661 295701
rect 298695 295559 298799 295667
rect 298660 295409 298799 295559
rect 298660 295375 298661 295409
rect 298695 295375 298753 295409
rect 298787 295375 298816 295409
rect 298660 295225 298799 295375
rect 298660 295083 298661 295191
rect 298695 295117 298799 295225
rect 298660 294865 298799 295083
rect 298660 294831 298661 294865
rect 298695 294831 298753 294865
rect 298787 294831 298816 294865
rect 298660 294613 298799 294831
rect 298660 294505 298661 294613
rect 298695 294471 298799 294579
rect 298660 294321 298799 294471
rect 298660 294287 298661 294321
rect 298695 294287 298753 294321
rect 298787 294287 298816 294321
rect 298660 294137 298799 294287
rect 298660 293995 298661 294103
rect 298695 294029 298799 294137
rect 298660 293777 298799 293995
rect 298660 293743 298661 293777
rect 298695 293743 298753 293777
rect 298787 293743 298816 293777
rect 298660 293525 298799 293743
rect 298660 293417 298661 293525
rect 298695 293383 298799 293491
rect 298660 293233 298799 293383
rect 298660 293199 298661 293233
rect 298695 293199 298753 293233
rect 298787 293199 298816 293233
rect 298660 293049 298799 293199
rect 298660 292907 298661 293015
rect 298695 292941 298799 293049
rect 298660 292689 298799 292907
rect 298660 292655 298661 292689
rect 298695 292655 298753 292689
rect 298787 292655 298816 292689
rect 298660 292437 298799 292655
rect 298660 292329 298661 292437
rect 298695 292295 298799 292403
rect 298660 292145 298799 292295
rect 298660 292111 298661 292145
rect 298695 292111 298753 292145
rect 298787 292111 298816 292145
rect 298660 291961 298799 292111
rect 298660 291819 298661 291927
rect 298695 291853 298799 291961
rect 298660 291601 298799 291819
rect 298660 291567 298661 291601
rect 298695 291567 298753 291601
rect 298787 291567 298816 291601
rect 298660 291349 298799 291567
rect 298660 291241 298661 291349
rect 298695 291207 298799 291315
rect 298660 291057 298799 291207
rect 298660 291023 298661 291057
rect 298695 291023 298753 291057
rect 298787 291023 298816 291057
rect 298660 290873 298799 291023
rect 298660 290731 298661 290839
rect 298695 290765 298799 290873
rect 298660 290513 298799 290731
rect 298660 290479 298661 290513
rect 298695 290479 298753 290513
rect 298787 290479 298816 290513
rect 298660 290261 298799 290479
rect 298660 290153 298661 290261
rect 298695 290119 298799 290227
rect 298660 289969 298799 290119
rect 298660 289935 298661 289969
rect 298695 289935 298753 289969
rect 298787 289935 298816 289969
rect 298660 289785 298799 289935
rect 298660 289643 298661 289751
rect 298695 289677 298799 289785
rect 298660 289425 298799 289643
rect 298660 289391 298661 289425
rect 298695 289391 298753 289425
rect 298787 289391 298816 289425
rect 298660 289173 298799 289391
rect 298660 289065 298661 289173
rect 298695 289031 298799 289139
rect 298660 288881 298799 289031
rect 298660 288847 298661 288881
rect 298695 288847 298753 288881
rect 298787 288847 298816 288881
rect 298660 288697 298799 288847
rect 298660 288555 298661 288663
rect 298695 288589 298799 288697
rect 298660 288337 298799 288555
rect 298660 288303 298661 288337
rect 298695 288303 298753 288337
rect 298787 288303 298816 288337
rect 298660 288085 298799 288303
rect 298660 287977 298661 288085
rect 298695 287943 298799 288051
rect 298660 287793 298799 287943
rect 298660 287759 298661 287793
rect 298695 287759 298753 287793
rect 298787 287759 298816 287793
rect 298660 287609 298799 287759
rect 298660 287467 298661 287575
rect 298695 287501 298799 287609
rect 298660 287249 298799 287467
rect 298660 287215 298661 287249
rect 298695 287215 298753 287249
rect 298787 287215 298816 287249
rect 298660 286997 298799 287215
rect 298660 286889 298661 286997
rect 298695 286855 298799 286963
rect 298660 286705 298799 286855
rect 298660 286671 298661 286705
rect 298695 286671 298753 286705
rect 298787 286671 298816 286705
rect 298660 286521 298799 286671
rect 298660 286379 298661 286487
rect 298695 286413 298799 286521
rect 298660 286161 298799 286379
rect 298660 286127 298661 286161
rect 298695 286127 298753 286161
rect 298787 286127 298816 286161
rect 298660 285909 298799 286127
rect 298660 285801 298661 285909
rect 298695 285767 298799 285875
rect 298660 285617 298799 285767
rect 298660 285583 298661 285617
rect 298695 285583 298753 285617
rect 298787 285583 298816 285617
rect 298660 285433 298799 285583
rect 298660 285291 298661 285399
rect 298695 285325 298799 285433
rect 298660 285073 298799 285291
rect 298660 285039 298661 285073
rect 298695 285039 298753 285073
rect 298787 285039 298816 285073
rect 298660 284821 298799 285039
rect 298660 284713 298661 284821
rect 298695 284679 298799 284787
rect 298660 284529 298799 284679
rect 298660 284495 298661 284529
rect 298695 284495 298753 284529
rect 298787 284495 298816 284529
rect 298660 284345 298799 284495
rect 298660 284203 298661 284311
rect 298695 284237 298799 284345
rect 298660 283985 298799 284203
rect 298660 283951 298661 283985
rect 298695 283951 298753 283985
rect 298787 283951 298816 283985
rect 298660 283733 298799 283951
rect 298660 283625 298661 283733
rect 298695 283591 298799 283699
rect 298660 283441 298799 283591
rect 298660 283407 298661 283441
rect 298695 283407 298753 283441
rect 298787 283407 298816 283441
rect 298660 283257 298799 283407
rect 298660 283115 298661 283223
rect 298695 283149 298799 283257
rect 298660 282897 298799 283115
rect 298660 282863 298661 282897
rect 298695 282863 298753 282897
rect 298787 282863 298816 282897
rect 298660 282645 298799 282863
rect 298660 282537 298661 282645
rect 298695 282503 298799 282611
rect 298660 282353 298799 282503
rect 298660 282319 298661 282353
rect 298695 282319 298753 282353
rect 298787 282319 298816 282353
rect 298660 282169 298799 282319
rect 298660 282027 298661 282135
rect 298695 282061 298799 282169
rect 298660 281809 298799 282027
rect 298660 281775 298661 281809
rect 298695 281775 298753 281809
rect 298787 281775 298816 281809
rect 298660 281557 298799 281775
rect 298660 281449 298661 281557
rect 298695 281415 298799 281523
rect 298660 281265 298799 281415
rect 298660 281231 298661 281265
rect 298695 281231 298753 281265
rect 298787 281231 298816 281265
rect 298660 281081 298799 281231
rect 298660 280939 298661 281047
rect 298695 280973 298799 281081
rect 298660 280721 298799 280939
rect 298660 280687 298661 280721
rect 298695 280687 298753 280721
rect 298787 280687 298816 280721
rect 298660 280469 298799 280687
rect 298660 280361 298661 280469
rect 298695 280327 298799 280435
rect 298660 280177 298799 280327
rect 298660 280143 298661 280177
rect 298695 280143 298753 280177
rect 298787 280143 298816 280177
rect 298660 279993 298799 280143
rect 298660 279851 298661 279959
rect 298695 279885 298799 279993
rect 298660 279633 298799 279851
rect 298660 279599 298661 279633
rect 298695 279599 298753 279633
rect 298787 279599 298816 279633
rect 298660 279381 298799 279599
rect 298660 279273 298661 279381
rect 298695 279239 298799 279347
rect 298660 279089 298799 279239
rect 298660 279055 298661 279089
rect 298695 279055 298753 279089
rect 298787 279055 298816 279089
rect 298660 278905 298799 279055
rect 298660 278763 298661 278871
rect 298695 278797 298799 278905
rect 298660 278545 298799 278763
rect 298660 278511 298661 278545
rect 298695 278511 298753 278545
rect 298787 278511 298816 278545
rect 298660 278293 298799 278511
rect 298660 278185 298661 278293
rect 298695 278151 298799 278259
rect 298660 278001 298799 278151
rect 298660 277967 298661 278001
rect 298695 277967 298753 278001
rect 298787 277967 298816 278001
rect 298660 277817 298799 277967
rect 298660 277675 298661 277783
rect 298695 277709 298799 277817
rect 298660 277457 298799 277675
rect 298660 277423 298661 277457
rect 298695 277423 298753 277457
rect 298787 277423 298816 277457
rect 298660 277205 298799 277423
rect 298660 277097 298661 277205
rect 298695 277063 298799 277171
rect 298660 276913 298799 277063
rect 298660 276879 298661 276913
rect 298695 276879 298753 276913
rect 298787 276879 298816 276913
rect 298660 276729 298799 276879
rect 298660 276587 298661 276695
rect 298695 276621 298799 276729
rect 298660 276369 298799 276587
rect 298660 276335 298661 276369
rect 298695 276335 298753 276369
rect 298787 276335 298816 276369
rect 298660 276117 298799 276335
rect 298660 276009 298661 276117
rect 298695 275975 298799 276083
rect 298660 275825 298799 275975
rect 298660 275791 298661 275825
rect 298695 275791 298753 275825
rect 298787 275791 298816 275825
rect 298660 275641 298799 275791
rect 298660 275499 298661 275607
rect 298695 275533 298799 275641
rect 298660 275281 298799 275499
rect 298660 275247 298661 275281
rect 298695 275247 298753 275281
rect 298787 275247 298816 275281
rect 298660 275029 298799 275247
rect 298660 274921 298661 275029
rect 298695 274887 298799 274995
rect 298660 274737 298799 274887
rect 298660 274703 298661 274737
rect 298695 274703 298753 274737
rect 298787 274703 298816 274737
rect 298660 274553 298799 274703
rect 298660 274411 298661 274519
rect 298695 274445 298799 274553
rect 298660 274193 298799 274411
rect 298660 274159 298661 274193
rect 298695 274159 298753 274193
rect 298787 274159 298816 274193
rect 298660 273941 298799 274159
rect 298660 273833 298661 273941
rect 298695 273799 298799 273907
rect 298660 273649 298799 273799
rect 298660 273615 298661 273649
rect 298695 273615 298753 273649
rect 298787 273615 298816 273649
rect 298660 273465 298799 273615
rect 298660 273323 298661 273431
rect 298695 273357 298799 273465
rect 298660 273105 298799 273323
rect 298660 273071 298661 273105
rect 298695 273071 298753 273105
rect 298787 273071 298816 273105
rect 298660 272853 298799 273071
rect 298660 272745 298661 272853
rect 298695 272711 298799 272819
rect 298660 272561 298799 272711
rect 298660 272527 298661 272561
rect 298695 272527 298753 272561
rect 298787 272527 298816 272561
rect 298660 272377 298799 272527
rect 298660 272235 298661 272343
rect 298695 272269 298799 272377
rect 298660 272017 298799 272235
rect 298660 271983 298661 272017
rect 298695 271983 298753 272017
rect 298787 271983 298816 272017
rect 298660 271765 298799 271983
rect 298660 271657 298661 271765
rect 298695 271623 298799 271731
rect 298660 271473 298799 271623
rect 298660 271439 298661 271473
rect 298695 271439 298753 271473
rect 298787 271439 298816 271473
rect 298660 271289 298799 271439
rect 298660 271147 298661 271255
rect 298695 271181 298799 271289
rect 298660 270929 298799 271147
rect 298660 270895 298661 270929
rect 298695 270895 298753 270929
rect 298787 270895 298816 270929
rect 298660 270677 298799 270895
rect 298660 270569 298661 270677
rect 298695 270535 298799 270643
rect 298660 270385 298799 270535
rect 298660 270351 298661 270385
rect 298695 270351 298753 270385
rect 298787 270351 298816 270385
rect 298660 270201 298799 270351
rect 298660 270059 298661 270167
rect 298695 270093 298799 270201
rect 298660 269841 298799 270059
rect 298660 269807 298661 269841
rect 298695 269807 298753 269841
rect 298787 269807 298816 269841
rect 298660 269589 298799 269807
rect 298660 269481 298661 269589
rect 298695 269447 298799 269555
rect 298660 269297 298799 269447
rect 298660 269263 298661 269297
rect 298695 269263 298753 269297
rect 298787 269263 298816 269297
rect 298660 269113 298799 269263
rect 298660 268971 298661 269079
rect 298695 269005 298799 269113
rect 298660 268753 298799 268971
rect 298660 268719 298661 268753
rect 298695 268719 298753 268753
rect 298787 268719 298816 268753
rect 298660 268501 298799 268719
rect 298660 268393 298661 268501
rect 298695 268359 298799 268467
rect 298660 268209 298799 268359
rect 298660 268175 298661 268209
rect 298695 268175 298753 268209
rect 298787 268175 298816 268209
rect 298660 268025 298799 268175
rect 298660 267883 298661 267991
rect 298695 267917 298799 268025
rect 298660 267665 298799 267883
rect 298660 267631 298661 267665
rect 298695 267631 298753 267665
rect 298787 267631 298816 267665
rect 298660 267413 298799 267631
rect 298660 267305 298661 267413
rect 298695 267271 298799 267379
rect 298660 267121 298799 267271
rect 298660 267087 298661 267121
rect 298695 267087 298753 267121
rect 298787 267087 298816 267121
rect 298660 266937 298799 267087
rect 298660 266795 298661 266903
rect 298695 266829 298799 266937
rect 298660 266577 298799 266795
rect 298660 266543 298661 266577
rect 298695 266543 298753 266577
rect 298787 266543 298816 266577
rect 298660 266325 298799 266543
rect 298660 266217 298661 266325
rect 298695 266183 298799 266291
rect 298660 266033 298799 266183
rect 298660 265999 298661 266033
rect 298695 265999 298753 266033
rect 298787 265999 298816 266033
rect 298660 265849 298799 265999
rect 298660 265707 298661 265815
rect 298695 265741 298799 265849
rect 298660 265489 298799 265707
rect 298660 265455 298661 265489
rect 298695 265455 298753 265489
rect 298787 265455 298816 265489
rect 298660 265237 298799 265455
rect 298660 265129 298661 265237
rect 298695 265095 298799 265203
rect 298660 264945 298799 265095
rect 298660 264911 298661 264945
rect 298695 264911 298753 264945
rect 298787 264911 298816 264945
rect 298660 264761 298799 264911
rect 298660 264619 298661 264727
rect 298695 264653 298799 264761
rect 298660 264401 298799 264619
rect 298660 264367 298661 264401
rect 298695 264367 298753 264401
rect 298787 264367 298816 264401
rect 298660 264149 298799 264367
rect 298660 264041 298661 264149
rect 298695 264007 298799 264115
rect 298660 263857 298799 264007
rect 298660 263823 298661 263857
rect 298695 263823 298753 263857
rect 298787 263823 298816 263857
rect 298660 263673 298799 263823
rect 298660 263531 298661 263639
rect 298695 263565 298799 263673
rect 298660 263313 298799 263531
rect 298660 263279 298661 263313
rect 298695 263279 298753 263313
rect 298787 263279 298816 263313
rect 298660 263061 298799 263279
rect 298660 262953 298661 263061
rect 298695 262919 298799 263027
rect 298660 262769 298799 262919
rect 298660 262735 298661 262769
rect 298695 262735 298753 262769
rect 298787 262735 298816 262769
rect 298660 262585 298799 262735
rect 298660 262443 298661 262551
rect 298695 262477 298799 262585
rect 298660 262225 298799 262443
rect 298660 262191 298661 262225
rect 298695 262191 298753 262225
rect 298787 262191 298816 262225
rect 298660 261973 298799 262191
rect 298660 261865 298661 261973
rect 298695 261831 298799 261939
rect 298660 261681 298799 261831
rect 298660 261647 298661 261681
rect 298695 261647 298753 261681
rect 298787 261647 298816 261681
rect 298660 261497 298799 261647
rect 298660 261355 298661 261463
rect 298695 261389 298799 261497
rect 298660 261137 298799 261355
rect 298660 261103 298661 261137
rect 298695 261103 298753 261137
rect 298787 261103 298816 261137
rect 298660 260885 298799 261103
rect 298660 260777 298661 260885
rect 298695 260743 298799 260851
rect 298660 260593 298799 260743
rect 298660 260559 298661 260593
rect 298695 260559 298753 260593
rect 298787 260559 298816 260593
rect 298660 260409 298799 260559
rect 298660 260267 298661 260375
rect 298695 260301 298799 260409
rect 298660 260049 298799 260267
rect 298660 260015 298661 260049
rect 298695 260015 298753 260049
rect 298787 260015 298816 260049
rect 298660 259797 298799 260015
rect 298660 259689 298661 259797
rect 298695 259655 298799 259763
rect 298660 259505 298799 259655
rect 298660 259471 298661 259505
rect 298695 259471 298753 259505
rect 298787 259471 298816 259505
rect 298660 259321 298799 259471
rect 298660 259179 298661 259287
rect 298695 259213 298799 259321
rect 298660 258961 298799 259179
rect 298660 258927 298661 258961
rect 298695 258927 298753 258961
rect 298787 258927 298816 258961
rect 298660 258709 298799 258927
rect 298660 258601 298661 258709
rect 298695 258567 298799 258675
rect 298660 258417 298799 258567
rect 298660 258383 298661 258417
rect 298695 258383 298753 258417
rect 298787 258383 298816 258417
rect 298660 258233 298799 258383
rect 298660 258091 298661 258199
rect 298695 258125 298799 258233
rect 298660 257873 298799 258091
rect 298660 257839 298661 257873
rect 298695 257839 298753 257873
rect 298787 257839 298816 257873
rect 298660 257621 298799 257839
rect 298660 257513 298661 257621
rect 298695 257479 298799 257587
rect 298660 257329 298799 257479
rect 298660 257295 298661 257329
rect 298695 257295 298753 257329
rect 298787 257295 298816 257329
rect 298660 257145 298799 257295
rect 298660 257003 298661 257111
rect 298695 257037 298799 257145
rect 298660 256785 298799 257003
rect 298660 256751 298661 256785
rect 298695 256751 298753 256785
rect 298787 256751 298816 256785
rect 298660 256533 298799 256751
rect 298660 256425 298661 256533
rect 298695 256391 298799 256499
rect 298660 256241 298799 256391
rect 298660 256207 298661 256241
rect 298695 256207 298753 256241
rect 298787 256207 298816 256241
rect 298660 256057 298799 256207
rect 298660 255915 298661 256023
rect 298695 255949 298799 256057
rect 298660 255697 298799 255915
rect 298660 255663 298661 255697
rect 298695 255663 298753 255697
rect 298787 255663 298816 255697
rect 298660 255445 298799 255663
rect 298660 255337 298661 255445
rect 298695 255303 298799 255411
rect 298660 255153 298799 255303
rect 298660 255119 298661 255153
rect 298695 255119 298753 255153
rect 298787 255119 298816 255153
rect 298660 254969 298799 255119
rect 298660 254827 298661 254935
rect 298695 254861 298799 254969
rect 298660 254609 298799 254827
rect 298660 254575 298661 254609
rect 298695 254575 298753 254609
rect 298787 254575 298816 254609
rect 298660 254357 298799 254575
rect 298660 254249 298661 254357
rect 298695 254215 298799 254323
rect 298660 254065 298799 254215
rect 298660 254031 298661 254065
rect 298695 254031 298753 254065
rect 298787 254031 298816 254065
rect 298660 253881 298799 254031
rect 298660 253739 298661 253847
rect 298695 253773 298799 253881
rect 298660 253521 298799 253739
rect 298660 253487 298661 253521
rect 298695 253487 298753 253521
rect 298787 253487 298816 253521
rect 298660 253269 298799 253487
rect 298660 253161 298661 253269
rect 298695 253127 298799 253235
rect 298660 252977 298799 253127
rect 298660 252943 298661 252977
rect 298695 252943 298753 252977
rect 298787 252943 298816 252977
rect 298660 252793 298799 252943
rect 298660 252651 298661 252759
rect 298695 252685 298799 252793
rect 298660 252433 298799 252651
rect 298660 252399 298661 252433
rect 298695 252399 298753 252433
rect 298787 252399 298816 252433
rect 298660 252181 298799 252399
rect 298660 252073 298661 252181
rect 298695 252039 298799 252147
rect 298660 251889 298799 252039
rect 298660 251855 298661 251889
rect 298695 251855 298753 251889
rect 298787 251855 298816 251889
rect 298660 251705 298799 251855
rect 298660 251563 298661 251671
rect 298695 251597 298799 251705
rect 298660 251345 298799 251563
rect 298660 251311 298661 251345
rect 298695 251311 298753 251345
rect 298787 251311 298816 251345
rect 298660 251093 298799 251311
rect 298660 250985 298661 251093
rect 298695 250951 298799 251059
rect 298660 250801 298799 250951
rect 298660 250767 298661 250801
rect 298695 250767 298753 250801
rect 298787 250767 298816 250801
rect 298660 250617 298799 250767
rect 298660 250475 298661 250583
rect 298695 250509 298799 250617
rect 298660 250257 298799 250475
rect 298660 250223 298661 250257
rect 298695 250223 298753 250257
rect 298787 250223 298816 250257
rect 298660 250005 298799 250223
rect 298660 249897 298661 250005
rect 298695 249863 298799 249971
rect 298660 249713 298799 249863
rect 298660 249679 298661 249713
rect 298695 249679 298753 249713
rect 298787 249679 298816 249713
rect 298660 249529 298799 249679
rect 298660 249387 298661 249495
rect 298695 249421 298799 249529
rect 298660 249169 298799 249387
rect 298660 249135 298661 249169
rect 298695 249135 298753 249169
rect 298787 249135 298816 249169
rect 298660 248917 298799 249135
rect 298660 248809 298661 248917
rect 298695 248775 298799 248883
rect 298660 248625 298799 248775
rect 298660 248591 298661 248625
rect 298695 248591 298753 248625
rect 298787 248591 298816 248625
rect 298660 248441 298799 248591
rect 298660 248299 298661 248407
rect 298695 248333 298799 248441
rect 298660 248081 298799 248299
rect 298660 248047 298661 248081
rect 298695 248047 298753 248081
rect 298787 248047 298816 248081
rect 298660 247829 298799 248047
rect 298660 247721 298661 247829
rect 298695 247687 298799 247795
rect 298660 247537 298799 247687
rect 298660 247503 298661 247537
rect 298695 247503 298753 247537
rect 298787 247503 298816 247537
rect 298660 247353 298799 247503
rect 298660 247211 298661 247319
rect 298695 247245 298799 247353
rect 298660 246993 298799 247211
rect 298660 246959 298661 246993
rect 298695 246959 298753 246993
rect 298787 246959 298816 246993
rect 298660 246741 298799 246959
rect 298660 246633 298661 246741
rect 298695 246599 298799 246707
rect 298660 246449 298799 246599
rect 298660 246415 298661 246449
rect 298695 246415 298753 246449
rect 298787 246415 298816 246449
rect 298660 246265 298799 246415
rect 298660 246123 298661 246231
rect 298695 246157 298799 246265
rect 298660 245905 298799 246123
rect 298660 245871 298661 245905
rect 298695 245871 298753 245905
rect 298787 245871 298816 245905
rect 298660 245653 298799 245871
rect 298660 245545 298661 245653
rect 298695 245511 298799 245619
rect 298660 245361 298799 245511
rect 298660 245327 298661 245361
rect 298695 245327 298753 245361
rect 298787 245327 298816 245361
rect 298660 245177 298799 245327
rect 298660 245035 298661 245143
rect 298695 245069 298799 245177
rect 298660 244817 298799 245035
rect 298660 244783 298661 244817
rect 298695 244783 298753 244817
rect 298787 244783 298816 244817
rect 298660 244565 298799 244783
rect 298660 244457 298661 244565
rect 298695 244423 298799 244531
rect 298660 244273 298799 244423
rect 298660 244239 298661 244273
rect 298695 244239 298753 244273
rect 298787 244239 298816 244273
rect 298660 244089 298799 244239
rect 298660 243947 298661 244055
rect 298695 243981 298799 244089
rect 298660 243729 298799 243947
rect 298660 243695 298661 243729
rect 298695 243695 298753 243729
rect 298787 243695 298816 243729
rect 298660 243477 298799 243695
rect 298660 243369 298661 243477
rect 298695 243335 298799 243443
rect 298660 243185 298799 243335
rect 298660 243151 298661 243185
rect 298695 243151 298753 243185
rect 298787 243151 298816 243185
rect 298660 243001 298799 243151
rect 298660 242859 298661 242967
rect 298695 242893 298799 243001
rect 298660 242641 298799 242859
rect 298660 242607 298661 242641
rect 298695 242607 298753 242641
rect 298787 242607 298816 242641
rect 298660 242389 298799 242607
rect 298660 242281 298661 242389
rect 298695 242247 298799 242355
rect 298660 242097 298799 242247
rect 298660 242063 298661 242097
rect 298695 242063 298753 242097
rect 298787 242063 298816 242097
rect 298660 241913 298799 242063
rect 298660 241771 298661 241879
rect 298695 241805 298799 241913
rect 298660 241553 298799 241771
rect 298660 241519 298661 241553
rect 298695 241519 298753 241553
rect 298787 241519 298816 241553
rect 298660 241301 298799 241519
rect 298660 241193 298661 241301
rect 298695 241159 298799 241267
rect 298660 241009 298799 241159
rect 298660 240975 298661 241009
rect 298695 240975 298753 241009
rect 298787 240975 298816 241009
rect 298660 240825 298799 240975
rect 298660 240683 298661 240791
rect 298695 240717 298799 240825
rect 298660 240465 298799 240683
rect 298660 240431 298661 240465
rect 298695 240431 298753 240465
rect 298787 240431 298816 240465
rect 298660 240213 298799 240431
rect 298660 240105 298661 240213
rect 298695 240071 298799 240179
rect 298660 239921 298799 240071
rect 298660 239887 298661 239921
rect 298695 239887 298753 239921
rect 298787 239887 298816 239921
rect 298660 239737 298799 239887
rect 298660 239595 298661 239703
rect 298695 239629 298799 239737
rect 298660 239377 298799 239595
rect 298660 239343 298661 239377
rect 298695 239343 298753 239377
rect 298787 239343 298816 239377
rect 298660 239125 298799 239343
rect 298660 239017 298661 239125
rect 298695 238983 298799 239091
rect 298660 238833 298799 238983
rect 298660 238799 298661 238833
rect 298695 238799 298753 238833
rect 298787 238799 298816 238833
rect 298660 238649 298799 238799
rect 298660 238507 298661 238615
rect 298695 238541 298799 238649
rect 298660 238289 298799 238507
rect 298660 238255 298661 238289
rect 298695 238255 298753 238289
rect 298787 238255 298816 238289
rect 298660 238037 298799 238255
rect 298660 237929 298661 238037
rect 298695 237895 298799 238003
rect 298660 237745 298799 237895
rect 298660 237711 298661 237745
rect 298695 237711 298753 237745
rect 298787 237711 298816 237745
rect 298660 237561 298799 237711
rect 298660 237419 298661 237527
rect 298695 237453 298799 237561
rect 298660 237201 298799 237419
rect 298660 237167 298661 237201
rect 298695 237167 298753 237201
rect 298787 237167 298816 237201
rect 298660 236949 298799 237167
rect 298660 236841 298661 236949
rect 298695 236807 298799 236915
rect 298660 236657 298799 236807
rect 298660 236623 298661 236657
rect 298695 236623 298753 236657
rect 298787 236623 298816 236657
rect 298660 236473 298799 236623
rect 298660 236331 298661 236439
rect 298695 236365 298799 236473
rect 298660 236113 298799 236331
rect 298660 236079 298661 236113
rect 298695 236079 298753 236113
rect 298787 236079 298816 236113
rect 298660 235861 298799 236079
rect 298660 235753 298661 235861
rect 298695 235719 298799 235827
rect 298660 235569 298799 235719
rect 298660 235535 298661 235569
rect 298695 235535 298753 235569
rect 298787 235535 298816 235569
rect 298660 235385 298799 235535
rect 298660 235243 298661 235351
rect 298695 235277 298799 235385
rect 298660 235025 298799 235243
rect 298660 234991 298661 235025
rect 298695 234991 298753 235025
rect 298787 234991 298816 235025
rect 298660 234773 298799 234991
rect 298660 234665 298661 234773
rect 298695 234631 298799 234739
rect 298660 234481 298799 234631
rect 298660 234447 298661 234481
rect 298695 234447 298753 234481
rect 298787 234447 298816 234481
rect 298660 234297 298799 234447
rect 298660 234155 298661 234263
rect 298695 234189 298799 234297
rect 298660 233937 298799 234155
rect 298660 233903 298661 233937
rect 298695 233903 298753 233937
rect 298787 233903 298816 233937
rect 298660 233685 298799 233903
rect 298660 233577 298661 233685
rect 298695 233543 298799 233651
rect 298660 233393 298799 233543
rect 298660 233359 298661 233393
rect 298695 233359 298753 233393
rect 298787 233359 298816 233393
rect 298660 233209 298799 233359
rect 298660 233067 298661 233175
rect 298695 233101 298799 233209
rect 298660 232849 298799 233067
rect 298660 232815 298661 232849
rect 298695 232815 298753 232849
rect 298787 232815 298816 232849
rect 298660 232597 298799 232815
rect 298660 232489 298661 232597
rect 298695 232455 298799 232563
rect 298660 232305 298799 232455
rect 298660 232271 298661 232305
rect 298695 232271 298753 232305
rect 298787 232271 298816 232305
rect 298660 232121 298799 232271
rect 298660 231979 298661 232087
rect 298695 232013 298799 232121
rect 298660 231761 298799 231979
rect 298660 231727 298661 231761
rect 298695 231727 298753 231761
rect 298787 231727 298816 231761
rect 298660 231509 298799 231727
rect 298660 231401 298661 231509
rect 298695 231367 298799 231475
rect 298660 231217 298799 231367
rect 298660 231183 298661 231217
rect 298695 231183 298753 231217
rect 298787 231183 298816 231217
rect 298660 231033 298799 231183
rect 298660 230891 298661 230999
rect 298695 230925 298799 231033
rect 298660 230673 298799 230891
rect 298660 230639 298661 230673
rect 298695 230639 298753 230673
rect 298787 230639 298816 230673
rect 298660 230421 298799 230639
rect 298660 230313 298661 230421
rect 298695 230279 298799 230387
rect 298660 230129 298799 230279
rect 298660 230095 298661 230129
rect 298695 230095 298753 230129
rect 298787 230095 298816 230129
rect 298660 229945 298799 230095
rect 298660 229803 298661 229911
rect 298695 229837 298799 229945
rect 298660 229585 298799 229803
rect 298660 229551 298661 229585
rect 298695 229551 298753 229585
rect 298787 229551 298816 229585
rect 298660 229333 298799 229551
rect 298660 229225 298661 229333
rect 298695 229191 298799 229299
rect 298660 229041 298799 229191
rect 298660 229007 298661 229041
rect 298695 229007 298753 229041
rect 298787 229007 298816 229041
rect 298660 228857 298799 229007
rect 298660 228715 298661 228823
rect 298695 228749 298799 228857
rect 298660 228497 298799 228715
rect 298660 228463 298661 228497
rect 298695 228463 298753 228497
rect 298787 228463 298816 228497
rect 298660 228245 298799 228463
rect 298660 228137 298661 228245
rect 298695 228103 298799 228211
rect 298660 227953 298799 228103
rect 298660 227919 298661 227953
rect 298695 227919 298753 227953
rect 298787 227919 298816 227953
rect 298660 227769 298799 227919
rect 298660 227627 298661 227735
rect 298695 227661 298799 227769
rect 298660 227409 298799 227627
rect 298660 227375 298661 227409
rect 298695 227375 298753 227409
rect 298787 227375 298816 227409
rect 298660 227157 298799 227375
rect 298660 227049 298661 227157
rect 298695 227015 298799 227123
rect 298660 226865 298799 227015
rect 298660 226831 298661 226865
rect 298695 226831 298753 226865
rect 298787 226831 298816 226865
rect 298660 226681 298799 226831
rect 298660 226539 298661 226647
rect 298695 226573 298799 226681
rect 298660 226321 298799 226539
rect 298660 226287 298661 226321
rect 298695 226287 298753 226321
rect 298787 226287 298816 226321
rect 298660 226069 298799 226287
rect 298660 225961 298661 226069
rect 298695 225927 298799 226035
rect 298660 225777 298799 225927
rect 298660 225743 298661 225777
rect 298695 225743 298753 225777
rect 298787 225743 298816 225777
rect 298660 225593 298799 225743
rect 298660 225451 298661 225559
rect 298695 225485 298799 225593
rect 298660 225233 298799 225451
rect 298660 225199 298661 225233
rect 298695 225199 298753 225233
rect 298787 225199 298816 225233
rect 298660 224981 298799 225199
rect 298660 224873 298661 224981
rect 298695 224839 298799 224947
rect 298660 224689 298799 224839
rect 298660 224655 298661 224689
rect 298695 224655 298753 224689
rect 298787 224655 298816 224689
rect 298660 224505 298799 224655
rect 298660 224363 298661 224471
rect 298695 224397 298799 224505
rect 298660 224145 298799 224363
rect 298660 224111 298661 224145
rect 298695 224111 298753 224145
rect 298787 224111 298816 224145
rect 298660 223893 298799 224111
rect 298660 223785 298661 223893
rect 298695 223751 298799 223859
rect 298660 223601 298799 223751
rect 298660 223567 298661 223601
rect 298695 223567 298753 223601
rect 298787 223567 298816 223601
rect 298660 223417 298799 223567
rect 298660 223275 298661 223383
rect 298695 223309 298799 223417
rect 298660 223057 298799 223275
rect 298660 223023 298661 223057
rect 298695 223023 298753 223057
rect 298787 223023 298816 223057
rect 298660 222805 298799 223023
rect 298660 222697 298661 222805
rect 298695 222663 298799 222771
rect 298660 222513 298799 222663
rect 298660 222479 298661 222513
rect 298695 222479 298753 222513
rect 298787 222479 298816 222513
rect 298660 222329 298799 222479
rect 298660 222187 298661 222295
rect 298695 222221 298799 222329
rect 298660 221969 298799 222187
rect 298660 221935 298661 221969
rect 298695 221935 298753 221969
rect 298787 221935 298816 221969
rect 298660 221717 298799 221935
rect 298660 221609 298661 221717
rect 298695 221575 298799 221683
rect 298660 221425 298799 221575
rect 298660 221391 298661 221425
rect 298695 221391 298753 221425
rect 298787 221391 298816 221425
rect 298660 221241 298799 221391
rect 298660 221099 298661 221207
rect 298695 221133 298799 221241
rect 298660 220881 298799 221099
rect 298660 220847 298661 220881
rect 298695 220847 298753 220881
rect 298787 220847 298816 220881
rect 298660 220629 298799 220847
rect 298660 220521 298661 220629
rect 298695 220487 298799 220595
rect 298660 220337 298799 220487
rect 298660 220303 298661 220337
rect 298695 220303 298753 220337
rect 298787 220303 298816 220337
rect 298660 220153 298799 220303
rect 298660 220011 298661 220119
rect 298695 220045 298799 220153
rect 298660 219793 298799 220011
rect 298660 219759 298661 219793
rect 298695 219759 298753 219793
rect 298787 219759 298816 219793
rect 298660 219541 298799 219759
rect 298660 219433 298661 219541
rect 298695 219399 298799 219507
rect 298660 219249 298799 219399
rect 298660 219215 298661 219249
rect 298695 219215 298753 219249
rect 298787 219215 298816 219249
rect 298660 219065 298799 219215
rect 298660 218923 298661 219031
rect 298695 218957 298799 219065
rect 298660 218705 298799 218923
rect 298660 218671 298661 218705
rect 298695 218671 298753 218705
rect 298787 218671 298816 218705
rect 298660 218453 298799 218671
rect 298660 218345 298661 218453
rect 298695 218311 298799 218419
rect 298660 218161 298799 218311
rect 298660 218127 298661 218161
rect 298695 218127 298753 218161
rect 298787 218127 298816 218161
rect 298660 217977 298799 218127
rect 298660 217835 298661 217943
rect 298695 217869 298799 217977
rect 298660 217617 298799 217835
rect 298660 217583 298661 217617
rect 298695 217583 298753 217617
rect 298787 217583 298816 217617
rect 298660 217365 298799 217583
rect 298660 217257 298661 217365
rect 298695 217223 298799 217331
rect 298660 217073 298799 217223
rect 298660 217039 298661 217073
rect 298695 217039 298753 217073
rect 298787 217039 298816 217073
rect 298660 216889 298799 217039
rect 298660 216747 298661 216855
rect 298695 216781 298799 216889
rect 298660 216529 298799 216747
rect 298660 216495 298661 216529
rect 298695 216495 298753 216529
rect 298787 216495 298816 216529
rect 298660 216277 298799 216495
rect 298660 216169 298661 216277
rect 298695 216135 298799 216243
rect 298660 215985 298799 216135
rect 298660 215951 298661 215985
rect 298695 215951 298753 215985
rect 298787 215951 298816 215985
rect 298660 215801 298799 215951
rect 298660 215659 298661 215767
rect 298695 215693 298799 215801
rect 298660 215441 298799 215659
rect 298660 215407 298661 215441
rect 298695 215407 298753 215441
rect 298787 215407 298816 215441
rect 298660 215189 298799 215407
rect 298660 215081 298661 215189
rect 298695 215047 298799 215155
rect 298660 214897 298799 215047
rect 298660 214863 298661 214897
rect 298695 214863 298753 214897
rect 298787 214863 298816 214897
rect 298660 214713 298799 214863
rect 298660 214571 298661 214679
rect 298695 214605 298799 214713
rect 298660 214353 298799 214571
rect 298660 214319 298661 214353
rect 298695 214319 298753 214353
rect 298787 214319 298816 214353
rect 298660 214101 298799 214319
rect 298660 213993 298661 214101
rect 298695 213959 298799 214067
rect 298660 213809 298799 213959
rect 298660 213775 298661 213809
rect 298695 213775 298753 213809
rect 298787 213775 298816 213809
rect 298660 213625 298799 213775
rect 298660 213483 298661 213591
rect 298695 213517 298799 213625
rect 298660 213265 298799 213483
rect 298660 213231 298661 213265
rect 298695 213231 298753 213265
rect 298787 213231 298816 213265
rect 298660 213013 298799 213231
rect 298660 212905 298661 213013
rect 298695 212871 298799 212979
rect 298660 212721 298799 212871
rect 298660 212687 298661 212721
rect 298695 212687 298753 212721
rect 298787 212687 298816 212721
rect 298660 212537 298799 212687
rect 298660 212395 298661 212503
rect 298695 212429 298799 212537
rect 298660 212177 298799 212395
rect 298660 212143 298661 212177
rect 298695 212143 298753 212177
rect 298787 212143 298816 212177
rect 298660 211925 298799 212143
rect 298660 211817 298661 211925
rect 298695 211783 298799 211891
rect 298660 211633 298799 211783
rect 298660 211599 298661 211633
rect 298695 211599 298753 211633
rect 298787 211599 298816 211633
rect 298660 211449 298799 211599
rect 298660 211307 298661 211415
rect 298695 211341 298799 211449
rect 298660 211089 298799 211307
rect 298660 211055 298661 211089
rect 298695 211055 298753 211089
rect 298787 211055 298816 211089
rect 298660 210837 298799 211055
rect 298660 210729 298661 210837
rect 298695 210695 298799 210803
rect 298660 210545 298799 210695
rect 298660 210511 298661 210545
rect 298695 210511 298753 210545
rect 298787 210511 298816 210545
rect 298660 210361 298799 210511
rect 298660 210219 298661 210327
rect 298695 210253 298799 210361
rect 298660 210001 298799 210219
rect 298660 209967 298661 210001
rect 298695 209967 298753 210001
rect 298787 209967 298816 210001
rect 298660 209749 298799 209967
rect 298660 209641 298661 209749
rect 298695 209607 298799 209715
rect 298660 209457 298799 209607
rect 298660 209423 298661 209457
rect 298695 209423 298753 209457
rect 298787 209423 298816 209457
rect 298660 209273 298799 209423
rect 298660 209131 298661 209239
rect 298695 209165 298799 209273
rect 298660 208913 298799 209131
rect 298660 208879 298661 208913
rect 298695 208879 298753 208913
rect 298787 208879 298816 208913
rect 298660 208661 298799 208879
rect 298660 208553 298661 208661
rect 298695 208519 298799 208627
rect 298660 208369 298799 208519
rect 298660 208335 298661 208369
rect 298695 208335 298753 208369
rect 298787 208335 298816 208369
rect 298660 208185 298799 208335
rect 298660 208043 298661 208151
rect 298695 208077 298799 208185
rect 298660 207825 298799 208043
rect 298660 207791 298661 207825
rect 298695 207791 298753 207825
rect 298787 207791 298816 207825
rect 298660 207573 298799 207791
rect 298660 207465 298661 207573
rect 298695 207431 298799 207539
rect 298660 207281 298799 207431
rect 298660 207247 298661 207281
rect 298695 207247 298753 207281
rect 298787 207247 298816 207281
rect 298660 207097 298799 207247
rect 298660 206955 298661 207063
rect 298695 206989 298799 207097
rect 298660 206737 298799 206955
rect 298660 206703 298661 206737
rect 298695 206703 298753 206737
rect 298787 206703 298816 206737
rect 298660 206485 298799 206703
rect 298660 206377 298661 206485
rect 298695 206343 298799 206451
rect 298660 206193 298799 206343
rect 298660 206159 298661 206193
rect 298695 206159 298753 206193
rect 298787 206159 298816 206193
rect 298660 206009 298799 206159
rect 298660 205867 298661 205975
rect 298695 205901 298799 206009
rect 298660 205649 298799 205867
rect 298660 205615 298661 205649
rect 298695 205615 298753 205649
rect 298787 205615 298816 205649
rect 298660 205397 298799 205615
rect 298660 205289 298661 205397
rect 298695 205255 298799 205363
rect 298660 205105 298799 205255
rect 298660 205071 298661 205105
rect 298695 205071 298753 205105
rect 298787 205071 298816 205105
rect 298660 204921 298799 205071
rect 298660 204779 298661 204887
rect 298695 204813 298799 204921
rect 298660 204561 298799 204779
rect 298660 204527 298661 204561
rect 298695 204527 298753 204561
rect 298787 204527 298816 204561
rect 298660 204309 298799 204527
rect 298660 204201 298661 204309
rect 298695 204167 298799 204275
rect 298660 204017 298799 204167
rect 298660 203983 298661 204017
rect 298695 203983 298753 204017
rect 298787 203983 298816 204017
rect 298660 203833 298799 203983
rect 298660 203691 298661 203799
rect 298695 203725 298799 203833
rect 298660 203473 298799 203691
rect 298660 203439 298661 203473
rect 298695 203439 298753 203473
rect 298787 203439 298816 203473
rect 298660 203221 298799 203439
rect 298660 203113 298661 203221
rect 298695 203079 298799 203187
rect 298660 202929 298799 203079
rect 298660 202895 298661 202929
rect 298695 202895 298753 202929
rect 298787 202895 298816 202929
rect 298660 202745 298799 202895
rect 298660 202603 298661 202711
rect 298695 202637 298799 202745
rect 298660 202385 298799 202603
rect 298660 202351 298661 202385
rect 298695 202351 298753 202385
rect 298787 202351 298816 202385
rect 298660 202133 298799 202351
rect 298660 202025 298661 202133
rect 298695 201991 298799 202099
rect 298660 201841 298799 201991
rect 298660 201807 298661 201841
rect 298695 201807 298753 201841
rect 298787 201807 298816 201841
rect 298660 201657 298799 201807
rect 298660 201515 298661 201623
rect 298695 201549 298799 201657
rect 298660 201297 298799 201515
rect 298660 201263 298661 201297
rect 298695 201263 298753 201297
rect 298787 201263 298816 201297
rect 298660 201045 298799 201263
rect 298660 200937 298661 201045
rect 298695 200903 298799 201011
rect 298660 200753 298799 200903
rect 298660 200719 298661 200753
rect 298695 200719 298753 200753
rect 298787 200719 298816 200753
rect 298660 200569 298799 200719
rect 298660 200427 298661 200535
rect 298695 200461 298799 200569
rect 298660 200209 298799 200427
rect 298660 200175 298661 200209
rect 298695 200175 298753 200209
rect 298787 200175 298816 200209
rect 298660 199957 298799 200175
rect 298660 199849 298661 199957
rect 298695 199815 298799 199923
rect 298660 199665 298799 199815
rect 298660 199631 298661 199665
rect 298695 199631 298753 199665
rect 298787 199631 298816 199665
rect 298660 199481 298799 199631
rect 298660 199339 298661 199447
rect 298695 199373 298799 199481
rect 298660 199121 298799 199339
rect 298660 199087 298661 199121
rect 298695 199087 298753 199121
rect 298787 199087 298816 199121
rect 298660 198869 298799 199087
rect 298660 198761 298661 198869
rect 298695 198727 298799 198835
rect 298660 198577 298799 198727
rect 298660 198543 298661 198577
rect 298695 198543 298753 198577
rect 298787 198543 298816 198577
rect 298660 198393 298799 198543
rect 298660 198251 298661 198359
rect 298695 198285 298799 198393
rect 298660 198033 298799 198251
rect 298660 197999 298661 198033
rect 298695 197999 298753 198033
rect 298787 197999 298816 198033
rect 298660 197781 298799 197999
rect 298660 197673 298661 197781
rect 298695 197639 298799 197747
rect 298660 197489 298799 197639
rect 298660 197455 298661 197489
rect 298695 197455 298753 197489
rect 298787 197455 298816 197489
rect 298660 197305 298799 197455
rect 298660 197163 298661 197271
rect 298695 197197 298799 197305
rect 298660 196945 298799 197163
rect 298660 196911 298661 196945
rect 298695 196911 298753 196945
rect 298787 196911 298816 196945
rect 298660 196693 298799 196911
rect 298660 196585 298661 196693
rect 298695 196551 298799 196659
rect 298660 196401 298799 196551
rect 298660 196367 298661 196401
rect 298695 196367 298753 196401
rect 298787 196367 298816 196401
rect 298660 196217 298799 196367
rect 298660 196075 298661 196183
rect 298695 196109 298799 196217
rect 298660 195857 298799 196075
rect 298660 195823 298661 195857
rect 298695 195823 298753 195857
rect 298787 195823 298816 195857
rect 298660 195605 298799 195823
rect 298660 195497 298661 195605
rect 298695 195463 298799 195571
rect 298660 195313 298799 195463
rect 298660 195279 298661 195313
rect 298695 195279 298753 195313
rect 298787 195279 298816 195313
rect 298660 195129 298799 195279
rect 298660 194987 298661 195095
rect 298695 195021 298799 195129
rect 298660 194769 298799 194987
rect 298660 194735 298661 194769
rect 298695 194735 298753 194769
rect 298787 194735 298816 194769
rect 298660 194517 298799 194735
rect 298660 194409 298661 194517
rect 298695 194375 298799 194483
rect 298660 194225 298799 194375
rect 298660 194191 298661 194225
rect 298695 194191 298753 194225
rect 298787 194191 298816 194225
rect 298660 194041 298799 194191
rect 298660 193899 298661 194007
rect 298695 193933 298799 194041
rect 298660 193681 298799 193899
rect 298660 193647 298661 193681
rect 298695 193647 298753 193681
rect 298787 193647 298816 193681
rect 298660 193429 298799 193647
rect 298660 193321 298661 193429
rect 298695 193287 298799 193395
rect 298660 193137 298799 193287
rect 298660 193103 298661 193137
rect 298695 193103 298753 193137
rect 298787 193103 298816 193137
rect 298660 192953 298799 193103
rect 298660 192811 298661 192919
rect 298695 192845 298799 192953
rect 298660 192593 298799 192811
rect 298660 192559 298661 192593
rect 298695 192559 298753 192593
rect 298787 192559 298816 192593
rect 298660 192341 298799 192559
rect 298660 192233 298661 192341
rect 298695 192199 298799 192307
rect 298660 192049 298799 192199
rect 298660 192015 298661 192049
rect 298695 192015 298753 192049
rect 298787 192015 298816 192049
rect 298660 191865 298799 192015
rect 298660 191723 298661 191831
rect 298695 191757 298799 191865
rect 298660 191505 298799 191723
rect 298660 191471 298661 191505
rect 298695 191471 298753 191505
rect 298787 191471 298816 191505
rect 298660 191253 298799 191471
rect 298660 191145 298661 191253
rect 298695 191111 298799 191219
rect 298660 190961 298799 191111
rect 298660 190927 298661 190961
rect 298695 190927 298753 190961
rect 298787 190927 298816 190961
rect 298660 190777 298799 190927
rect 298660 190635 298661 190743
rect 298695 190669 298799 190777
rect 298660 190417 298799 190635
rect 298660 190383 298661 190417
rect 298695 190383 298753 190417
rect 298787 190383 298816 190417
rect 298660 190165 298799 190383
rect 298660 190057 298661 190165
rect 298695 190023 298799 190131
rect 298660 189873 298799 190023
rect 298660 189839 298661 189873
rect 298695 189839 298753 189873
rect 298787 189839 298816 189873
rect 298660 189689 298799 189839
rect 298660 189547 298661 189655
rect 298695 189581 298799 189689
rect 298660 189329 298799 189547
rect 298660 189295 298661 189329
rect 298695 189295 298753 189329
rect 298787 189295 298816 189329
rect 298660 189077 298799 189295
rect 298660 188969 298661 189077
rect 298695 188935 298799 189043
rect 298660 188785 298799 188935
rect 298660 188751 298661 188785
rect 298695 188751 298753 188785
rect 298787 188751 298816 188785
rect 298660 188601 298799 188751
rect 298660 188459 298661 188567
rect 298695 188493 298799 188601
rect 298660 188241 298799 188459
rect 298660 188207 298661 188241
rect 298695 188207 298753 188241
rect 298787 188207 298816 188241
rect 298660 187989 298799 188207
rect 298660 187881 298661 187989
rect 298695 187847 298799 187955
rect 298660 187697 298799 187847
rect 298660 187663 298661 187697
rect 298695 187663 298753 187697
rect 298787 187663 298816 187697
rect 298660 187513 298799 187663
rect 298660 187371 298661 187479
rect 298695 187405 298799 187513
rect 298660 187153 298799 187371
rect 298660 187119 298661 187153
rect 298695 187119 298753 187153
rect 298787 187119 298816 187153
rect 298660 186901 298799 187119
rect 298660 186793 298661 186901
rect 298695 186759 298799 186867
rect 298660 186609 298799 186759
rect 298660 186575 298661 186609
rect 298695 186575 298753 186609
rect 298787 186575 298816 186609
rect 298660 186425 298799 186575
rect 298660 186283 298661 186391
rect 298695 186317 298799 186425
rect 298660 186065 298799 186283
rect 298660 186031 298661 186065
rect 298695 186031 298753 186065
rect 298787 186031 298816 186065
rect 298660 185813 298799 186031
rect 298660 185705 298661 185813
rect 298695 185671 298799 185779
rect 298660 185521 298799 185671
rect 298660 185487 298661 185521
rect 298695 185487 298753 185521
rect 298787 185487 298816 185521
rect 298660 185337 298799 185487
rect 298660 185195 298661 185303
rect 298695 185229 298799 185337
rect 298660 184977 298799 185195
rect 298660 184943 298661 184977
rect 298695 184943 298753 184977
rect 298787 184943 298816 184977
rect 298660 184725 298799 184943
rect 298660 184617 298661 184725
rect 298695 184583 298799 184691
rect 298660 184433 298799 184583
rect 298660 184399 298661 184433
rect 298695 184399 298753 184433
rect 298787 184399 298816 184433
rect 298660 184249 298799 184399
rect 298660 184107 298661 184215
rect 298695 184141 298799 184249
rect 298660 183889 298799 184107
rect 298660 183855 298661 183889
rect 298695 183855 298753 183889
rect 298787 183855 298816 183889
rect 298660 183637 298799 183855
rect 298660 183529 298661 183637
rect 298695 183495 298799 183603
rect 298660 183345 298799 183495
rect 298660 183311 298661 183345
rect 298695 183311 298753 183345
rect 298787 183311 298816 183345
rect 298660 183161 298799 183311
rect 298660 183019 298661 183127
rect 298695 183053 298799 183161
rect 298660 182801 298799 183019
rect 298660 182767 298661 182801
rect 298695 182767 298753 182801
rect 298787 182767 298816 182801
rect 298660 182549 298799 182767
rect 298660 182441 298661 182549
rect 298695 182407 298799 182515
rect 298660 182257 298799 182407
rect 298660 182223 298661 182257
rect 298695 182223 298753 182257
rect 298787 182223 298816 182257
rect 298660 182073 298799 182223
rect 298660 181931 298661 182039
rect 298695 181965 298799 182073
rect 298660 181713 298799 181931
rect 298660 181679 298661 181713
rect 298695 181679 298753 181713
rect 298787 181679 298816 181713
rect 298660 181461 298799 181679
rect 298660 181353 298661 181461
rect 298695 181319 298799 181427
rect 298660 181169 298799 181319
rect 298660 181135 298661 181169
rect 298695 181135 298753 181169
rect 298787 181135 298816 181169
rect 298660 180985 298799 181135
rect 298660 180843 298661 180951
rect 298695 180877 298799 180985
rect 298660 180625 298799 180843
rect 298660 180591 298661 180625
rect 298695 180591 298753 180625
rect 298787 180591 298816 180625
rect 298660 180373 298799 180591
rect 298660 180265 298661 180373
rect 298695 180231 298799 180339
rect 298660 180081 298799 180231
rect 298660 180047 298661 180081
rect 298695 180047 298753 180081
rect 298787 180047 298816 180081
rect 298660 179897 298799 180047
rect 298660 179755 298661 179863
rect 298695 179789 298799 179897
rect 298660 179537 298799 179755
rect 298660 179503 298661 179537
rect 298695 179503 298753 179537
rect 298787 179503 298816 179537
rect 298660 179285 298799 179503
rect 298660 179177 298661 179285
rect 298695 179143 298799 179251
rect 298660 178993 298799 179143
rect 298660 178959 298661 178993
rect 298695 178959 298753 178993
rect 298787 178959 298816 178993
rect 298660 178809 298799 178959
rect 298660 178667 298661 178775
rect 298695 178701 298799 178809
rect 298660 178449 298799 178667
rect 298660 178415 298661 178449
rect 298695 178415 298753 178449
rect 298787 178415 298816 178449
rect 298660 178197 298799 178415
rect 298660 178089 298661 178197
rect 298695 178055 298799 178163
rect 298660 177905 298799 178055
rect 298660 177871 298661 177905
rect 298695 177871 298753 177905
rect 298787 177871 298816 177905
rect 298660 177721 298799 177871
rect 298660 177579 298661 177687
rect 298695 177613 298799 177721
rect 298660 177361 298799 177579
rect 298660 177327 298661 177361
rect 298695 177327 298753 177361
rect 298787 177327 298816 177361
rect 298660 177109 298799 177327
rect 298660 177001 298661 177109
rect 298695 176967 298799 177075
rect 298660 176817 298799 176967
rect 298660 176783 298661 176817
rect 298695 176783 298753 176817
rect 298787 176783 298816 176817
rect 298660 176633 298799 176783
rect 298660 176491 298661 176599
rect 298695 176525 298799 176633
rect 298660 176273 298799 176491
rect 298660 176239 298661 176273
rect 298695 176239 298753 176273
rect 298787 176239 298816 176273
rect 298660 176021 298799 176239
rect 298660 175913 298661 176021
rect 298695 175879 298799 175987
rect 298660 175729 298799 175879
rect 298660 175695 298661 175729
rect 298695 175695 298753 175729
rect 298787 175695 298816 175729
rect 298660 175545 298799 175695
rect 298660 175403 298661 175511
rect 298695 175437 298799 175545
rect 298660 175185 298799 175403
rect 298660 175151 298661 175185
rect 298695 175151 298753 175185
rect 298787 175151 298816 175185
rect 298660 174933 298799 175151
rect 298660 174825 298661 174933
rect 298695 174791 298799 174899
rect 298660 174641 298799 174791
rect 298660 174607 298661 174641
rect 298695 174607 298753 174641
rect 298787 174607 298816 174641
rect 298660 174457 298799 174607
rect 298660 174315 298661 174423
rect 298695 174349 298799 174457
rect 298660 174097 298799 174315
rect 298660 174063 298661 174097
rect 298695 174063 298753 174097
rect 298787 174063 298816 174097
rect 298660 173845 298799 174063
rect 298660 173737 298661 173845
rect 298695 173703 298799 173811
rect 298660 173553 298799 173703
rect 298660 173519 298661 173553
rect 298695 173519 298753 173553
rect 298787 173519 298816 173553
rect 298660 173369 298799 173519
rect 298660 173227 298661 173335
rect 298695 173261 298799 173369
rect 298660 173009 298799 173227
rect 298660 172975 298661 173009
rect 298695 172975 298753 173009
rect 298787 172975 298816 173009
rect 298660 172757 298799 172975
rect 298660 172649 298661 172757
rect 298695 172615 298799 172723
rect 298660 172465 298799 172615
rect 298660 172431 298661 172465
rect 298695 172431 298753 172465
rect 298787 172431 298816 172465
rect 298660 172281 298799 172431
rect 298660 172139 298661 172247
rect 298695 172173 298799 172281
rect 298660 171921 298799 172139
rect 298660 171887 298661 171921
rect 298695 171887 298753 171921
rect 298787 171887 298816 171921
rect 298660 171669 298799 171887
rect 298660 171561 298661 171669
rect 298695 171527 298799 171635
rect 298660 171377 298799 171527
rect 298660 171343 298661 171377
rect 298695 171343 298753 171377
rect 298787 171343 298816 171377
rect 298660 171193 298799 171343
rect 298660 171051 298661 171159
rect 298695 171085 298799 171193
rect 298660 170833 298799 171051
rect 298660 170799 298661 170833
rect 298695 170799 298753 170833
rect 298787 170799 298816 170833
rect 298660 170581 298799 170799
rect 298660 170473 298661 170581
rect 298695 170439 298799 170547
rect 298660 170289 298799 170439
rect 298660 170255 298661 170289
rect 298695 170255 298753 170289
rect 298787 170255 298816 170289
rect 298660 170105 298799 170255
rect 298660 169963 298661 170071
rect 298695 169997 298799 170105
rect 298660 169745 298799 169963
rect 298660 169711 298661 169745
rect 298695 169711 298753 169745
rect 298787 169711 298816 169745
rect 298660 169493 298799 169711
rect 298660 169385 298661 169493
rect 298695 169351 298799 169459
rect 298660 169201 298799 169351
rect 298660 169167 298661 169201
rect 298695 169167 298753 169201
rect 298787 169167 298816 169201
rect 298660 169017 298799 169167
rect 298660 168875 298661 168983
rect 298695 168909 298799 169017
rect 298660 168657 298799 168875
rect 298660 168623 298661 168657
rect 298695 168623 298753 168657
rect 298787 168623 298816 168657
rect 298660 168405 298799 168623
rect 298660 168297 298661 168405
rect 298695 168263 298799 168371
rect 298660 168113 298799 168263
rect 298660 168079 298661 168113
rect 298695 168079 298753 168113
rect 298787 168079 298816 168113
rect 298660 167929 298799 168079
rect 298660 167787 298661 167895
rect 298695 167821 298799 167929
rect 298660 167569 298799 167787
rect 298660 167535 298661 167569
rect 298695 167535 298753 167569
rect 298787 167535 298816 167569
rect 298660 167317 298799 167535
rect 298660 167209 298661 167317
rect 298695 167175 298799 167283
rect 298660 167025 298799 167175
rect 298660 166991 298661 167025
rect 298695 166991 298753 167025
rect 298787 166991 298816 167025
rect 298660 166841 298799 166991
rect 298660 166699 298661 166807
rect 298695 166733 298799 166841
rect 298660 166481 298799 166699
rect 298660 166447 298661 166481
rect 298695 166447 298753 166481
rect 298787 166447 298816 166481
rect 298660 166229 298799 166447
rect 298660 166121 298661 166229
rect 298695 166087 298799 166195
rect 298660 165937 298799 166087
rect 298660 165903 298661 165937
rect 298695 165903 298753 165937
rect 298787 165903 298816 165937
rect 298660 165753 298799 165903
rect 298660 165611 298661 165719
rect 298695 165645 298799 165753
rect 298660 165393 298799 165611
rect 298660 165359 298661 165393
rect 298695 165359 298753 165393
rect 298787 165359 298816 165393
rect 298660 165141 298799 165359
rect 298660 165033 298661 165141
rect 298695 164999 298799 165107
rect 298660 164849 298799 164999
rect 298660 164815 298661 164849
rect 298695 164815 298753 164849
rect 298787 164815 298816 164849
rect 298660 164665 298799 164815
rect 298660 164523 298661 164631
rect 298695 164557 298799 164665
rect 298660 164305 298799 164523
rect 298660 164271 298661 164305
rect 298695 164271 298753 164305
rect 298787 164271 298816 164305
rect 298660 164053 298799 164271
rect 298660 163945 298661 164053
rect 298695 163911 298799 164019
rect 298660 163761 298799 163911
rect 298660 163727 298661 163761
rect 298695 163727 298753 163761
rect 298787 163727 298816 163761
rect 298660 163577 298799 163727
rect 298660 163435 298661 163543
rect 298695 163469 298799 163577
rect 298660 163217 298799 163435
rect 298660 163183 298661 163217
rect 298695 163183 298753 163217
rect 298787 163183 298816 163217
rect 298660 162965 298799 163183
rect 298660 162857 298661 162965
rect 298695 162823 298799 162931
rect 298660 162673 298799 162823
rect 298660 162639 298661 162673
rect 298695 162639 298753 162673
rect 298787 162639 298816 162673
rect 298660 162489 298799 162639
rect 298660 162347 298661 162455
rect 298695 162381 298799 162489
rect 298660 162129 298799 162347
rect 298660 162095 298661 162129
rect 298695 162095 298753 162129
rect 298787 162095 298816 162129
rect 298660 161877 298799 162095
rect 298660 161769 298661 161877
rect 298695 161735 298799 161843
rect 298660 161585 298799 161735
rect 298660 161551 298661 161585
rect 298695 161551 298753 161585
rect 298787 161551 298816 161585
rect 298660 161401 298799 161551
rect 298660 161259 298661 161367
rect 298695 161293 298799 161401
rect 298660 161041 298799 161259
rect 298660 161007 298661 161041
rect 298695 161007 298753 161041
rect 298787 161007 298816 161041
rect 298660 160789 298799 161007
rect 298660 160681 298661 160789
rect 298695 160647 298799 160755
rect 298660 160497 298799 160647
rect 298660 160463 298661 160497
rect 298695 160463 298753 160497
rect 298787 160463 298816 160497
rect 298660 160313 298799 160463
rect 298660 160171 298661 160279
rect 298695 160205 298799 160313
rect 298660 159953 298799 160171
rect 298660 159919 298661 159953
rect 298695 159919 298753 159953
rect 298787 159919 298816 159953
rect 298660 159701 298799 159919
rect 298660 159593 298661 159701
rect 298695 159559 298799 159667
rect 298660 159409 298799 159559
rect 298660 159375 298661 159409
rect 298695 159375 298753 159409
rect 298787 159375 298816 159409
rect 298660 159225 298799 159375
rect 298660 159083 298661 159191
rect 298695 159117 298799 159225
rect 298660 158865 298799 159083
rect 298660 158831 298661 158865
rect 298695 158831 298753 158865
rect 298787 158831 298816 158865
rect 298660 158613 298799 158831
rect 298660 158505 298661 158613
rect 298695 158471 298799 158579
rect 298660 158321 298799 158471
rect 298660 158287 298661 158321
rect 298695 158287 298753 158321
rect 298787 158287 298816 158321
rect 298660 158137 298799 158287
rect 298660 157995 298661 158103
rect 298695 158029 298799 158137
rect 298660 157777 298799 157995
rect 298660 157743 298661 157777
rect 298695 157743 298753 157777
rect 298787 157743 298816 157777
rect 298660 157525 298799 157743
rect 298660 157417 298661 157525
rect 298695 157383 298799 157491
rect 298660 157233 298799 157383
rect 298660 157199 298661 157233
rect 298695 157199 298753 157233
rect 298787 157199 298816 157233
rect 298660 157049 298799 157199
rect 298660 156907 298661 157015
rect 298695 156941 298799 157049
rect 298660 156689 298799 156907
rect 298660 156655 298661 156689
rect 298695 156655 298753 156689
rect 298787 156655 298816 156689
rect 298660 156437 298799 156655
rect 298660 156329 298661 156437
rect 298695 156295 298799 156403
rect 298660 156145 298799 156295
rect 298660 156111 298661 156145
rect 298695 156111 298753 156145
rect 298787 156111 298816 156145
rect 298660 155961 298799 156111
rect 298660 155819 298661 155927
rect 298695 155853 298799 155961
rect 298660 155601 298799 155819
rect 298660 155567 298661 155601
rect 298695 155567 298753 155601
rect 298787 155567 298816 155601
rect 298660 155349 298799 155567
rect 298660 155241 298661 155349
rect 298695 155207 298799 155315
rect 298660 155057 298799 155207
rect 298660 155023 298661 155057
rect 298695 155023 298753 155057
rect 298787 155023 298816 155057
rect 298660 154873 298799 155023
rect 298660 154731 298661 154839
rect 298695 154765 298799 154873
rect 298660 154513 298799 154731
rect 298660 154479 298661 154513
rect 298695 154479 298753 154513
rect 298787 154479 298816 154513
rect 298660 154261 298799 154479
rect 298660 154153 298661 154261
rect 298695 154119 298799 154227
rect 298660 153969 298799 154119
rect 298660 153935 298661 153969
rect 298695 153935 298753 153969
rect 298787 153935 298816 153969
rect 298660 153785 298799 153935
rect 298660 153643 298661 153751
rect 298695 153677 298799 153785
rect 298660 153425 298799 153643
rect 298660 153391 298661 153425
rect 298695 153391 298753 153425
rect 298787 153391 298816 153425
rect 298660 153173 298799 153391
rect 298660 153065 298661 153173
rect 298695 153031 298799 153139
rect 298660 152881 298799 153031
rect 298660 152847 298661 152881
rect 298695 152847 298753 152881
rect 298787 152847 298816 152881
rect 298660 152697 298799 152847
rect 298660 152555 298661 152663
rect 298695 152589 298799 152697
rect 298660 152337 298799 152555
rect 298660 152303 298661 152337
rect 298695 152303 298753 152337
rect 298787 152303 298816 152337
rect 298660 152085 298799 152303
rect 298660 151977 298661 152085
rect 298695 151943 298799 152051
rect 298660 151793 298799 151943
rect 298660 151759 298661 151793
rect 298695 151759 298753 151793
rect 298787 151759 298816 151793
rect 298660 151609 298799 151759
rect 298660 151467 298661 151575
rect 298695 151501 298799 151609
rect 298660 151249 298799 151467
rect 298660 151215 298661 151249
rect 298695 151215 298753 151249
rect 298787 151215 298816 151249
rect 298660 150997 298799 151215
rect 298660 150889 298661 150997
rect 298695 150855 298799 150963
rect 298660 150705 298799 150855
rect 298660 150671 298661 150705
rect 298695 150671 298753 150705
rect 298787 150671 298816 150705
rect 298660 150521 298799 150671
rect 298660 150379 298661 150487
rect 298695 150413 298799 150521
rect 298660 150161 298799 150379
rect 298660 150127 298661 150161
rect 298695 150127 298753 150161
rect 298787 150127 298816 150161
rect 298660 149909 298799 150127
rect 298660 149801 298661 149909
rect 298695 149767 298799 149875
rect 298660 149617 298799 149767
rect 298660 149583 298661 149617
rect 298695 149583 298753 149617
rect 298787 149583 298816 149617
rect 298660 149433 298799 149583
rect 298660 149291 298661 149399
rect 298695 149325 298799 149433
rect 298660 149073 298799 149291
rect 298660 149039 298661 149073
rect 298695 149039 298753 149073
rect 298787 149039 298816 149073
rect 298660 148821 298799 149039
rect 298660 148713 298661 148821
rect 298695 148679 298799 148787
rect 298660 148529 298799 148679
rect 298660 148495 298661 148529
rect 298695 148495 298753 148529
rect 298787 148495 298816 148529
rect 298660 148345 298799 148495
rect 298660 148203 298661 148311
rect 298695 148237 298799 148345
rect 298660 147985 298799 148203
rect 298660 147951 298661 147985
rect 298695 147951 298753 147985
rect 298787 147951 298816 147985
rect 298660 147733 298799 147951
rect 298660 147625 298661 147733
rect 298695 147591 298799 147699
rect 298660 147441 298799 147591
rect 298660 147407 298661 147441
rect 298695 147407 298753 147441
rect 298787 147407 298816 147441
rect 298660 147257 298799 147407
rect 298660 147115 298661 147223
rect 298695 147149 298799 147257
rect 298660 146897 298799 147115
rect 298660 146863 298661 146897
rect 298695 146863 298753 146897
rect 298787 146863 298816 146897
rect 298660 146645 298799 146863
rect 298660 146537 298661 146645
rect 298695 146503 298799 146611
rect 298660 146353 298799 146503
rect 298660 146319 298661 146353
rect 298695 146319 298753 146353
rect 298787 146319 298816 146353
rect 298660 146169 298799 146319
rect 298660 146027 298661 146135
rect 298695 146061 298799 146169
rect 298660 145809 298799 146027
rect 298660 145775 298661 145809
rect 298695 145775 298753 145809
rect 298787 145775 298816 145809
rect 298660 145557 298799 145775
rect 298660 145449 298661 145557
rect 298695 145415 298799 145523
rect 298660 145265 298799 145415
rect 298660 145231 298661 145265
rect 298695 145231 298753 145265
rect 298787 145231 298816 145265
rect 298660 145081 298799 145231
rect 298660 144939 298661 145047
rect 298695 144973 298799 145081
rect 298660 144721 298799 144939
rect 298660 144687 298661 144721
rect 298695 144687 298753 144721
rect 298787 144687 298816 144721
rect 298660 144469 298799 144687
rect 298660 144361 298661 144469
rect 298695 144327 298799 144435
rect 298660 144177 298799 144327
rect 298660 144143 298661 144177
rect 298695 144143 298753 144177
rect 298787 144143 298816 144177
rect 298660 143993 298799 144143
rect 298660 143851 298661 143959
rect 298695 143885 298799 143993
rect 298660 143633 298799 143851
rect 298660 143599 298661 143633
rect 298695 143599 298753 143633
rect 298787 143599 298816 143633
rect 298660 143381 298799 143599
rect 298660 143273 298661 143381
rect 298695 143239 298799 143347
rect 298660 143089 298799 143239
rect 298660 143055 298661 143089
rect 298695 143055 298753 143089
rect 298787 143055 298816 143089
rect 298660 142905 298799 143055
rect 298660 142763 298661 142871
rect 298695 142797 298799 142905
rect 298660 142545 298799 142763
rect 298660 142511 298661 142545
rect 298695 142511 298753 142545
rect 298787 142511 298816 142545
rect 298660 142293 298799 142511
rect 298660 142185 298661 142293
rect 298695 142151 298799 142259
rect 298660 142001 298799 142151
rect 298660 141967 298661 142001
rect 298695 141967 298753 142001
rect 298787 141967 298816 142001
rect 298660 141817 298799 141967
rect 298660 141675 298661 141783
rect 298695 141709 298799 141817
rect 298660 141457 298799 141675
rect 298660 141423 298661 141457
rect 298695 141423 298753 141457
rect 298787 141423 298816 141457
rect 298660 141205 298799 141423
rect 298660 141097 298661 141205
rect 298695 141063 298799 141171
rect 298660 140913 298799 141063
rect 298660 140879 298661 140913
rect 298695 140879 298753 140913
rect 298787 140879 298816 140913
rect 298660 140729 298799 140879
rect 298660 140587 298661 140695
rect 298695 140621 298799 140729
rect 298660 140369 298799 140587
rect 298660 140335 298661 140369
rect 298695 140335 298753 140369
rect 298787 140335 298816 140369
rect 298660 140117 298799 140335
rect 298660 140009 298661 140117
rect 298695 139975 298799 140083
rect 298660 139825 298799 139975
rect 298660 139791 298661 139825
rect 298695 139791 298753 139825
rect 298787 139791 298816 139825
rect 298660 139641 298799 139791
rect 298660 139499 298661 139607
rect 298695 139533 298799 139641
rect 298660 139281 298799 139499
rect 298660 139247 298661 139281
rect 298695 139247 298753 139281
rect 298787 139247 298816 139281
rect 298660 139029 298799 139247
rect 298660 138921 298661 139029
rect 298695 138887 298799 138995
rect 298660 138737 298799 138887
rect 298660 138703 298661 138737
rect 298695 138703 298753 138737
rect 298787 138703 298816 138737
rect 298660 138553 298799 138703
rect 298660 138411 298661 138519
rect 298695 138445 298799 138553
rect 298660 138193 298799 138411
rect 298660 138159 298661 138193
rect 298695 138159 298753 138193
rect 298787 138159 298816 138193
rect 298660 137941 298799 138159
rect 298660 137833 298661 137941
rect 298695 137799 298799 137907
rect 298660 137649 298799 137799
rect 298660 137615 298661 137649
rect 298695 137615 298753 137649
rect 298787 137615 298816 137649
rect 298660 137465 298799 137615
rect 298660 137323 298661 137431
rect 298695 137357 298799 137465
rect 298660 137105 298799 137323
rect 298660 137071 298661 137105
rect 298695 137071 298753 137105
rect 298787 137071 298816 137105
rect 298660 136853 298799 137071
rect 298660 136745 298661 136853
rect 298695 136711 298799 136819
rect 298660 136561 298799 136711
rect 298660 136527 298661 136561
rect 298695 136527 298753 136561
rect 298787 136527 298816 136561
rect 298660 136377 298799 136527
rect 298660 136235 298661 136343
rect 298695 136269 298799 136377
rect 298660 136017 298799 136235
rect 298660 135983 298661 136017
rect 298695 135983 298753 136017
rect 298787 135983 298816 136017
rect 298660 135765 298799 135983
rect 298660 135657 298661 135765
rect 298695 135623 298799 135731
rect 298660 135473 298799 135623
rect 298660 135439 298661 135473
rect 298695 135439 298753 135473
rect 298787 135439 298816 135473
rect 298660 135289 298799 135439
rect 298660 135147 298661 135255
rect 298695 135181 298799 135289
rect 298660 134929 298799 135147
rect 298660 134895 298661 134929
rect 298695 134895 298753 134929
rect 298787 134895 298816 134929
rect 298660 134677 298799 134895
rect 298660 134569 298661 134677
rect 298695 134535 298799 134643
rect 298660 134385 298799 134535
rect 298660 134351 298661 134385
rect 298695 134351 298753 134385
rect 298787 134351 298816 134385
rect 298660 134201 298799 134351
rect 298660 134059 298661 134167
rect 298695 134093 298799 134201
rect 298660 133841 298799 134059
rect 298660 133807 298661 133841
rect 298695 133807 298753 133841
rect 298787 133807 298816 133841
rect 298660 133589 298799 133807
rect 298660 133481 298661 133589
rect 298695 133447 298799 133555
rect 298660 133297 298799 133447
rect 298660 133263 298661 133297
rect 298695 133263 298753 133297
rect 298787 133263 298816 133297
rect 298660 133113 298799 133263
rect 298660 132971 298661 133079
rect 298695 133005 298799 133113
rect 298660 132753 298799 132971
rect 298660 132719 298661 132753
rect 298695 132719 298753 132753
rect 298787 132719 298816 132753
rect 298660 132501 298799 132719
rect 298660 132393 298661 132501
rect 298695 132359 298799 132467
rect 298660 132209 298799 132359
rect 298660 132175 298661 132209
rect 298695 132175 298753 132209
rect 298787 132175 298816 132209
rect 298660 132025 298799 132175
rect 298660 131883 298661 131991
rect 298695 131917 298799 132025
rect 298660 131665 298799 131883
rect 298660 131631 298661 131665
rect 298695 131631 298753 131665
rect 298787 131631 298816 131665
rect 298660 131413 298799 131631
rect 298660 131305 298661 131413
rect 298695 131271 298799 131379
rect 298660 131121 298799 131271
rect 298660 131087 298661 131121
rect 298695 131087 298753 131121
rect 298787 131087 298816 131121
rect 298660 130937 298799 131087
rect 298660 130795 298661 130903
rect 298695 130829 298799 130937
rect 298660 130577 298799 130795
rect 298660 130543 298661 130577
rect 298695 130543 298753 130577
rect 298787 130543 298816 130577
rect 298660 130325 298799 130543
rect 298660 130217 298661 130325
rect 298695 130183 298799 130291
rect 298660 130033 298799 130183
rect 298660 129999 298661 130033
rect 298695 129999 298753 130033
rect 298787 129999 298816 130033
rect 298660 129849 298799 129999
rect 298660 129707 298661 129815
rect 298695 129741 298799 129849
rect 298660 129489 298799 129707
rect 298660 129455 298661 129489
rect 298695 129455 298753 129489
rect 298787 129455 298816 129489
rect 298660 129237 298799 129455
rect 298660 129129 298661 129237
rect 298695 129095 298799 129203
rect 298660 128945 298799 129095
rect 298660 128911 298661 128945
rect 298695 128911 298753 128945
rect 298787 128911 298816 128945
rect 298660 128761 298799 128911
rect 298660 128619 298661 128727
rect 298695 128653 298799 128761
rect 298660 128401 298799 128619
rect 298660 128367 298661 128401
rect 298695 128367 298753 128401
rect 298787 128367 298816 128401
rect 298660 128149 298799 128367
rect 298660 128041 298661 128149
rect 298695 128007 298799 128115
rect 298660 127857 298799 128007
rect 298660 127823 298661 127857
rect 298695 127823 298753 127857
rect 298787 127823 298816 127857
rect 298660 127673 298799 127823
rect 298660 127531 298661 127639
rect 298695 127565 298799 127673
rect 298660 127313 298799 127531
rect 298660 127279 298661 127313
rect 298695 127279 298753 127313
rect 298787 127279 298816 127313
rect 298660 127061 298799 127279
rect 298660 126953 298661 127061
rect 298695 126919 298799 127027
rect 298660 126769 298799 126919
rect 298660 126735 298661 126769
rect 298695 126735 298753 126769
rect 298787 126735 298816 126769
rect 298660 126585 298799 126735
rect 298660 126443 298661 126551
rect 298695 126477 298799 126585
rect 298660 126225 298799 126443
rect 298660 126191 298661 126225
rect 298695 126191 298753 126225
rect 298787 126191 298816 126225
rect 298660 125973 298799 126191
rect 298660 125865 298661 125973
rect 298695 125831 298799 125939
rect 298660 125681 298799 125831
rect 298660 125647 298661 125681
rect 298695 125647 298753 125681
rect 298787 125647 298816 125681
rect 298660 125497 298799 125647
rect 298660 125355 298661 125463
rect 298695 125389 298799 125497
rect 298660 125137 298799 125355
rect 298660 125103 298661 125137
rect 298695 125103 298753 125137
rect 298787 125103 298816 125137
rect 298660 124885 298799 125103
rect 298660 124777 298661 124885
rect 298695 124743 298799 124851
rect 298660 124593 298799 124743
rect 298660 124559 298661 124593
rect 298695 124559 298753 124593
rect 298787 124559 298816 124593
rect 298660 124409 298799 124559
rect 298660 124267 298661 124375
rect 298695 124301 298799 124409
rect 298660 124049 298799 124267
rect 298660 124015 298661 124049
rect 298695 124015 298753 124049
rect 298787 124015 298816 124049
rect 298660 123797 298799 124015
rect 298660 123689 298661 123797
rect 298695 123655 298799 123763
rect 298660 123505 298799 123655
rect 298660 123471 298661 123505
rect 298695 123471 298753 123505
rect 298787 123471 298816 123505
rect 298660 123321 298799 123471
rect 298660 123179 298661 123287
rect 298695 123213 298799 123321
rect 298660 122961 298799 123179
rect 298660 122927 298661 122961
rect 298695 122927 298753 122961
rect 298787 122927 298816 122961
rect 298660 122709 298799 122927
rect 298660 122601 298661 122709
rect 298695 122567 298799 122675
rect 298660 122417 298799 122567
rect 298660 122383 298661 122417
rect 298695 122383 298753 122417
rect 298787 122383 298816 122417
rect 298660 122233 298799 122383
rect 298660 122091 298661 122199
rect 298695 122125 298799 122233
rect 298660 121873 298799 122091
rect 298660 121839 298661 121873
rect 298695 121839 298753 121873
rect 298787 121839 298816 121873
rect 298660 121621 298799 121839
rect 298660 121513 298661 121621
rect 298695 121479 298799 121587
rect 298660 121329 298799 121479
rect 298660 121295 298661 121329
rect 298695 121295 298753 121329
rect 298787 121295 298816 121329
rect 298660 121145 298799 121295
rect 298660 121003 298661 121111
rect 298695 121037 298799 121145
rect 298660 120785 298799 121003
rect 298660 120751 298661 120785
rect 298695 120751 298753 120785
rect 298787 120751 298816 120785
rect 298660 120533 298799 120751
rect 298660 120425 298661 120533
rect 298695 120391 298799 120499
rect 298660 120241 298799 120391
rect 298660 120207 298661 120241
rect 298695 120207 298753 120241
rect 298787 120207 298816 120241
rect 298660 120057 298799 120207
rect 298660 119915 298661 120023
rect 298695 119949 298799 120057
rect 298660 119697 298799 119915
rect 298660 119663 298661 119697
rect 298695 119663 298753 119697
rect 298787 119663 298816 119697
rect 298660 119445 298799 119663
rect 298660 119337 298661 119445
rect 298695 119303 298799 119411
rect 298660 119153 298799 119303
rect 298660 119119 298661 119153
rect 298695 119119 298753 119153
rect 298787 119119 298816 119153
rect 298660 118969 298799 119119
rect 298660 118827 298661 118935
rect 298695 118861 298799 118969
rect 298660 118609 298799 118827
rect 298660 118575 298661 118609
rect 298695 118575 298753 118609
rect 298787 118575 298816 118609
rect 298660 118357 298799 118575
rect 298660 118249 298661 118357
rect 298695 118215 298799 118323
rect 298660 118065 298799 118215
rect 298660 118031 298661 118065
rect 298695 118031 298753 118065
rect 298787 118031 298816 118065
rect 298660 117881 298799 118031
rect 298660 117739 298661 117847
rect 298695 117773 298799 117881
rect 298660 117521 298799 117739
rect 298660 117487 298661 117521
rect 298695 117487 298753 117521
rect 298787 117487 298816 117521
rect 298660 117269 298799 117487
rect 298660 117161 298661 117269
rect 298695 117127 298799 117235
rect 298660 116977 298799 117127
rect 298660 116943 298661 116977
rect 298695 116943 298753 116977
rect 298787 116943 298816 116977
rect 298660 116793 298799 116943
rect 298660 116651 298661 116759
rect 298695 116685 298799 116793
rect 298660 116433 298799 116651
rect 298660 116399 298661 116433
rect 298695 116399 298753 116433
rect 298787 116399 298816 116433
rect 298660 116181 298799 116399
rect 298660 116073 298661 116181
rect 298695 116039 298799 116147
rect 298660 115889 298799 116039
rect 298660 115855 298661 115889
rect 298695 115855 298753 115889
rect 298787 115855 298816 115889
rect 298660 115705 298799 115855
rect 298660 115563 298661 115671
rect 298695 115597 298799 115705
rect 298660 115345 298799 115563
rect 298660 115311 298661 115345
rect 298695 115311 298753 115345
rect 298787 115311 298816 115345
rect 298660 115093 298799 115311
rect 298660 114985 298661 115093
rect 298695 114951 298799 115059
rect 298660 114801 298799 114951
rect 298660 114767 298661 114801
rect 298695 114767 298753 114801
rect 298787 114767 298816 114801
rect 298660 114617 298799 114767
rect 298660 114475 298661 114583
rect 298695 114509 298799 114617
rect 298660 114257 298799 114475
rect 298660 114223 298661 114257
rect 298695 114223 298753 114257
rect 298787 114223 298816 114257
rect 298660 114005 298799 114223
rect 298660 113897 298661 114005
rect 298695 113863 298799 113971
rect 298660 113713 298799 113863
rect 298660 113679 298661 113713
rect 298695 113679 298753 113713
rect 298787 113679 298816 113713
rect 298660 113529 298799 113679
rect 298660 113387 298661 113495
rect 298695 113421 298799 113529
rect 298660 113169 298799 113387
rect 298660 113135 298661 113169
rect 298695 113135 298753 113169
rect 298787 113135 298816 113169
rect 298660 112917 298799 113135
rect 298660 112809 298661 112917
rect 298695 112775 298799 112883
rect 298660 112625 298799 112775
rect 298660 112591 298661 112625
rect 298695 112591 298753 112625
rect 298787 112591 298816 112625
rect 298660 112441 298799 112591
rect 298660 112299 298661 112407
rect 298695 112333 298799 112441
rect 298660 112081 298799 112299
rect 298660 112047 298661 112081
rect 298695 112047 298753 112081
rect 298787 112047 298816 112081
rect 298660 111829 298799 112047
rect 298660 111721 298661 111829
rect 298695 111687 298799 111795
rect 298660 111537 298799 111687
rect 298660 111503 298661 111537
rect 298695 111503 298753 111537
rect 298787 111503 298816 111537
rect 298660 111353 298799 111503
rect 298660 111211 298661 111319
rect 298695 111245 298799 111353
rect 298660 110993 298799 111211
rect 298660 110959 298661 110993
rect 298695 110959 298753 110993
rect 298787 110959 298816 110993
rect 298660 110741 298799 110959
rect 298660 110633 298661 110741
rect 298695 110599 298799 110707
rect 298660 110449 298799 110599
rect 298660 110415 298661 110449
rect 298695 110415 298753 110449
rect 298787 110415 298816 110449
rect 298660 110265 298799 110415
rect 298660 110123 298661 110231
rect 298695 110157 298799 110265
rect 298660 109905 298799 110123
rect 298660 109871 298661 109905
rect 298695 109871 298753 109905
rect 298787 109871 298816 109905
rect 298660 109653 298799 109871
rect 298660 109545 298661 109653
rect 298695 109511 298799 109619
rect 298660 109361 298799 109511
rect 298660 109327 298661 109361
rect 298695 109327 298753 109361
rect 298787 109327 298816 109361
rect 298660 109177 298799 109327
rect 298660 109035 298661 109143
rect 298695 109069 298799 109177
rect 298660 108817 298799 109035
rect 298660 108783 298661 108817
rect 298695 108783 298753 108817
rect 298787 108783 298816 108817
rect 298660 108565 298799 108783
rect 298660 108457 298661 108565
rect 298695 108423 298799 108531
rect 298660 108273 298799 108423
rect 298660 108239 298661 108273
rect 298695 108239 298753 108273
rect 298787 108239 298816 108273
rect 298660 108089 298799 108239
rect 298660 107947 298661 108055
rect 298695 107981 298799 108089
rect 298660 107729 298799 107947
rect 298660 107695 298661 107729
rect 298695 107695 298753 107729
rect 298787 107695 298816 107729
rect 298660 107477 298799 107695
rect 298660 107369 298661 107477
rect 298695 107335 298799 107443
rect 298660 107185 298799 107335
rect 298660 107151 298661 107185
rect 298695 107151 298753 107185
rect 298787 107151 298816 107185
rect 298660 107001 298799 107151
rect 298660 106859 298661 106967
rect 298695 106893 298799 107001
rect 298660 106641 298799 106859
rect 298660 106607 298661 106641
rect 298695 106607 298753 106641
rect 298787 106607 298816 106641
rect 298660 106389 298799 106607
rect 298660 106281 298661 106389
rect 298695 106247 298799 106355
rect 298660 106097 298799 106247
rect 298660 106063 298661 106097
rect 298695 106063 298753 106097
rect 298787 106063 298816 106097
rect 298660 105913 298799 106063
rect 298660 105771 298661 105879
rect 298695 105805 298799 105913
rect 298660 105553 298799 105771
rect 298660 105519 298661 105553
rect 298695 105519 298753 105553
rect 298787 105519 298816 105553
rect 298660 105301 298799 105519
rect 298660 105193 298661 105301
rect 298695 105159 298799 105267
rect 298660 105009 298799 105159
rect 298660 104975 298661 105009
rect 298695 104975 298753 105009
rect 298787 104975 298816 105009
rect 298660 104825 298799 104975
rect 298660 104683 298661 104791
rect 298695 104717 298799 104825
rect 298660 104465 298799 104683
rect 298660 104431 298661 104465
rect 298695 104431 298753 104465
rect 298787 104431 298816 104465
rect 298660 104213 298799 104431
rect 298660 104105 298661 104213
rect 298695 104071 298799 104179
rect 298660 103921 298799 104071
rect 298660 103887 298661 103921
rect 298695 103887 298753 103921
rect 298787 103887 298816 103921
rect 298660 103737 298799 103887
rect 298660 103595 298661 103703
rect 298695 103629 298799 103737
rect 298660 103377 298799 103595
rect 298660 103343 298661 103377
rect 298695 103343 298753 103377
rect 298787 103343 298816 103377
rect 298660 103125 298799 103343
rect 298660 103017 298661 103125
rect 298695 102983 298799 103091
rect 298660 102833 298799 102983
rect 298660 102799 298661 102833
rect 298695 102799 298753 102833
rect 298787 102799 298816 102833
rect 298660 102649 298799 102799
rect 298660 102507 298661 102615
rect 298695 102541 298799 102649
rect 298660 102289 298799 102507
rect 298660 102255 298661 102289
rect 298695 102255 298753 102289
rect 298787 102255 298816 102289
rect 298660 102037 298799 102255
rect 298660 101929 298661 102037
rect 298695 101895 298799 102003
rect 298660 101745 298799 101895
rect 298660 101711 298661 101745
rect 298695 101711 298753 101745
rect 298787 101711 298816 101745
rect 298660 101561 298799 101711
rect 298660 101419 298661 101527
rect 298695 101453 298799 101561
rect 298660 101201 298799 101419
rect 298660 101167 298661 101201
rect 298695 101167 298753 101201
rect 298787 101167 298816 101201
rect 298660 100949 298799 101167
rect 298660 100841 298661 100949
rect 298695 100807 298799 100915
rect 298660 100657 298799 100807
rect 298660 100623 298661 100657
rect 298695 100623 298753 100657
rect 298787 100623 298816 100657
rect 298660 100473 298799 100623
rect 298660 100331 298661 100439
rect 298695 100365 298799 100473
rect 298660 100113 298799 100331
rect 298660 100079 298661 100113
rect 298695 100079 298753 100113
rect 298787 100079 298816 100113
rect 298660 99861 298799 100079
rect 298660 99753 298661 99861
rect 298695 99719 298799 99827
rect 298660 99569 298799 99719
rect 298660 99535 298661 99569
rect 298695 99535 298753 99569
rect 298787 99535 298816 99569
rect 298660 99385 298799 99535
rect 298660 99243 298661 99351
rect 298695 99277 298799 99385
rect 298660 99025 298799 99243
rect 298660 98991 298661 99025
rect 298695 98991 298753 99025
rect 298787 98991 298816 99025
rect 298660 98773 298799 98991
rect 298660 98665 298661 98773
rect 298695 98631 298799 98739
rect 298660 98481 298799 98631
rect 298660 98447 298661 98481
rect 298695 98447 298753 98481
rect 298787 98447 298816 98481
rect 298660 98297 298799 98447
rect 298660 98155 298661 98263
rect 298695 98189 298799 98297
rect 298660 97937 298799 98155
rect 298660 97903 298661 97937
rect 298695 97903 298753 97937
rect 298787 97903 298816 97937
rect 298660 97685 298799 97903
rect 298660 97577 298661 97685
rect 298695 97543 298799 97651
rect 298660 97393 298799 97543
rect 298660 97359 298661 97393
rect 298695 97359 298753 97393
rect 298787 97359 298816 97393
rect 298660 97209 298799 97359
rect 298660 97067 298661 97175
rect 298695 97101 298799 97209
rect 298660 96849 298799 97067
rect 298660 96815 298661 96849
rect 298695 96815 298753 96849
rect 298787 96815 298816 96849
rect 298660 96597 298799 96815
rect 298660 96489 298661 96597
rect 298695 96455 298799 96563
rect 298660 96305 298799 96455
rect 298660 96271 298661 96305
rect 298695 96271 298753 96305
rect 298787 96271 298816 96305
rect 298660 96121 298799 96271
rect 298660 95979 298661 96087
rect 298695 96013 298799 96121
rect 298660 95761 298799 95979
rect 298660 95727 298661 95761
rect 298695 95727 298753 95761
rect 298787 95727 298816 95761
rect 298660 95509 298799 95727
rect 298660 95401 298661 95509
rect 298695 95367 298799 95475
rect 298660 95217 298799 95367
rect 298660 95183 298661 95217
rect 298695 95183 298753 95217
rect 298787 95183 298816 95217
rect 298660 95033 298799 95183
rect 298660 94891 298661 94999
rect 298695 94925 298799 95033
rect 298660 94673 298799 94891
rect 298660 94639 298661 94673
rect 298695 94639 298753 94673
rect 298787 94639 298816 94673
rect 298660 94421 298799 94639
rect 298660 94313 298661 94421
rect 298695 94279 298799 94387
rect 298660 94129 298799 94279
rect 298660 94095 298661 94129
rect 298695 94095 298753 94129
rect 298787 94095 298816 94129
rect 298660 93945 298799 94095
rect 298660 93803 298661 93911
rect 298695 93837 298799 93945
rect 298660 93585 298799 93803
rect 298660 93551 298661 93585
rect 298695 93551 298753 93585
rect 298787 93551 298816 93585
rect 298660 93333 298799 93551
rect 298660 93225 298661 93333
rect 298695 93191 298799 93299
rect 298660 93041 298799 93191
rect 298660 93007 298661 93041
rect 298695 93007 298753 93041
rect 298787 93007 298816 93041
rect 298660 92857 298799 93007
rect 298660 92715 298661 92823
rect 298695 92749 298799 92857
rect 298660 92497 298799 92715
rect 298660 92463 298661 92497
rect 298695 92463 298753 92497
rect 298787 92463 298816 92497
rect 298660 92245 298799 92463
rect 298660 92137 298661 92245
rect 298695 92103 298799 92211
rect 298660 91953 298799 92103
rect 298660 91919 298661 91953
rect 298695 91919 298753 91953
rect 298787 91919 298816 91953
rect 298660 91769 298799 91919
rect 298660 91627 298661 91735
rect 298695 91661 298799 91769
rect 298660 91409 298799 91627
rect 298660 91375 298661 91409
rect 298695 91375 298753 91409
rect 298787 91375 298816 91409
rect 298660 91157 298799 91375
rect 298660 91049 298661 91157
rect 298695 91015 298799 91123
rect 298660 90865 298799 91015
rect 298660 90831 298661 90865
rect 298695 90831 298753 90865
rect 298787 90831 298816 90865
rect 298660 90681 298799 90831
rect 298660 90539 298661 90647
rect 298695 90573 298799 90681
rect 298660 90321 298799 90539
rect 298660 90287 298661 90321
rect 298695 90287 298753 90321
rect 298787 90287 298816 90321
rect 298660 90069 298799 90287
rect 298660 89961 298661 90069
rect 298695 89927 298799 90035
rect 298660 89777 298799 89927
rect 298660 89743 298661 89777
rect 298695 89743 298753 89777
rect 298787 89743 298816 89777
rect 298660 89593 298799 89743
rect 298660 89451 298661 89559
rect 298695 89485 298799 89593
rect 298660 89233 298799 89451
rect 298660 89199 298661 89233
rect 298695 89199 298753 89233
rect 298787 89199 298816 89233
rect 298660 88981 298799 89199
rect 298660 88873 298661 88981
rect 298695 88839 298799 88947
rect 298660 88689 298799 88839
rect 298660 88655 298661 88689
rect 298695 88655 298753 88689
rect 298787 88655 298816 88689
rect 298660 88505 298799 88655
rect 298660 88363 298661 88471
rect 298695 88397 298799 88505
rect 298660 88145 298799 88363
rect 298660 88111 298661 88145
rect 298695 88111 298753 88145
rect 298787 88111 298816 88145
rect 298660 87893 298799 88111
rect 298660 87785 298661 87893
rect 298695 87751 298799 87859
rect 298660 87601 298799 87751
rect 298660 87567 298661 87601
rect 298695 87567 298753 87601
rect 298787 87567 298816 87601
rect 298660 87417 298799 87567
rect 298660 87275 298661 87383
rect 298695 87309 298799 87417
rect 298660 87057 298799 87275
rect 298660 87023 298661 87057
rect 298695 87023 298753 87057
rect 298787 87023 298816 87057
rect 298660 86805 298799 87023
rect 298660 86697 298661 86805
rect 298695 86663 298799 86771
rect 298660 86513 298799 86663
rect 298660 86479 298661 86513
rect 298695 86479 298753 86513
rect 298787 86479 298816 86513
rect 298660 86329 298799 86479
rect 298660 86187 298661 86295
rect 298695 86221 298799 86329
rect 298660 85969 298799 86187
rect 298660 85935 298661 85969
rect 298695 85935 298753 85969
rect 298787 85935 298816 85969
rect 298660 85717 298799 85935
rect 298660 85609 298661 85717
rect 298695 85575 298799 85683
rect 298660 85425 298799 85575
rect 298660 85391 298661 85425
rect 298695 85391 298753 85425
rect 298787 85391 298816 85425
rect 298660 85241 298799 85391
rect 298660 85099 298661 85207
rect 298695 85133 298799 85241
rect 298660 84881 298799 85099
rect 298660 84847 298661 84881
rect 298695 84847 298753 84881
rect 298787 84847 298816 84881
rect 298660 84629 298799 84847
rect 298660 84521 298661 84629
rect 298695 84487 298799 84595
rect 298660 84337 298799 84487
rect 298660 84303 298661 84337
rect 298695 84303 298753 84337
rect 298787 84303 298816 84337
rect 298660 84153 298799 84303
rect 298660 84011 298661 84119
rect 298695 84045 298799 84153
rect 298660 83793 298799 84011
rect 298660 83759 298661 83793
rect 298695 83759 298753 83793
rect 298787 83759 298816 83793
rect 298660 83541 298799 83759
rect 298660 83433 298661 83541
rect 298695 83399 298799 83507
rect 298660 83249 298799 83399
rect 298660 83215 298661 83249
rect 298695 83215 298753 83249
rect 298787 83215 298816 83249
rect 298660 83065 298799 83215
rect 298660 82923 298661 83031
rect 298695 82957 298799 83065
rect 298660 82705 298799 82923
rect 298660 82671 298661 82705
rect 298695 82671 298753 82705
rect 298787 82671 298816 82705
rect 298660 82453 298799 82671
rect 298660 82345 298661 82453
rect 298695 82311 298799 82419
rect 298660 82161 298799 82311
rect 298660 82127 298661 82161
rect 298695 82127 298753 82161
rect 298787 82127 298816 82161
rect 298660 81977 298799 82127
rect 298660 81835 298661 81943
rect 298695 81869 298799 81977
rect 298660 81617 298799 81835
rect 298660 81583 298661 81617
rect 298695 81583 298753 81617
rect 298787 81583 298816 81617
rect 298660 81365 298799 81583
rect 298660 81257 298661 81365
rect 298695 81223 298799 81331
rect 298660 81073 298799 81223
rect 298660 81039 298661 81073
rect 298695 81039 298753 81073
rect 298787 81039 298816 81073
rect 298660 80889 298799 81039
rect 298660 80747 298661 80855
rect 298695 80781 298799 80889
rect 298660 80529 298799 80747
rect 298660 80495 298661 80529
rect 298695 80495 298753 80529
rect 298787 80495 298816 80529
rect 298660 80277 298799 80495
rect 298660 80169 298661 80277
rect 298695 80135 298799 80243
rect 298660 79985 298799 80135
rect 298660 79951 298661 79985
rect 298695 79951 298753 79985
rect 298787 79951 298816 79985
rect 298660 79801 298799 79951
rect 298660 79659 298661 79767
rect 298695 79693 298799 79801
rect 298660 79441 298799 79659
rect 298660 79407 298661 79441
rect 298695 79407 298753 79441
rect 298787 79407 298816 79441
rect 298660 79189 298799 79407
rect 298660 79081 298661 79189
rect 298695 79047 298799 79155
rect 298660 78897 298799 79047
rect 298660 78863 298661 78897
rect 298695 78863 298753 78897
rect 298787 78863 298816 78897
rect 298660 78713 298799 78863
rect 298660 78571 298661 78679
rect 298695 78605 298799 78713
rect 298660 78353 298799 78571
rect 298660 78319 298661 78353
rect 298695 78319 298753 78353
rect 298787 78319 298816 78353
rect 298660 78101 298799 78319
rect 298660 77993 298661 78101
rect 298695 77959 298799 78067
rect 298660 77809 298799 77959
rect 298660 77775 298661 77809
rect 298695 77775 298753 77809
rect 298787 77775 298816 77809
rect 298660 77625 298799 77775
rect 298660 77483 298661 77591
rect 298695 77517 298799 77625
rect 298660 77265 298799 77483
rect 298660 77231 298661 77265
rect 298695 77231 298753 77265
rect 298787 77231 298816 77265
rect 298660 77013 298799 77231
rect 298660 76905 298661 77013
rect 298695 76871 298799 76979
rect 298660 76721 298799 76871
rect 298660 76687 298661 76721
rect 298695 76687 298753 76721
rect 298787 76687 298816 76721
rect 298660 76537 298799 76687
rect 298660 76395 298661 76503
rect 298695 76429 298799 76537
rect 298660 76177 298799 76395
rect 298660 76143 298661 76177
rect 298695 76143 298753 76177
rect 298787 76143 298816 76177
rect 298660 75925 298799 76143
rect 298660 75817 298661 75925
rect 298695 75783 298799 75891
rect 298660 75633 298799 75783
rect 298660 75599 298661 75633
rect 298695 75599 298753 75633
rect 298787 75599 298816 75633
rect 298660 75449 298799 75599
rect 298660 75307 298661 75415
rect 298695 75341 298799 75449
rect 298660 75089 298799 75307
rect 298660 75055 298661 75089
rect 298695 75055 298753 75089
rect 298787 75055 298816 75089
rect 298660 74837 298799 75055
rect 298660 74729 298661 74837
rect 298695 74695 298799 74803
rect 298660 74545 298799 74695
rect 298660 74511 298661 74545
rect 298695 74511 298753 74545
rect 298787 74511 298816 74545
rect 298660 74361 298799 74511
rect 298660 74219 298661 74327
rect 298695 74253 298799 74361
rect 298660 74001 298799 74219
rect 298660 73967 298661 74001
rect 298695 73967 298753 74001
rect 298787 73967 298816 74001
rect 298660 73749 298799 73967
rect 298660 73641 298661 73749
rect 298695 73607 298799 73715
rect 298660 73457 298799 73607
rect 298660 73423 298661 73457
rect 298695 73423 298753 73457
rect 298787 73423 298816 73457
rect 298660 73273 298799 73423
rect 298660 73131 298661 73239
rect 298695 73165 298799 73273
rect 298660 72913 298799 73131
rect 298660 72879 298661 72913
rect 298695 72879 298753 72913
rect 298787 72879 298816 72913
rect 298660 72661 298799 72879
rect 298660 72553 298661 72661
rect 298695 72519 298799 72627
rect 298660 72369 298799 72519
rect 298660 72335 298661 72369
rect 298695 72335 298753 72369
rect 298787 72335 298816 72369
rect 298660 72185 298799 72335
rect 298660 72043 298661 72151
rect 298695 72077 298799 72185
rect 298660 71825 298799 72043
rect 298660 71791 298661 71825
rect 298695 71791 298753 71825
rect 298787 71791 298816 71825
rect 298660 71573 298799 71791
rect 298660 71465 298661 71573
rect 298695 71431 298799 71539
rect 298660 71281 298799 71431
rect 298660 71247 298661 71281
rect 298695 71247 298753 71281
rect 298787 71247 298816 71281
rect 298660 71097 298799 71247
rect 298660 70955 298661 71063
rect 298695 70989 298799 71097
rect 298660 70737 298799 70955
rect 298660 70703 298661 70737
rect 298695 70703 298753 70737
rect 298787 70703 298816 70737
rect 298660 70485 298799 70703
rect 298660 70377 298661 70485
rect 298695 70343 298799 70451
rect 298660 70193 298799 70343
rect 298660 70159 298661 70193
rect 298695 70159 298753 70193
rect 298787 70159 298816 70193
rect 298660 70009 298799 70159
rect 298660 69867 298661 69975
rect 298695 69901 298799 70009
rect 298660 69649 298799 69867
rect 298660 69615 298661 69649
rect 298695 69615 298753 69649
rect 298787 69615 298816 69649
rect 298660 69397 298799 69615
rect 298660 69289 298661 69397
rect 298695 69255 298799 69363
rect 298660 69105 298799 69255
rect 298660 69071 298661 69105
rect 298695 69071 298753 69105
rect 298787 69071 298816 69105
rect 298660 68921 298799 69071
rect 298660 68779 298661 68887
rect 298695 68813 298799 68921
rect 298660 68561 298799 68779
rect 298660 68527 298661 68561
rect 298695 68527 298753 68561
rect 298787 68527 298816 68561
rect 298660 68309 298799 68527
rect 298660 68201 298661 68309
rect 298695 68167 298799 68275
rect 298660 68017 298799 68167
rect 298660 67983 298661 68017
rect 298695 67983 298753 68017
rect 298787 67983 298816 68017
rect 298660 67833 298799 67983
rect 298660 67691 298661 67799
rect 298695 67725 298799 67833
rect 298660 67473 298799 67691
rect 298660 67439 298661 67473
rect 298695 67439 298753 67473
rect 298787 67439 298816 67473
rect 298660 67221 298799 67439
rect 298660 67113 298661 67221
rect 298695 67079 298799 67187
rect 298660 66929 298799 67079
rect 298660 66895 298661 66929
rect 298695 66895 298753 66929
rect 298787 66895 298816 66929
rect 298660 66745 298799 66895
rect 298660 66603 298661 66711
rect 298695 66637 298799 66745
rect 298660 66385 298799 66603
rect 298660 66351 298661 66385
rect 298695 66351 298753 66385
rect 298787 66351 298816 66385
rect 298660 66133 298799 66351
rect 298660 66025 298661 66133
rect 298695 65991 298799 66099
rect 298660 65841 298799 65991
rect 298660 65807 298661 65841
rect 298695 65807 298753 65841
rect 298787 65807 298816 65841
rect 298660 65657 298799 65807
rect 298660 65515 298661 65623
rect 298695 65549 298799 65657
rect 298660 65297 298799 65515
rect 298660 65263 298661 65297
rect 298695 65263 298753 65297
rect 298787 65263 298816 65297
rect 298660 65045 298799 65263
rect 298660 64937 298661 65045
rect 298695 64903 298799 65011
rect 298660 64753 298799 64903
rect 298660 64719 298661 64753
rect 298695 64719 298753 64753
rect 298787 64719 298816 64753
rect 298660 64569 298799 64719
rect 298660 64427 298661 64535
rect 298695 64461 298799 64569
rect 298660 64209 298799 64427
rect 298660 64175 298661 64209
rect 298695 64175 298753 64209
rect 298787 64175 298816 64209
rect 298660 63957 298799 64175
rect 298660 63849 298661 63957
rect 298695 63815 298799 63923
rect 298660 63665 298799 63815
rect 298660 63631 298661 63665
rect 298695 63631 298753 63665
rect 298787 63631 298816 63665
rect 298660 63481 298799 63631
rect 298660 63339 298661 63447
rect 298695 63373 298799 63481
rect 298660 63121 298799 63339
rect 298660 63087 298661 63121
rect 298695 63087 298753 63121
rect 298787 63087 298816 63121
rect 298660 62869 298799 63087
rect 298660 62761 298661 62869
rect 298695 62727 298799 62835
rect 298660 62577 298799 62727
rect 298660 62543 298661 62577
rect 298695 62543 298753 62577
rect 298787 62543 298816 62577
rect 298660 62393 298799 62543
rect 298660 62251 298661 62359
rect 298695 62285 298799 62393
rect 298660 62033 298799 62251
rect 298660 61999 298661 62033
rect 298695 61999 298753 62033
rect 298787 61999 298816 62033
rect 298660 61781 298799 61999
rect 298660 61673 298661 61781
rect 298695 61639 298799 61747
rect 298660 61489 298799 61639
rect 298660 61455 298661 61489
rect 298695 61455 298753 61489
rect 298787 61455 298816 61489
rect 298660 61305 298799 61455
rect 298660 61163 298661 61271
rect 298695 61197 298799 61305
rect 298660 60945 298799 61163
rect 298660 60911 298661 60945
rect 298695 60911 298753 60945
rect 298787 60911 298816 60945
rect 298660 60693 298799 60911
rect 298660 60585 298661 60693
rect 298695 60551 298799 60659
rect 298660 60401 298799 60551
rect 298660 60367 298661 60401
rect 298695 60367 298753 60401
rect 298787 60367 298816 60401
rect 298660 60217 298799 60367
rect 298660 60075 298661 60183
rect 298695 60109 298799 60217
rect 298660 59857 298799 60075
rect 298660 59823 298661 59857
rect 298695 59823 298753 59857
rect 298787 59823 298816 59857
rect 298660 59605 298799 59823
rect 298660 59497 298661 59605
rect 298695 59463 298799 59571
rect 298660 59313 298799 59463
rect 298660 59279 298661 59313
rect 298695 59279 298753 59313
rect 298787 59279 298816 59313
rect 298660 59129 298799 59279
rect 298660 58987 298661 59095
rect 298695 59021 298799 59129
rect 298660 58769 298799 58987
rect 298660 58735 298661 58769
rect 298695 58735 298753 58769
rect 298787 58735 298816 58769
rect 298660 58517 298799 58735
rect 298660 58409 298661 58517
rect 298695 58375 298799 58483
rect 298660 58225 298799 58375
rect 298660 58191 298661 58225
rect 298695 58191 298753 58225
rect 298787 58191 298816 58225
rect 298660 58041 298799 58191
rect 298660 57899 298661 58007
rect 298695 57933 298799 58041
rect 298660 57681 298799 57899
rect 298660 57647 298661 57681
rect 298695 57647 298753 57681
rect 298787 57647 298816 57681
rect 298660 57429 298799 57647
rect 298660 57321 298661 57429
rect 298695 57287 298799 57395
rect 298660 57137 298799 57287
rect 298660 57103 298661 57137
rect 298695 57103 298753 57137
rect 298787 57103 298816 57137
rect 298660 56953 298799 57103
rect 298660 56811 298661 56919
rect 298695 56845 298799 56953
rect 298660 56593 298799 56811
rect 298660 56559 298661 56593
rect 298695 56559 298753 56593
rect 298787 56559 298816 56593
rect 298660 56341 298799 56559
rect 298660 56233 298661 56341
rect 298695 56199 298799 56307
rect 298660 56049 298799 56199
rect 298660 56015 298661 56049
rect 298695 56015 298753 56049
rect 298787 56015 298816 56049
rect 298660 55865 298799 56015
rect 298660 55723 298661 55831
rect 298695 55757 298799 55865
rect 298660 55505 298799 55723
rect 298660 55471 298661 55505
rect 298695 55471 298753 55505
rect 298787 55471 298816 55505
rect 298660 55253 298799 55471
rect 298660 55145 298661 55253
rect 298695 55111 298799 55219
rect 298660 54961 298799 55111
rect 298660 54927 298661 54961
rect 298695 54927 298753 54961
rect 298787 54927 298816 54961
rect 298660 54777 298799 54927
rect 298660 54635 298661 54743
rect 298695 54669 298799 54777
rect 298660 54417 298799 54635
rect 298660 54383 298661 54417
rect 298695 54383 298753 54417
rect 298787 54383 298816 54417
rect 298660 54165 298799 54383
rect 298660 54057 298661 54165
rect 298695 54023 298799 54131
rect 298660 53873 298799 54023
rect 298660 53839 298661 53873
rect 298695 53839 298753 53873
rect 298787 53839 298816 53873
rect 298660 53689 298799 53839
rect 298660 53547 298661 53655
rect 298695 53581 298799 53689
rect 298660 53329 298799 53547
rect 298660 53295 298661 53329
rect 298695 53295 298753 53329
rect 298787 53295 298816 53329
rect 298660 53077 298799 53295
rect 298660 52969 298661 53077
rect 298695 52935 298799 53043
rect 298660 52785 298799 52935
rect 298660 52751 298661 52785
rect 298695 52751 298753 52785
rect 298787 52751 298816 52785
rect 298660 52601 298799 52751
rect 298660 52459 298661 52567
rect 298695 52493 298799 52601
rect 298660 52241 298799 52459
rect 298660 52207 298661 52241
rect 298695 52207 298753 52241
rect 298787 52207 298816 52241
rect 298660 51989 298799 52207
rect 298660 51881 298661 51989
rect 298695 51847 298799 51955
rect 298660 51697 298799 51847
rect 298660 51663 298661 51697
rect 298695 51663 298753 51697
rect 298787 51663 298816 51697
rect 298660 51513 298799 51663
rect 298660 51371 298661 51479
rect 298695 51405 298799 51513
rect 298660 51153 298799 51371
rect 298660 51119 298661 51153
rect 298695 51119 298753 51153
rect 298787 51119 298816 51153
rect 298660 50901 298799 51119
rect 298660 50793 298661 50901
rect 298695 50759 298799 50867
rect 298660 50609 298799 50759
rect 298660 50575 298661 50609
rect 298695 50575 298753 50609
rect 298787 50575 298816 50609
rect 298660 50425 298799 50575
rect 298660 50283 298661 50391
rect 298695 50317 298799 50425
rect 298660 50065 298799 50283
rect 298660 50031 298661 50065
rect 298695 50031 298753 50065
rect 298787 50031 298816 50065
rect 298660 49813 298799 50031
rect 298660 49705 298661 49813
rect 298695 49671 298799 49779
rect 298660 49521 298799 49671
rect 298660 49487 298661 49521
rect 298695 49487 298753 49521
rect 298787 49487 298816 49521
rect 298660 49337 298799 49487
rect 298660 49195 298661 49303
rect 298695 49229 298799 49337
rect 298660 48977 298799 49195
rect 298660 48943 298661 48977
rect 298695 48943 298753 48977
rect 298787 48943 298816 48977
rect 298660 48725 298799 48943
rect 298660 48617 298661 48725
rect 298695 48583 298799 48691
rect 298660 48433 298799 48583
rect 298660 48399 298661 48433
rect 298695 48399 298753 48433
rect 298787 48399 298816 48433
rect 298660 48249 298799 48399
rect 298660 48107 298661 48215
rect 298695 48141 298799 48249
rect 298660 47889 298799 48107
rect 298660 47855 298661 47889
rect 298695 47855 298753 47889
rect 298787 47855 298816 47889
rect 298660 47637 298799 47855
rect 298660 47529 298661 47637
rect 298695 47495 298799 47603
rect 298660 47345 298799 47495
rect 298660 47311 298661 47345
rect 298695 47311 298753 47345
rect 298787 47311 298816 47345
rect 298660 47161 298799 47311
rect 298660 47019 298661 47127
rect 298695 47053 298799 47161
rect 298660 46801 298799 47019
rect 298660 46767 298661 46801
rect 298695 46767 298753 46801
rect 298787 46767 298816 46801
rect 298660 46549 298799 46767
rect 298660 46441 298661 46549
rect 298695 46407 298799 46515
rect 298660 46257 298799 46407
rect 298660 46223 298661 46257
rect 298695 46223 298753 46257
rect 298787 46223 298816 46257
rect 298660 46073 298799 46223
rect 298660 45931 298661 46039
rect 298695 45965 298799 46073
rect 298660 45713 298799 45931
rect 298660 45679 298661 45713
rect 298695 45679 298753 45713
rect 298787 45679 298816 45713
rect 298660 45461 298799 45679
rect 298660 45353 298661 45461
rect 298695 45319 298799 45427
rect 298660 45169 298799 45319
rect 298660 45135 298661 45169
rect 298695 45135 298753 45169
rect 298787 45135 298816 45169
rect 298660 44985 298799 45135
rect 298660 44843 298661 44951
rect 298695 44877 298799 44985
rect 298660 44625 298799 44843
rect 298660 44591 298661 44625
rect 298695 44591 298753 44625
rect 298787 44591 298816 44625
rect 298660 44373 298799 44591
rect 298660 44265 298661 44373
rect 298695 44231 298799 44339
rect 298660 44081 298799 44231
rect 298660 44047 298661 44081
rect 298695 44047 298753 44081
rect 298787 44047 298816 44081
rect 298660 43897 298799 44047
rect 298660 43755 298661 43863
rect 298695 43789 298799 43897
rect 298660 43537 298799 43755
rect 298660 43503 298661 43537
rect 298695 43503 298753 43537
rect 298787 43503 298816 43537
rect 298660 43285 298799 43503
rect 298660 43177 298661 43285
rect 298695 43143 298799 43251
rect 298660 42993 298799 43143
rect 298660 42959 298661 42993
rect 298695 42959 298753 42993
rect 298787 42959 298816 42993
rect 298660 42809 298799 42959
rect 298660 42667 298661 42775
rect 298695 42701 298799 42809
rect 298660 42449 298799 42667
rect 298660 42415 298661 42449
rect 298695 42415 298753 42449
rect 298787 42415 298816 42449
rect 298660 42197 298799 42415
rect 298660 42089 298661 42197
rect 298695 42055 298799 42163
rect 298660 41905 298799 42055
rect 298660 41871 298661 41905
rect 298695 41871 298753 41905
rect 298787 41871 298816 41905
rect 298660 41721 298799 41871
rect 298660 41579 298661 41687
rect 298695 41613 298799 41721
rect 298660 41361 298799 41579
rect 298660 41327 298661 41361
rect 298695 41327 298753 41361
rect 298787 41327 298816 41361
rect 298660 41109 298799 41327
rect 298660 41001 298661 41109
rect 298695 40967 298799 41075
rect 298660 40817 298799 40967
rect 298660 40783 298661 40817
rect 298695 40783 298753 40817
rect 298787 40783 298816 40817
rect 298660 40633 298799 40783
rect 298660 40491 298661 40599
rect 298695 40525 298799 40633
rect 298660 40273 298799 40491
rect 298660 40239 298661 40273
rect 298695 40239 298753 40273
rect 298787 40239 298816 40273
rect 298660 40021 298799 40239
rect 298660 39913 298661 40021
rect 298695 39879 298799 39987
rect 298660 39729 298799 39879
rect 298660 39695 298661 39729
rect 298695 39695 298753 39729
rect 298787 39695 298816 39729
rect 298660 39545 298799 39695
rect 298660 39403 298661 39511
rect 298695 39437 298799 39545
rect 298660 39185 298799 39403
rect 298660 39151 298661 39185
rect 298695 39151 298753 39185
rect 298787 39151 298816 39185
rect 298660 38933 298799 39151
rect 298660 38825 298661 38933
rect 298695 38791 298799 38899
rect 298660 38641 298799 38791
rect 298660 38607 298661 38641
rect 298695 38607 298753 38641
rect 298787 38607 298816 38641
rect 298660 38457 298799 38607
rect 298660 38315 298661 38423
rect 298695 38349 298799 38457
rect 298660 38097 298799 38315
rect 298660 38063 298661 38097
rect 298695 38063 298753 38097
rect 298787 38063 298816 38097
rect 298660 37845 298799 38063
rect 298660 37737 298661 37845
rect 298695 37703 298799 37811
rect 298660 37553 298799 37703
rect 298660 37519 298661 37553
rect 298695 37519 298753 37553
rect 298787 37519 298816 37553
rect 298660 37369 298799 37519
rect 298660 37227 298661 37335
rect 298695 37261 298799 37369
rect 298660 37009 298799 37227
rect 298660 36975 298661 37009
rect 298695 36975 298753 37009
rect 298787 36975 298816 37009
rect 298660 36757 298799 36975
rect 298660 36649 298661 36757
rect 298695 36615 298799 36723
rect 298660 36465 298799 36615
rect 298660 36431 298661 36465
rect 298695 36431 298753 36465
rect 298787 36431 298816 36465
rect 298660 36281 298799 36431
rect 298660 36139 298661 36247
rect 298695 36173 298799 36281
rect 298660 35921 298799 36139
rect 298660 35887 298661 35921
rect 298695 35887 298753 35921
rect 298787 35887 298816 35921
rect 298660 35669 298799 35887
rect 298660 35561 298661 35669
rect 298695 35527 298799 35635
rect 298660 35377 298799 35527
rect 298660 35343 298661 35377
rect 298695 35343 298753 35377
rect 298787 35343 298816 35377
rect 298660 35193 298799 35343
rect 298660 35051 298661 35159
rect 298695 35085 298799 35193
rect 298660 34833 298799 35051
rect 298660 34799 298661 34833
rect 298695 34799 298753 34833
rect 298787 34799 298816 34833
rect 298660 34581 298799 34799
rect 298660 34473 298661 34581
rect 298695 34439 298799 34547
rect 298660 34289 298799 34439
rect 298660 34255 298661 34289
rect 298695 34255 298753 34289
rect 298787 34255 298816 34289
rect 298660 34105 298799 34255
rect 298660 33963 298661 34071
rect 298695 33997 298799 34105
rect 298660 33745 298799 33963
rect 298660 33711 298661 33745
rect 298695 33711 298753 33745
rect 298787 33711 298816 33745
rect 298660 33493 298799 33711
rect 298660 33385 298661 33493
rect 298695 33351 298799 33459
rect 298660 33201 298799 33351
rect 298660 33167 298661 33201
rect 298695 33167 298753 33201
rect 298787 33167 298816 33201
rect 298660 33017 298799 33167
rect 298660 32875 298661 32983
rect 298695 32909 298799 33017
rect 298660 32657 298799 32875
rect 298660 32623 298661 32657
rect 298695 32623 298753 32657
rect 298787 32623 298816 32657
rect 298660 32405 298799 32623
rect 298660 32297 298661 32405
rect 298695 32263 298799 32371
rect 298660 32113 298799 32263
rect 298660 32079 298661 32113
rect 298695 32079 298753 32113
rect 298787 32079 298816 32113
rect 298660 31929 298799 32079
rect 298660 31787 298661 31895
rect 298695 31821 298799 31929
rect 298660 31569 298799 31787
rect 298660 31535 298661 31569
rect 298695 31535 298753 31569
rect 298787 31535 298816 31569
rect 298660 31317 298799 31535
rect 298660 31209 298661 31317
rect 298695 31175 298799 31283
rect 298660 31025 298799 31175
rect 298660 30991 298661 31025
rect 298695 30991 298753 31025
rect 298787 30991 298816 31025
rect 298660 30841 298799 30991
rect 298660 30699 298661 30807
rect 298695 30733 298799 30841
rect 298660 30481 298799 30699
rect 298660 30447 298661 30481
rect 298695 30447 298753 30481
rect 298787 30447 298816 30481
rect 298660 30229 298799 30447
rect 298660 30121 298661 30229
rect 298695 30087 298799 30195
rect 298660 29937 298799 30087
rect 298660 29903 298661 29937
rect 298695 29903 298753 29937
rect 298787 29903 298816 29937
rect 298660 29753 298799 29903
rect 298660 29611 298661 29719
rect 298695 29645 298799 29753
rect 298660 29393 298799 29611
rect 298660 29359 298661 29393
rect 298695 29359 298753 29393
rect 298787 29359 298816 29393
rect 298660 29141 298799 29359
rect 298660 29033 298661 29141
rect 298695 28999 298799 29107
rect 298660 28849 298799 28999
rect 298660 28815 298661 28849
rect 298695 28815 298753 28849
rect 298787 28815 298816 28849
rect 298660 28665 298799 28815
rect 298660 28523 298661 28631
rect 298695 28557 298799 28665
rect 298660 28305 298799 28523
rect 298660 28271 298661 28305
rect 298695 28271 298753 28305
rect 298787 28271 298816 28305
rect 298660 28053 298799 28271
rect 298660 27945 298661 28053
rect 298695 27911 298799 28019
rect 298660 27761 298799 27911
rect 298660 27727 298661 27761
rect 298695 27727 298753 27761
rect 298787 27727 298816 27761
rect 298660 27577 298799 27727
rect 298660 27435 298661 27543
rect 298695 27469 298799 27577
rect 298660 27217 298799 27435
rect 298660 27183 298661 27217
rect 298695 27183 298753 27217
rect 298787 27183 298816 27217
rect 298660 26965 298799 27183
rect 298660 26857 298661 26965
rect 298695 26823 298799 26931
rect 298660 26673 298799 26823
rect 298660 26639 298661 26673
rect 298695 26639 298753 26673
rect 298787 26639 298816 26673
rect 298660 26489 298799 26639
rect 298660 26347 298661 26455
rect 298695 26381 298799 26489
rect 298660 26129 298799 26347
rect 298660 26095 298661 26129
rect 298695 26095 298753 26129
rect 298787 26095 298816 26129
rect 298660 25877 298799 26095
rect 298660 25769 298661 25877
rect 298695 25735 298799 25843
rect 298660 25585 298799 25735
rect 298660 25551 298661 25585
rect 298695 25551 298753 25585
rect 298787 25551 298816 25585
rect 298660 25401 298799 25551
rect 298660 25259 298661 25367
rect 298695 25293 298799 25401
rect 298660 25041 298799 25259
rect 298660 25007 298661 25041
rect 298695 25007 298753 25041
rect 298787 25007 298816 25041
rect 298660 24789 298799 25007
rect 298660 24681 298661 24789
rect 298695 24647 298799 24755
rect 298660 24497 298799 24647
rect 298660 24463 298661 24497
rect 298695 24463 298753 24497
rect 298787 24463 298816 24497
rect 298660 24313 298799 24463
rect 298660 24171 298661 24279
rect 298695 24205 298799 24313
rect 298660 23953 298799 24171
rect 298660 23919 298661 23953
rect 298695 23919 298753 23953
rect 298787 23919 298816 23953
rect 298660 23701 298799 23919
rect 298660 23593 298661 23701
rect 298695 23559 298799 23667
rect 298660 23409 298799 23559
rect 298660 23375 298661 23409
rect 298695 23375 298753 23409
rect 298787 23375 298816 23409
rect 298660 23225 298799 23375
rect 298660 23083 298661 23191
rect 298695 23117 298799 23225
rect 298660 22865 298799 23083
rect 298660 22831 298661 22865
rect 298695 22831 298753 22865
rect 298787 22831 298816 22865
rect 298660 22613 298799 22831
rect 298660 22505 298661 22613
rect 298695 22471 298799 22579
rect 298660 22321 298799 22471
rect 298660 22287 298661 22321
rect 298695 22287 298753 22321
rect 298787 22287 298816 22321
rect 298660 22137 298799 22287
rect 298660 21995 298661 22103
rect 298695 22029 298799 22137
rect 298660 21777 298799 21995
rect 298660 21743 298661 21777
rect 298695 21743 298753 21777
rect 298787 21743 298816 21777
rect 298660 21525 298799 21743
rect 298660 21417 298661 21525
rect 298695 21383 298799 21491
rect 298660 21233 298799 21383
rect 298660 21199 298661 21233
rect 298695 21199 298753 21233
rect 298787 21199 298816 21233
rect 298660 21049 298799 21199
rect 298660 20907 298661 21015
rect 298695 20941 298799 21049
rect 298660 20689 298799 20907
rect 298660 20655 298661 20689
rect 298695 20655 298753 20689
rect 298787 20655 298816 20689
rect 298660 20437 298799 20655
rect 298660 20329 298661 20437
rect 298695 20295 298799 20403
rect 298660 20145 298799 20295
rect 298660 20111 298661 20145
rect 298695 20111 298753 20145
rect 298787 20111 298816 20145
rect 298660 19961 298799 20111
rect 298660 19819 298661 19927
rect 298695 19853 298799 19961
rect 298660 19601 298799 19819
rect 298660 19567 298661 19601
rect 298695 19567 298753 19601
rect 298787 19567 298816 19601
rect 298660 19349 298799 19567
rect 298660 19241 298661 19349
rect 298695 19207 298799 19315
rect 298660 19057 298799 19207
rect 298660 19023 298661 19057
rect 298695 19023 298753 19057
rect 298787 19023 298816 19057
rect 298660 18873 298799 19023
rect 298660 18731 298661 18839
rect 298695 18765 298799 18873
rect 298660 18513 298799 18731
rect 298660 18479 298661 18513
rect 298695 18479 298753 18513
rect 298787 18479 298816 18513
rect 298660 18261 298799 18479
rect 298660 18153 298661 18261
rect 298695 18119 298799 18227
rect 298660 17969 298799 18119
rect 298660 17935 298661 17969
rect 298695 17935 298753 17969
rect 298787 17935 298816 17969
rect 298660 17785 298799 17935
rect 298660 17643 298661 17751
rect 298695 17677 298799 17785
rect 298660 17425 298799 17643
rect 298660 17391 298661 17425
rect 298695 17391 298753 17425
rect 298787 17391 298816 17425
rect 298660 17173 298799 17391
rect 298660 17065 298661 17173
rect 298695 17031 298799 17139
rect 298660 16881 298799 17031
rect 298660 16847 298661 16881
rect 298695 16847 298753 16881
rect 298787 16847 298816 16881
rect 298660 16697 298799 16847
rect 298660 16555 298661 16663
rect 298695 16589 298799 16697
rect 298660 16337 298799 16555
rect 298660 16303 298661 16337
rect 298695 16303 298753 16337
rect 298787 16303 298816 16337
rect 298660 16085 298799 16303
rect 298660 15977 298661 16085
rect 298695 15943 298799 16051
rect 298660 15793 298799 15943
rect 298660 15759 298661 15793
rect 298695 15759 298753 15793
rect 298787 15759 298816 15793
rect 298660 15609 298799 15759
rect 298660 15467 298661 15575
rect 298695 15501 298799 15609
rect 298660 15249 298799 15467
rect 298660 15215 298661 15249
rect 298695 15215 298753 15249
rect 298787 15215 298816 15249
rect 298660 14997 298799 15215
rect 298660 14889 298661 14997
rect 298695 14855 298799 14963
rect 298660 14705 298799 14855
rect 298660 14671 298661 14705
rect 298695 14671 298753 14705
rect 298787 14671 298816 14705
rect 298660 14521 298799 14671
rect 298660 14379 298661 14487
rect 298695 14413 298799 14521
rect 298660 14161 298799 14379
rect 298660 14127 298661 14161
rect 298695 14127 298753 14161
rect 298787 14127 298816 14161
rect 298660 13909 298799 14127
rect 298660 13801 298661 13909
rect 298695 13767 298799 13875
rect 298660 13617 298799 13767
rect 298660 13583 298661 13617
rect 298695 13583 298753 13617
rect 298787 13583 298816 13617
rect 298660 13433 298799 13583
rect 298660 13291 298661 13399
rect 298695 13325 298799 13433
rect 298660 13073 298799 13291
rect 298660 13039 298661 13073
rect 298695 13039 298753 13073
rect 298787 13039 298816 13073
rect 298660 12821 298799 13039
rect 298660 12713 298661 12821
rect 298695 12679 298799 12787
rect 298660 12529 298799 12679
rect 298660 12495 298661 12529
rect 298695 12495 298753 12529
rect 298787 12495 298816 12529
rect 298660 12345 298799 12495
rect 298660 12203 298661 12311
rect 298695 12237 298799 12345
rect 298660 11985 298799 12203
rect 298660 11951 298661 11985
rect 298695 11951 298753 11985
rect 298787 11951 298816 11985
rect 298660 11733 298799 11951
rect 298660 11625 298661 11733
rect 298695 11591 298799 11699
rect 298660 11441 298799 11591
rect 298660 11407 298661 11441
rect 298695 11407 298753 11441
rect 298787 11407 298816 11441
rect 298660 11257 298799 11407
rect 298660 11115 298661 11223
rect 298695 11149 298799 11257
rect 298660 10897 298799 11115
rect 298660 10863 298661 10897
rect 298695 10863 298753 10897
rect 298787 10863 298816 10897
rect 298660 10645 298799 10863
rect 298660 10537 298661 10645
rect 298695 10503 298799 10611
rect 298660 10353 298799 10503
rect 298660 10319 298661 10353
rect 298695 10319 298753 10353
rect 298787 10319 298816 10353
rect 298660 10169 298799 10319
rect 298660 10027 298661 10135
rect 298695 10061 298799 10169
rect 298660 9809 298799 10027
rect 298660 9775 298661 9809
rect 298695 9775 298753 9809
rect 298787 9775 298816 9809
rect 298660 9557 298799 9775
rect 298660 9449 298661 9557
rect 298695 9415 298799 9523
rect 298660 9265 298799 9415
rect 298660 9231 298661 9265
rect 298695 9231 298753 9265
rect 298787 9231 298816 9265
rect 298660 9081 298799 9231
rect 298660 8939 298661 9047
rect 298695 8973 298799 9081
rect 298660 8721 298799 8939
rect 298660 8687 298661 8721
rect 298695 8687 298753 8721
rect 298787 8687 298816 8721
rect 298660 8469 298799 8687
rect 298660 8361 298661 8469
rect 298695 8327 298799 8435
rect 298660 8177 298799 8327
rect 298660 8143 298661 8177
rect 298695 8143 298753 8177
rect 298787 8143 298816 8177
rect 298660 7993 298799 8143
rect 298660 7851 298661 7959
rect 298695 7885 298799 7993
rect 298660 7633 298799 7851
rect 298660 7599 298661 7633
rect 298695 7599 298753 7633
rect 298787 7599 298816 7633
rect 298660 7381 298799 7599
rect 298660 7273 298661 7381
rect 298695 7239 298799 7347
rect 298660 7089 298799 7239
rect 298660 7055 298661 7089
rect 298695 7055 298753 7089
rect 298787 7055 298816 7089
rect 298660 6905 298799 7055
rect 298660 6763 298661 6871
rect 298695 6797 298799 6905
rect 298660 6545 298799 6763
rect 298660 6511 298661 6545
rect 298695 6511 298753 6545
rect 298787 6511 298816 6545
rect 298660 6293 298799 6511
rect 298660 6185 298661 6293
rect 298695 6151 298799 6259
rect 298660 6001 298799 6151
rect 298660 5967 298661 6001
rect 298695 5967 298753 6001
rect 298787 5967 298816 6001
rect 298660 5817 298799 5967
rect 298660 5675 298661 5783
rect 298695 5709 298799 5817
rect 298660 5457 298799 5675
rect 298660 5423 298661 5457
rect 298695 5423 298753 5457
rect 298787 5423 298816 5457
rect 298660 5205 298799 5423
rect 298660 5097 298661 5205
rect 298695 5063 298799 5171
rect 298660 4913 298799 5063
rect 298660 4879 298661 4913
rect 298695 4879 298753 4913
rect 298787 4879 298816 4913
rect 298660 4729 298799 4879
rect 298660 4587 298661 4695
rect 298695 4621 298799 4729
rect 298660 4369 298799 4587
rect 298660 4335 298661 4369
rect 298695 4335 298753 4369
rect 298787 4335 298816 4369
rect 298660 4117 298799 4335
rect 298660 4009 298661 4117
rect 298695 3975 298799 4083
rect 298660 3825 298799 3975
rect 298660 3791 298661 3825
rect 298695 3791 298753 3825
rect 298787 3791 298816 3825
rect 298660 3641 298799 3791
rect 298660 3499 298661 3607
rect 298695 3533 298799 3641
rect 298660 3281 298799 3499
rect 298660 3247 298661 3281
rect 298695 3247 298753 3281
rect 298787 3247 298816 3281
rect 298660 3029 298799 3247
rect 298660 2921 298661 3029
rect 298695 2887 298799 2995
rect 298660 2737 298799 2887
rect 298660 2703 298661 2737
rect 298695 2703 298753 2737
rect 298787 2703 298816 2737
rect 298660 2553 298799 2703
rect 298660 2411 298661 2519
rect 298695 2445 298799 2553
rect 298660 2193 298799 2411
rect 298660 2159 298661 2193
rect 298695 2159 298753 2193
rect 298787 2159 298816 2193
<< viali >>
rect 1133 297551 1167 297585
rect 1225 297551 1259 297585
rect 1317 297551 1340 297585
rect 1133 297007 1167 297041
rect 1225 297007 1259 297041
rect 1317 297007 1340 297041
rect 1133 296463 1167 296497
rect 1225 296463 1259 296497
rect 1317 296463 1340 296497
rect 1133 295919 1167 295953
rect 1225 295919 1259 295953
rect 1317 295919 1340 295953
rect 1133 295375 1167 295409
rect 1225 295375 1259 295409
rect 1317 295375 1340 295409
rect 1133 294831 1167 294865
rect 1225 294831 1259 294865
rect 1317 294831 1340 294865
rect 1133 294287 1167 294321
rect 1225 294287 1259 294321
rect 1317 294287 1340 294321
rect 1133 293743 1167 293777
rect 1225 293743 1259 293777
rect 1317 293743 1340 293777
rect 1133 293199 1167 293233
rect 1225 293199 1259 293233
rect 1317 293199 1340 293233
rect 1133 292655 1167 292689
rect 1225 292655 1259 292689
rect 1317 292655 1340 292689
rect 1133 292111 1167 292145
rect 1225 292111 1259 292145
rect 1317 292111 1340 292145
rect 1133 291567 1167 291601
rect 1225 291567 1259 291601
rect 1317 291567 1340 291601
rect 1133 291023 1167 291057
rect 1225 291023 1259 291057
rect 1317 291023 1340 291057
rect 1133 290479 1167 290513
rect 1225 290479 1259 290513
rect 1317 290479 1340 290513
rect 1133 289935 1167 289969
rect 1225 289935 1259 289969
rect 1317 289935 1340 289969
rect 1133 289391 1167 289425
rect 1225 289391 1259 289425
rect 1317 289391 1340 289425
rect 1133 288847 1167 288881
rect 1225 288847 1259 288881
rect 1317 288847 1340 288881
rect 1133 288303 1167 288337
rect 1225 288303 1259 288337
rect 1317 288303 1340 288337
rect 1133 287759 1167 287793
rect 1225 287759 1259 287793
rect 1317 287759 1340 287793
rect 1133 287215 1167 287249
rect 1225 287215 1259 287249
rect 1317 287215 1340 287249
rect 1133 286671 1167 286705
rect 1225 286671 1259 286705
rect 1317 286671 1340 286705
rect 1133 286127 1167 286161
rect 1225 286127 1259 286161
rect 1317 286127 1340 286161
rect 1133 285583 1167 285617
rect 1225 285583 1259 285617
rect 1317 285583 1340 285617
rect 1133 285039 1167 285073
rect 1225 285039 1259 285073
rect 1317 285039 1340 285073
rect 1133 284495 1167 284529
rect 1225 284495 1259 284529
rect 1317 284495 1340 284529
rect 1133 283951 1167 283985
rect 1225 283951 1259 283985
rect 1317 283951 1340 283985
rect 1133 283407 1167 283441
rect 1225 283407 1259 283441
rect 1317 283407 1340 283441
rect 1133 282863 1167 282897
rect 1225 282863 1259 282897
rect 1317 282863 1340 282897
rect 1133 282319 1167 282353
rect 1225 282319 1259 282353
rect 1317 282319 1340 282353
rect 1133 281775 1167 281809
rect 1225 281775 1259 281809
rect 1317 281775 1340 281809
rect 1133 281231 1167 281265
rect 1225 281231 1259 281265
rect 1317 281231 1340 281265
rect 1133 280687 1167 280721
rect 1225 280687 1259 280721
rect 1317 280687 1340 280721
rect 1133 280143 1167 280177
rect 1225 280143 1259 280177
rect 1317 280143 1340 280177
rect 1133 279599 1167 279633
rect 1225 279599 1259 279633
rect 1317 279599 1340 279633
rect 1133 279055 1167 279089
rect 1225 279055 1259 279089
rect 1317 279055 1340 279089
rect 1133 278511 1167 278545
rect 1225 278511 1259 278545
rect 1317 278511 1340 278545
rect 1133 277967 1167 278001
rect 1225 277967 1259 278001
rect 1317 277967 1340 278001
rect 1133 277423 1167 277457
rect 1225 277423 1259 277457
rect 1317 277423 1340 277457
rect 1133 276879 1167 276913
rect 1225 276879 1259 276913
rect 1317 276879 1340 276913
rect 1133 276335 1167 276369
rect 1225 276335 1259 276369
rect 1317 276335 1340 276369
rect 1133 275791 1167 275825
rect 1225 275791 1259 275825
rect 1317 275791 1340 275825
rect 1133 275247 1167 275281
rect 1225 275247 1259 275281
rect 1317 275247 1340 275281
rect 1133 274703 1167 274737
rect 1225 274703 1259 274737
rect 1317 274703 1340 274737
rect 1133 274159 1167 274193
rect 1225 274159 1259 274193
rect 1317 274159 1340 274193
rect 1133 273615 1167 273649
rect 1225 273615 1259 273649
rect 1317 273615 1340 273649
rect 1133 273071 1167 273105
rect 1225 273071 1259 273105
rect 1317 273071 1340 273105
rect 1133 272527 1167 272561
rect 1225 272527 1259 272561
rect 1317 272527 1340 272561
rect 1133 271983 1167 272017
rect 1225 271983 1259 272017
rect 1317 271983 1340 272017
rect 1133 271439 1167 271473
rect 1225 271439 1259 271473
rect 1317 271439 1340 271473
rect 1133 270895 1167 270929
rect 1225 270895 1259 270929
rect 1317 270895 1340 270929
rect 1133 270351 1167 270385
rect 1225 270351 1259 270385
rect 1317 270351 1340 270385
rect 1133 269807 1167 269841
rect 1225 269807 1259 269841
rect 1317 269807 1340 269841
rect 1133 269263 1167 269297
rect 1225 269263 1259 269297
rect 1317 269263 1340 269297
rect 1133 268719 1167 268753
rect 1225 268719 1259 268753
rect 1317 268719 1340 268753
rect 1133 268175 1167 268209
rect 1225 268175 1259 268209
rect 1317 268175 1340 268209
rect 1133 267631 1167 267665
rect 1225 267631 1259 267665
rect 1317 267631 1340 267665
rect 1133 267087 1167 267121
rect 1225 267087 1259 267121
rect 1317 267087 1340 267121
rect 1133 266543 1167 266577
rect 1225 266543 1259 266577
rect 1317 266543 1340 266577
rect 1133 265999 1167 266033
rect 1225 265999 1259 266033
rect 1317 265999 1340 266033
rect 1133 265455 1167 265489
rect 1225 265455 1259 265489
rect 1317 265455 1340 265489
rect 1133 264911 1167 264945
rect 1225 264911 1259 264945
rect 1317 264911 1340 264945
rect 1133 264367 1167 264401
rect 1225 264367 1259 264401
rect 1317 264367 1340 264401
rect 1133 263823 1167 263857
rect 1225 263823 1259 263857
rect 1317 263823 1340 263857
rect 1133 263279 1167 263313
rect 1225 263279 1259 263313
rect 1317 263279 1340 263313
rect 1133 262735 1167 262769
rect 1225 262735 1259 262769
rect 1317 262735 1340 262769
rect 1133 262191 1167 262225
rect 1225 262191 1259 262225
rect 1317 262191 1340 262225
rect 1133 261647 1167 261681
rect 1225 261647 1259 261681
rect 1317 261647 1340 261681
rect 1133 261103 1167 261137
rect 1225 261103 1259 261137
rect 1317 261103 1340 261137
rect 1133 260559 1167 260593
rect 1225 260559 1259 260593
rect 1317 260559 1340 260593
rect 1133 260015 1167 260049
rect 1225 260015 1259 260049
rect 1317 260015 1340 260049
rect 1133 259471 1167 259505
rect 1225 259471 1259 259505
rect 1317 259471 1340 259505
rect 1133 258927 1167 258961
rect 1225 258927 1259 258961
rect 1317 258927 1340 258961
rect 1133 258383 1167 258417
rect 1225 258383 1259 258417
rect 1317 258383 1340 258417
rect 1133 257839 1167 257873
rect 1225 257839 1259 257873
rect 1317 257839 1340 257873
rect 1133 257295 1167 257329
rect 1225 257295 1259 257329
rect 1317 257295 1340 257329
rect 1133 256751 1167 256785
rect 1225 256751 1259 256785
rect 1317 256751 1340 256785
rect 1133 256207 1167 256241
rect 1225 256207 1259 256241
rect 1317 256207 1340 256241
rect 1133 255663 1167 255697
rect 1225 255663 1259 255697
rect 1317 255663 1340 255697
rect 1133 255119 1167 255153
rect 1225 255119 1259 255153
rect 1317 255119 1340 255153
rect 1133 254575 1167 254609
rect 1225 254575 1259 254609
rect 1317 254575 1340 254609
rect 1133 254031 1167 254065
rect 1225 254031 1259 254065
rect 1317 254031 1340 254065
rect 1133 253487 1167 253521
rect 1225 253487 1259 253521
rect 1317 253487 1340 253521
rect 1133 252943 1167 252977
rect 1225 252943 1259 252977
rect 1317 252943 1340 252977
rect 1133 252399 1167 252433
rect 1225 252399 1259 252433
rect 1317 252399 1340 252433
rect 1133 251855 1167 251889
rect 1225 251855 1259 251889
rect 1317 251855 1340 251889
rect 1133 251311 1167 251345
rect 1225 251311 1259 251345
rect 1317 251311 1340 251345
rect 1133 250767 1167 250801
rect 1225 250767 1259 250801
rect 1317 250767 1340 250801
rect 1133 250223 1167 250257
rect 1225 250223 1259 250257
rect 1317 250223 1340 250257
rect 1133 249679 1167 249713
rect 1225 249679 1259 249713
rect 1317 249679 1340 249713
rect 1133 249135 1167 249169
rect 1225 249135 1259 249169
rect 1317 249135 1340 249169
rect 1133 248591 1167 248625
rect 1225 248591 1259 248625
rect 1317 248591 1340 248625
rect 1133 248047 1167 248081
rect 1225 248047 1259 248081
rect 1317 248047 1340 248081
rect 1133 247503 1167 247537
rect 1225 247503 1259 247537
rect 1317 247503 1340 247537
rect 1133 246959 1167 246993
rect 1225 246959 1259 246993
rect 1317 246959 1340 246993
rect 1133 246415 1167 246449
rect 1225 246415 1259 246449
rect 1317 246415 1340 246449
rect 1133 245871 1167 245905
rect 1225 245871 1259 245905
rect 1317 245871 1340 245905
rect 1133 245327 1167 245361
rect 1225 245327 1259 245361
rect 1317 245327 1340 245361
rect 1133 244783 1167 244817
rect 1225 244783 1259 244817
rect 1317 244783 1340 244817
rect 1133 244239 1167 244273
rect 1225 244239 1259 244273
rect 1317 244239 1340 244273
rect 1133 243695 1167 243729
rect 1225 243695 1259 243729
rect 1317 243695 1340 243729
rect 1133 243151 1167 243185
rect 1225 243151 1259 243185
rect 1317 243151 1340 243185
rect 1133 242607 1167 242641
rect 1225 242607 1259 242641
rect 1317 242607 1340 242641
rect 1133 242063 1167 242097
rect 1225 242063 1259 242097
rect 1317 242063 1340 242097
rect 1133 241519 1167 241553
rect 1225 241519 1259 241553
rect 1317 241519 1340 241553
rect 1133 240975 1167 241009
rect 1225 240975 1259 241009
rect 1317 240975 1340 241009
rect 1133 240431 1167 240465
rect 1225 240431 1259 240465
rect 1317 240431 1340 240465
rect 1133 239887 1167 239921
rect 1225 239887 1259 239921
rect 1317 239887 1340 239921
rect 1133 239343 1167 239377
rect 1225 239343 1259 239377
rect 1317 239343 1340 239377
rect 1133 238799 1167 238833
rect 1225 238799 1259 238833
rect 1317 238799 1340 238833
rect 1133 238255 1167 238289
rect 1225 238255 1259 238289
rect 1317 238255 1340 238289
rect 1133 237711 1167 237745
rect 1225 237711 1259 237745
rect 1317 237711 1340 237745
rect 1133 237167 1167 237201
rect 1225 237167 1259 237201
rect 1317 237167 1340 237201
rect 1133 236623 1167 236657
rect 1225 236623 1259 236657
rect 1317 236623 1340 236657
rect 1133 236079 1167 236113
rect 1225 236079 1259 236113
rect 1317 236079 1340 236113
rect 1133 235535 1167 235569
rect 1225 235535 1259 235569
rect 1317 235535 1340 235569
rect 1133 234991 1167 235025
rect 1225 234991 1259 235025
rect 1317 234991 1340 235025
rect 1133 234447 1167 234481
rect 1225 234447 1259 234481
rect 1317 234447 1340 234481
rect 1133 233903 1167 233937
rect 1225 233903 1259 233937
rect 1317 233903 1340 233937
rect 1133 233359 1167 233393
rect 1225 233359 1259 233393
rect 1317 233359 1340 233393
rect 1133 232815 1167 232849
rect 1225 232815 1259 232849
rect 1317 232815 1340 232849
rect 1133 232271 1167 232305
rect 1225 232271 1259 232305
rect 1317 232271 1340 232305
rect 1133 231727 1167 231761
rect 1225 231727 1259 231761
rect 1317 231727 1340 231761
rect 1133 231183 1167 231217
rect 1225 231183 1259 231217
rect 1317 231183 1340 231217
rect 1133 230639 1167 230673
rect 1225 230639 1259 230673
rect 1317 230639 1340 230673
rect 1133 230095 1167 230129
rect 1225 230095 1259 230129
rect 1317 230095 1340 230129
rect 1133 229551 1167 229585
rect 1225 229551 1259 229585
rect 1317 229551 1340 229585
rect 1133 229007 1167 229041
rect 1225 229007 1259 229041
rect 1317 229007 1340 229041
rect 1133 228463 1167 228497
rect 1225 228463 1259 228497
rect 1317 228463 1340 228497
rect 1133 227919 1167 227953
rect 1225 227919 1259 227953
rect 1317 227919 1340 227953
rect 1133 227375 1167 227409
rect 1225 227375 1259 227409
rect 1317 227375 1340 227409
rect 1133 226831 1167 226865
rect 1225 226831 1259 226865
rect 1317 226831 1340 226865
rect 1133 226287 1167 226321
rect 1225 226287 1259 226321
rect 1317 226287 1340 226321
rect 1133 225743 1167 225777
rect 1225 225743 1259 225777
rect 1317 225743 1340 225777
rect 1133 225199 1167 225233
rect 1225 225199 1259 225233
rect 1317 225199 1340 225233
rect 1133 224655 1167 224689
rect 1225 224655 1259 224689
rect 1317 224655 1340 224689
rect 1133 224111 1167 224145
rect 1225 224111 1259 224145
rect 1317 224111 1340 224145
rect 1133 223567 1167 223601
rect 1225 223567 1259 223601
rect 1317 223567 1340 223601
rect 1133 223023 1167 223057
rect 1225 223023 1259 223057
rect 1317 223023 1340 223057
rect 1133 222479 1167 222513
rect 1225 222479 1259 222513
rect 1317 222479 1340 222513
rect 1133 221935 1167 221969
rect 1225 221935 1259 221969
rect 1317 221935 1340 221969
rect 1133 221391 1167 221425
rect 1225 221391 1259 221425
rect 1317 221391 1340 221425
rect 1133 220847 1167 220881
rect 1225 220847 1259 220881
rect 1317 220847 1340 220881
rect 1133 220303 1167 220337
rect 1225 220303 1259 220337
rect 1317 220303 1340 220337
rect 1133 219759 1167 219793
rect 1225 219759 1259 219793
rect 1317 219759 1340 219793
rect 1133 219215 1167 219249
rect 1225 219215 1259 219249
rect 1317 219215 1340 219249
rect 1133 218671 1167 218705
rect 1225 218671 1259 218705
rect 1317 218671 1340 218705
rect 1133 218127 1167 218161
rect 1225 218127 1259 218161
rect 1317 218127 1340 218161
rect 1133 217583 1167 217617
rect 1225 217583 1259 217617
rect 1317 217583 1340 217617
rect 1133 217039 1167 217073
rect 1225 217039 1259 217073
rect 1317 217039 1340 217073
rect 1133 216495 1167 216529
rect 1225 216495 1259 216529
rect 1317 216495 1340 216529
rect 1133 215951 1167 215985
rect 1225 215951 1259 215985
rect 1317 215951 1340 215985
rect 1133 215407 1167 215441
rect 1225 215407 1259 215441
rect 1317 215407 1340 215441
rect 1133 214863 1167 214897
rect 1225 214863 1259 214897
rect 1317 214863 1340 214897
rect 1133 214319 1167 214353
rect 1225 214319 1259 214353
rect 1317 214319 1340 214353
rect 1133 213775 1167 213809
rect 1225 213775 1259 213809
rect 1317 213775 1340 213809
rect 1133 213231 1167 213265
rect 1225 213231 1259 213265
rect 1317 213231 1340 213265
rect 1133 212687 1167 212721
rect 1225 212687 1259 212721
rect 1317 212687 1340 212721
rect 1133 212143 1167 212177
rect 1225 212143 1259 212177
rect 1317 212143 1340 212177
rect 1133 211599 1167 211633
rect 1225 211599 1259 211633
rect 1317 211599 1340 211633
rect 1133 211055 1167 211089
rect 1225 211055 1259 211089
rect 1317 211055 1340 211089
rect 1133 210511 1167 210545
rect 1225 210511 1259 210545
rect 1317 210511 1340 210545
rect 1133 209967 1167 210001
rect 1225 209967 1259 210001
rect 1317 209967 1340 210001
rect 1133 209423 1167 209457
rect 1225 209423 1259 209457
rect 1317 209423 1340 209457
rect 1133 208879 1167 208913
rect 1225 208879 1259 208913
rect 1317 208879 1340 208913
rect 1133 208335 1167 208369
rect 1225 208335 1259 208369
rect 1317 208335 1340 208369
rect 1133 207791 1167 207825
rect 1225 207791 1259 207825
rect 1317 207791 1340 207825
rect 1133 207247 1167 207281
rect 1225 207247 1259 207281
rect 1317 207247 1340 207281
rect 1133 206703 1167 206737
rect 1225 206703 1259 206737
rect 1317 206703 1340 206737
rect 1133 206159 1167 206193
rect 1225 206159 1259 206193
rect 1317 206159 1340 206193
rect 1133 205615 1167 205649
rect 1225 205615 1259 205649
rect 1317 205615 1340 205649
rect 1133 205071 1167 205105
rect 1225 205071 1259 205105
rect 1317 205071 1340 205105
rect 1133 204527 1167 204561
rect 1225 204527 1259 204561
rect 1317 204527 1340 204561
rect 1133 203983 1167 204017
rect 1225 203983 1259 204017
rect 1317 203983 1340 204017
rect 1133 203439 1167 203473
rect 1225 203439 1259 203473
rect 1317 203439 1340 203473
rect 1133 202895 1167 202929
rect 1225 202895 1259 202929
rect 1317 202895 1340 202929
rect 1133 202351 1167 202385
rect 1225 202351 1259 202385
rect 1317 202351 1340 202385
rect 1133 201807 1167 201841
rect 1225 201807 1259 201841
rect 1317 201807 1340 201841
rect 1133 201263 1167 201297
rect 1225 201263 1259 201297
rect 1317 201263 1340 201297
rect 1133 200719 1167 200753
rect 1225 200719 1259 200753
rect 1317 200719 1340 200753
rect 1133 200175 1167 200209
rect 1225 200175 1259 200209
rect 1317 200175 1340 200209
rect 1133 199631 1167 199665
rect 1225 199631 1259 199665
rect 1317 199631 1340 199665
rect 1133 199087 1167 199121
rect 1225 199087 1259 199121
rect 1317 199087 1340 199121
rect 1133 198543 1167 198577
rect 1225 198543 1259 198577
rect 1317 198543 1340 198577
rect 1133 197999 1167 198033
rect 1225 197999 1259 198033
rect 1317 197999 1340 198033
rect 1133 197455 1167 197489
rect 1225 197455 1259 197489
rect 1317 197455 1340 197489
rect 1133 196911 1167 196945
rect 1225 196911 1259 196945
rect 1317 196911 1340 196945
rect 1133 196367 1167 196401
rect 1225 196367 1259 196401
rect 1317 196367 1340 196401
rect 1133 195823 1167 195857
rect 1225 195823 1259 195857
rect 1317 195823 1340 195857
rect 1133 195279 1167 195313
rect 1225 195279 1259 195313
rect 1317 195279 1340 195313
rect 1133 194735 1167 194769
rect 1225 194735 1259 194769
rect 1317 194735 1340 194769
rect 1133 194191 1167 194225
rect 1225 194191 1259 194225
rect 1317 194191 1340 194225
rect 1133 193647 1167 193681
rect 1225 193647 1259 193681
rect 1317 193647 1340 193681
rect 1133 193103 1167 193137
rect 1225 193103 1259 193137
rect 1317 193103 1340 193137
rect 1133 192559 1167 192593
rect 1225 192559 1259 192593
rect 1317 192559 1340 192593
rect 1133 192015 1167 192049
rect 1225 192015 1259 192049
rect 1317 192015 1340 192049
rect 1133 191471 1167 191505
rect 1225 191471 1259 191505
rect 1317 191471 1340 191505
rect 1133 190927 1167 190961
rect 1225 190927 1259 190961
rect 1317 190927 1340 190961
rect 1133 190383 1167 190417
rect 1225 190383 1259 190417
rect 1317 190383 1340 190417
rect 1133 189839 1167 189873
rect 1225 189839 1259 189873
rect 1317 189839 1340 189873
rect 1133 189295 1167 189329
rect 1225 189295 1259 189329
rect 1317 189295 1340 189329
rect 1133 188751 1167 188785
rect 1225 188751 1259 188785
rect 1317 188751 1340 188785
rect 1133 188207 1167 188241
rect 1225 188207 1259 188241
rect 1317 188207 1340 188241
rect 1133 187663 1167 187697
rect 1225 187663 1259 187697
rect 1317 187663 1340 187697
rect 1133 187119 1167 187153
rect 1225 187119 1259 187153
rect 1317 187119 1340 187153
rect 1133 186575 1167 186609
rect 1225 186575 1259 186609
rect 1317 186575 1340 186609
rect 1133 186031 1167 186065
rect 1225 186031 1259 186065
rect 1317 186031 1340 186065
rect 1133 185487 1167 185521
rect 1225 185487 1259 185521
rect 1317 185487 1340 185521
rect 1133 184943 1167 184977
rect 1225 184943 1259 184977
rect 1317 184943 1340 184977
rect 1133 184399 1167 184433
rect 1225 184399 1259 184433
rect 1317 184399 1340 184433
rect 1133 183855 1167 183889
rect 1225 183855 1259 183889
rect 1317 183855 1340 183889
rect 1133 183311 1167 183345
rect 1225 183311 1259 183345
rect 1317 183311 1340 183345
rect 1133 182767 1167 182801
rect 1225 182767 1259 182801
rect 1317 182767 1340 182801
rect 1133 182223 1167 182257
rect 1225 182223 1259 182257
rect 1317 182223 1340 182257
rect 1133 181679 1167 181713
rect 1225 181679 1259 181713
rect 1317 181679 1340 181713
rect 1133 181135 1167 181169
rect 1225 181135 1259 181169
rect 1317 181135 1340 181169
rect 1133 180591 1167 180625
rect 1225 180591 1259 180625
rect 1317 180591 1340 180625
rect 1133 180047 1167 180081
rect 1225 180047 1259 180081
rect 1317 180047 1340 180081
rect 1133 179503 1167 179537
rect 1225 179503 1259 179537
rect 1317 179503 1340 179537
rect 1133 178959 1167 178993
rect 1225 178959 1259 178993
rect 1317 178959 1340 178993
rect 1133 178415 1167 178449
rect 1225 178415 1259 178449
rect 1317 178415 1340 178449
rect 1133 177871 1167 177905
rect 1225 177871 1259 177905
rect 1317 177871 1340 177905
rect 1133 177327 1167 177361
rect 1225 177327 1259 177361
rect 1317 177327 1340 177361
rect 1133 176783 1167 176817
rect 1225 176783 1259 176817
rect 1317 176783 1340 176817
rect 1133 176239 1167 176273
rect 1225 176239 1259 176273
rect 1317 176239 1340 176273
rect 1133 175695 1167 175729
rect 1225 175695 1259 175729
rect 1317 175695 1340 175729
rect 1133 175151 1167 175185
rect 1225 175151 1259 175185
rect 1317 175151 1340 175185
rect 1133 174607 1167 174641
rect 1225 174607 1259 174641
rect 1317 174607 1340 174641
rect 1133 174063 1167 174097
rect 1225 174063 1259 174097
rect 1317 174063 1340 174097
rect 1133 173519 1167 173553
rect 1225 173519 1259 173553
rect 1317 173519 1340 173553
rect 1133 172975 1167 173009
rect 1225 172975 1259 173009
rect 1317 172975 1340 173009
rect 1133 172431 1167 172465
rect 1225 172431 1259 172465
rect 1317 172431 1340 172465
rect 1133 171887 1167 171921
rect 1225 171887 1259 171921
rect 1317 171887 1340 171921
rect 1133 171343 1167 171377
rect 1225 171343 1259 171377
rect 1317 171343 1340 171377
rect 1133 170799 1167 170833
rect 1225 170799 1259 170833
rect 1317 170799 1340 170833
rect 1133 170255 1167 170289
rect 1225 170255 1259 170289
rect 1317 170255 1340 170289
rect 1133 169711 1167 169745
rect 1225 169711 1259 169745
rect 1317 169711 1340 169745
rect 1133 169167 1167 169201
rect 1225 169167 1259 169201
rect 1317 169167 1340 169201
rect 1133 168623 1167 168657
rect 1225 168623 1259 168657
rect 1317 168623 1340 168657
rect 1133 168079 1167 168113
rect 1225 168079 1259 168113
rect 1317 168079 1340 168113
rect 1133 167535 1167 167569
rect 1225 167535 1259 167569
rect 1317 167535 1340 167569
rect 1133 166991 1167 167025
rect 1225 166991 1259 167025
rect 1317 166991 1340 167025
rect 1133 166447 1167 166481
rect 1225 166447 1259 166481
rect 1317 166447 1340 166481
rect 1133 165903 1167 165937
rect 1225 165903 1259 165937
rect 1317 165903 1340 165937
rect 1133 165359 1167 165393
rect 1225 165359 1259 165393
rect 1317 165359 1340 165393
rect 1133 164815 1167 164849
rect 1225 164815 1259 164849
rect 1317 164815 1340 164849
rect 1133 164271 1167 164305
rect 1225 164271 1259 164305
rect 1317 164271 1340 164305
rect 1133 163727 1167 163761
rect 1225 163727 1259 163761
rect 1317 163727 1340 163761
rect 1133 163183 1167 163217
rect 1225 163183 1259 163217
rect 1317 163183 1340 163217
rect 1133 162639 1167 162673
rect 1225 162639 1259 162673
rect 1317 162639 1340 162673
rect 1133 162095 1167 162129
rect 1225 162095 1259 162129
rect 1317 162095 1340 162129
rect 1133 161551 1167 161585
rect 1225 161551 1259 161585
rect 1317 161551 1340 161585
rect 1133 161007 1167 161041
rect 1225 161007 1259 161041
rect 1317 161007 1340 161041
rect 1133 160463 1167 160497
rect 1225 160463 1259 160497
rect 1317 160463 1340 160497
rect 1133 159919 1167 159953
rect 1225 159919 1259 159953
rect 1317 159919 1340 159953
rect 1133 159375 1167 159409
rect 1225 159375 1259 159409
rect 1317 159375 1340 159409
rect 1133 158831 1167 158865
rect 1225 158831 1259 158865
rect 1317 158831 1340 158865
rect 1133 158287 1167 158321
rect 1225 158287 1259 158321
rect 1317 158287 1340 158321
rect 1133 157743 1167 157777
rect 1225 157743 1259 157777
rect 1317 157743 1340 157777
rect 1133 157199 1167 157233
rect 1225 157199 1259 157233
rect 1317 157199 1340 157233
rect 1133 156655 1167 156689
rect 1225 156655 1259 156689
rect 1317 156655 1340 156689
rect 1133 156111 1167 156145
rect 1225 156111 1259 156145
rect 1317 156111 1340 156145
rect 1133 155567 1167 155601
rect 1225 155567 1259 155601
rect 1317 155567 1340 155601
rect 1133 155023 1167 155057
rect 1225 155023 1259 155057
rect 1317 155023 1340 155057
rect 1133 154479 1167 154513
rect 1225 154479 1259 154513
rect 1317 154479 1340 154513
rect 1133 153935 1167 153969
rect 1225 153935 1259 153969
rect 1317 153935 1340 153969
rect 1133 153391 1167 153425
rect 1225 153391 1259 153425
rect 1317 153391 1340 153425
rect 1133 152847 1167 152881
rect 1225 152847 1259 152881
rect 1317 152847 1340 152881
rect 1133 152303 1167 152337
rect 1225 152303 1259 152337
rect 1317 152303 1340 152337
rect 1133 151759 1167 151793
rect 1225 151759 1259 151793
rect 1317 151759 1340 151793
rect 1133 151215 1167 151249
rect 1225 151215 1259 151249
rect 1317 151215 1340 151249
rect 1133 150671 1167 150705
rect 1225 150671 1259 150705
rect 1317 150671 1340 150705
rect 1133 150127 1167 150161
rect 1225 150127 1259 150161
rect 1317 150127 1340 150161
rect 1133 149583 1167 149617
rect 1225 149583 1259 149617
rect 1317 149583 1340 149617
rect 1133 149039 1167 149073
rect 1225 149039 1259 149073
rect 1317 149039 1340 149073
rect 1133 148495 1167 148529
rect 1225 148495 1259 148529
rect 1317 148495 1340 148529
rect 1133 147951 1167 147985
rect 1225 147951 1259 147985
rect 1317 147951 1340 147985
rect 1133 147407 1167 147441
rect 1225 147407 1259 147441
rect 1317 147407 1340 147441
rect 1133 146863 1167 146897
rect 1225 146863 1259 146897
rect 1317 146863 1340 146897
rect 1133 146319 1167 146353
rect 1225 146319 1259 146353
rect 1317 146319 1340 146353
rect 1133 145775 1167 145809
rect 1225 145775 1259 145809
rect 1317 145775 1340 145809
rect 1133 145231 1167 145265
rect 1225 145231 1259 145265
rect 1317 145231 1340 145265
rect 1133 144687 1167 144721
rect 1225 144687 1259 144721
rect 1317 144687 1340 144721
rect 1133 144143 1167 144177
rect 1225 144143 1259 144177
rect 1317 144143 1340 144177
rect 1133 143599 1167 143633
rect 1225 143599 1259 143633
rect 1317 143599 1340 143633
rect 1133 143055 1167 143089
rect 1225 143055 1259 143089
rect 1317 143055 1340 143089
rect 1133 142511 1167 142545
rect 1225 142511 1259 142545
rect 1317 142511 1340 142545
rect 1133 141967 1167 142001
rect 1225 141967 1259 142001
rect 1317 141967 1340 142001
rect 1133 141423 1167 141457
rect 1225 141423 1259 141457
rect 1317 141423 1340 141457
rect 1133 140879 1167 140913
rect 1225 140879 1259 140913
rect 1317 140879 1340 140913
rect 1133 140335 1167 140369
rect 1225 140335 1259 140369
rect 1317 140335 1340 140369
rect 1133 139791 1167 139825
rect 1225 139791 1259 139825
rect 1317 139791 1340 139825
rect 1133 139247 1167 139281
rect 1225 139247 1259 139281
rect 1317 139247 1340 139281
rect 1133 138703 1167 138737
rect 1225 138703 1259 138737
rect 1317 138703 1340 138737
rect 1133 138159 1167 138193
rect 1225 138159 1259 138193
rect 1317 138159 1340 138193
rect 1133 137615 1167 137649
rect 1225 137615 1259 137649
rect 1317 137615 1340 137649
rect 1133 137071 1167 137105
rect 1225 137071 1259 137105
rect 1317 137071 1340 137105
rect 1133 136527 1167 136561
rect 1225 136527 1259 136561
rect 1317 136527 1340 136561
rect 1133 135983 1167 136017
rect 1225 135983 1259 136017
rect 1317 135983 1340 136017
rect 1133 135439 1167 135473
rect 1225 135439 1259 135473
rect 1317 135439 1340 135473
rect 1133 134895 1167 134929
rect 1225 134895 1259 134929
rect 1317 134895 1340 134929
rect 1133 134351 1167 134385
rect 1225 134351 1259 134385
rect 1317 134351 1340 134385
rect 1133 133807 1167 133841
rect 1225 133807 1259 133841
rect 1317 133807 1340 133841
rect 1133 133263 1167 133297
rect 1225 133263 1259 133297
rect 1317 133263 1340 133297
rect 1133 132719 1167 132753
rect 1225 132719 1259 132753
rect 1317 132719 1340 132753
rect 1133 132175 1167 132209
rect 1225 132175 1259 132209
rect 1317 132175 1340 132209
rect 1133 131631 1167 131665
rect 1225 131631 1259 131665
rect 1317 131631 1340 131665
rect 1133 131087 1167 131121
rect 1225 131087 1259 131121
rect 1317 131087 1340 131121
rect 1133 130543 1167 130577
rect 1225 130543 1259 130577
rect 1317 130543 1340 130577
rect 1133 129999 1167 130033
rect 1225 129999 1259 130033
rect 1317 129999 1340 130033
rect 1133 129455 1167 129489
rect 1225 129455 1259 129489
rect 1317 129455 1340 129489
rect 1133 128911 1167 128945
rect 1225 128911 1259 128945
rect 1317 128911 1340 128945
rect 1133 128367 1167 128401
rect 1225 128367 1259 128401
rect 1317 128367 1340 128401
rect 1133 127823 1167 127857
rect 1225 127823 1259 127857
rect 1317 127823 1340 127857
rect 1133 127279 1167 127313
rect 1225 127279 1259 127313
rect 1317 127279 1340 127313
rect 1133 126735 1167 126769
rect 1225 126735 1259 126769
rect 1317 126735 1340 126769
rect 1133 126191 1167 126225
rect 1225 126191 1259 126225
rect 1317 126191 1340 126225
rect 1133 125647 1167 125681
rect 1225 125647 1259 125681
rect 1317 125647 1340 125681
rect 1133 125103 1167 125137
rect 1225 125103 1259 125137
rect 1317 125103 1340 125137
rect 1133 124559 1167 124593
rect 1225 124559 1259 124593
rect 1317 124559 1340 124593
rect 1133 124015 1167 124049
rect 1225 124015 1259 124049
rect 1317 124015 1340 124049
rect 1133 123471 1167 123505
rect 1225 123471 1259 123505
rect 1317 123471 1340 123505
rect 1133 122927 1167 122961
rect 1225 122927 1259 122961
rect 1317 122927 1340 122961
rect 1133 122383 1167 122417
rect 1225 122383 1259 122417
rect 1317 122383 1340 122417
rect 1133 121839 1167 121873
rect 1225 121839 1259 121873
rect 1317 121839 1340 121873
rect 1133 121295 1167 121329
rect 1225 121295 1259 121329
rect 1317 121295 1340 121329
rect 1133 120751 1167 120785
rect 1225 120751 1259 120785
rect 1317 120751 1340 120785
rect 1133 120207 1167 120241
rect 1225 120207 1259 120241
rect 1317 120207 1340 120241
rect 1133 119663 1167 119697
rect 1225 119663 1259 119697
rect 1317 119663 1340 119697
rect 1133 119119 1167 119153
rect 1225 119119 1259 119153
rect 1317 119119 1340 119153
rect 1133 118575 1167 118609
rect 1225 118575 1259 118609
rect 1317 118575 1340 118609
rect 1133 118031 1167 118065
rect 1225 118031 1259 118065
rect 1317 118031 1340 118065
rect 1133 117487 1167 117521
rect 1225 117487 1259 117521
rect 1317 117487 1340 117521
rect 1133 116943 1167 116977
rect 1225 116943 1259 116977
rect 1317 116943 1340 116977
rect 1133 116399 1167 116433
rect 1225 116399 1259 116433
rect 1317 116399 1340 116433
rect 1133 115855 1167 115889
rect 1225 115855 1259 115889
rect 1317 115855 1340 115889
rect 1133 115311 1167 115345
rect 1225 115311 1259 115345
rect 1317 115311 1340 115345
rect 1133 114767 1167 114801
rect 1225 114767 1259 114801
rect 1317 114767 1340 114801
rect 1133 114223 1167 114257
rect 1225 114223 1259 114257
rect 1317 114223 1340 114257
rect 1133 113679 1167 113713
rect 1225 113679 1259 113713
rect 1317 113679 1340 113713
rect 1133 113135 1167 113169
rect 1225 113135 1259 113169
rect 1317 113135 1340 113169
rect 1133 112591 1167 112625
rect 1225 112591 1259 112625
rect 1317 112591 1340 112625
rect 1133 112047 1167 112081
rect 1225 112047 1259 112081
rect 1317 112047 1340 112081
rect 1133 111503 1167 111537
rect 1225 111503 1259 111537
rect 1317 111503 1340 111537
rect 1133 110959 1167 110993
rect 1225 110959 1259 110993
rect 1317 110959 1340 110993
rect 1133 110415 1167 110449
rect 1225 110415 1259 110449
rect 1317 110415 1340 110449
rect 1133 109871 1167 109905
rect 1225 109871 1259 109905
rect 1317 109871 1340 109905
rect 1133 109327 1167 109361
rect 1225 109327 1259 109361
rect 1317 109327 1340 109361
rect 1133 108783 1167 108817
rect 1225 108783 1259 108817
rect 1317 108783 1340 108817
rect 1133 108239 1167 108273
rect 1225 108239 1259 108273
rect 1317 108239 1340 108273
rect 1133 107695 1167 107729
rect 1225 107695 1259 107729
rect 1317 107695 1340 107729
rect 1133 107151 1167 107185
rect 1225 107151 1259 107185
rect 1317 107151 1340 107185
rect 1133 106607 1167 106641
rect 1225 106607 1259 106641
rect 1317 106607 1340 106641
rect 1133 106063 1167 106097
rect 1225 106063 1259 106097
rect 1317 106063 1340 106097
rect 1133 105519 1167 105553
rect 1225 105519 1259 105553
rect 1317 105519 1340 105553
rect 1133 104975 1167 105009
rect 1225 104975 1259 105009
rect 1317 104975 1340 105009
rect 1133 104431 1167 104465
rect 1225 104431 1259 104465
rect 1317 104431 1340 104465
rect 1133 103887 1167 103921
rect 1225 103887 1259 103921
rect 1317 103887 1340 103921
rect 1133 103343 1167 103377
rect 1225 103343 1259 103377
rect 1317 103343 1340 103377
rect 1133 102799 1167 102833
rect 1225 102799 1259 102833
rect 1317 102799 1340 102833
rect 1133 102255 1167 102289
rect 1225 102255 1259 102289
rect 1317 102255 1340 102289
rect 1133 101711 1167 101745
rect 1225 101711 1259 101745
rect 1317 101711 1340 101745
rect 1133 101167 1167 101201
rect 1225 101167 1259 101201
rect 1317 101167 1340 101201
rect 1133 100623 1167 100657
rect 1225 100623 1259 100657
rect 1317 100623 1340 100657
rect 1133 100079 1167 100113
rect 1225 100079 1259 100113
rect 1317 100079 1340 100113
rect 1133 99535 1167 99569
rect 1225 99535 1259 99569
rect 1317 99535 1340 99569
rect 1133 98991 1167 99025
rect 1225 98991 1259 99025
rect 1317 98991 1340 99025
rect 1133 98447 1167 98481
rect 1225 98447 1259 98481
rect 1317 98447 1340 98481
rect 1133 97903 1167 97937
rect 1225 97903 1259 97937
rect 1317 97903 1340 97937
rect 1133 97359 1167 97393
rect 1225 97359 1259 97393
rect 1317 97359 1340 97393
rect 1133 96815 1167 96849
rect 1225 96815 1259 96849
rect 1317 96815 1340 96849
rect 1133 96271 1167 96305
rect 1225 96271 1259 96305
rect 1317 96271 1340 96305
rect 1133 95727 1167 95761
rect 1225 95727 1259 95761
rect 1317 95727 1340 95761
rect 1133 95183 1167 95217
rect 1225 95183 1259 95217
rect 1317 95183 1340 95217
rect 1133 94639 1167 94673
rect 1225 94639 1259 94673
rect 1317 94639 1340 94673
rect 1133 94095 1167 94129
rect 1225 94095 1259 94129
rect 1317 94095 1340 94129
rect 1133 93551 1167 93585
rect 1225 93551 1259 93585
rect 1317 93551 1340 93585
rect 1133 93007 1167 93041
rect 1225 93007 1259 93041
rect 1317 93007 1340 93041
rect 1133 92463 1167 92497
rect 1225 92463 1259 92497
rect 1317 92463 1340 92497
rect 1133 91919 1167 91953
rect 1225 91919 1259 91953
rect 1317 91919 1340 91953
rect 1133 91375 1167 91409
rect 1225 91375 1259 91409
rect 1317 91375 1340 91409
rect 1133 90831 1167 90865
rect 1225 90831 1259 90865
rect 1317 90831 1340 90865
rect 1133 90287 1167 90321
rect 1225 90287 1259 90321
rect 1317 90287 1340 90321
rect 1133 89743 1167 89777
rect 1225 89743 1259 89777
rect 1317 89743 1340 89777
rect 1133 89199 1167 89233
rect 1225 89199 1259 89233
rect 1317 89199 1340 89233
rect 1133 88655 1167 88689
rect 1225 88655 1259 88689
rect 1317 88655 1340 88689
rect 1133 88111 1167 88145
rect 1225 88111 1259 88145
rect 1317 88111 1340 88145
rect 1133 87567 1167 87601
rect 1225 87567 1259 87601
rect 1317 87567 1340 87601
rect 1133 87023 1167 87057
rect 1225 87023 1259 87057
rect 1317 87023 1340 87057
rect 1133 86479 1167 86513
rect 1225 86479 1259 86513
rect 1317 86479 1340 86513
rect 1133 85935 1167 85969
rect 1225 85935 1259 85969
rect 1317 85935 1340 85969
rect 1133 85391 1167 85425
rect 1225 85391 1259 85425
rect 1317 85391 1340 85425
rect 1133 84847 1167 84881
rect 1225 84847 1259 84881
rect 1317 84847 1340 84881
rect 1133 84303 1167 84337
rect 1225 84303 1259 84337
rect 1317 84303 1340 84337
rect 1133 83759 1167 83793
rect 1225 83759 1259 83793
rect 1317 83759 1340 83793
rect 1133 83215 1167 83249
rect 1225 83215 1259 83249
rect 1317 83215 1340 83249
rect 1133 82671 1167 82705
rect 1225 82671 1259 82705
rect 1317 82671 1340 82705
rect 1133 82127 1167 82161
rect 1225 82127 1259 82161
rect 1317 82127 1340 82161
rect 1133 81583 1167 81617
rect 1225 81583 1259 81617
rect 1317 81583 1340 81617
rect 1133 81039 1167 81073
rect 1225 81039 1259 81073
rect 1317 81039 1340 81073
rect 1133 80495 1167 80529
rect 1225 80495 1259 80529
rect 1317 80495 1340 80529
rect 1133 79951 1167 79985
rect 1225 79951 1259 79985
rect 1317 79951 1340 79985
rect 1133 79407 1167 79441
rect 1225 79407 1259 79441
rect 1317 79407 1340 79441
rect 1133 78863 1167 78897
rect 1225 78863 1259 78897
rect 1317 78863 1340 78897
rect 1133 78319 1167 78353
rect 1225 78319 1259 78353
rect 1317 78319 1340 78353
rect 1133 77775 1167 77809
rect 1225 77775 1259 77809
rect 1317 77775 1340 77809
rect 1133 77231 1167 77265
rect 1225 77231 1259 77265
rect 1317 77231 1340 77265
rect 1133 76687 1167 76721
rect 1225 76687 1259 76721
rect 1317 76687 1340 76721
rect 1133 76143 1167 76177
rect 1225 76143 1259 76177
rect 1317 76143 1340 76177
rect 1133 75599 1167 75633
rect 1225 75599 1259 75633
rect 1317 75599 1340 75633
rect 1133 75055 1167 75089
rect 1225 75055 1259 75089
rect 1317 75055 1340 75089
rect 1133 74511 1167 74545
rect 1225 74511 1259 74545
rect 1317 74511 1340 74545
rect 1133 73967 1167 74001
rect 1225 73967 1259 74001
rect 1317 73967 1340 74001
rect 1133 73423 1167 73457
rect 1225 73423 1259 73457
rect 1317 73423 1340 73457
rect 1133 72879 1167 72913
rect 1225 72879 1259 72913
rect 1317 72879 1340 72913
rect 1133 72335 1167 72369
rect 1225 72335 1259 72369
rect 1317 72335 1340 72369
rect 1133 71791 1167 71825
rect 1225 71791 1259 71825
rect 1317 71791 1340 71825
rect 1133 71247 1167 71281
rect 1225 71247 1259 71281
rect 1317 71247 1340 71281
rect 1133 70703 1167 70737
rect 1225 70703 1259 70737
rect 1317 70703 1340 70737
rect 1133 70159 1167 70193
rect 1225 70159 1259 70193
rect 1317 70159 1340 70193
rect 1133 69615 1167 69649
rect 1225 69615 1259 69649
rect 1317 69615 1340 69649
rect 1133 69071 1167 69105
rect 1225 69071 1259 69105
rect 1317 69071 1340 69105
rect 1133 68527 1167 68561
rect 1225 68527 1259 68561
rect 1317 68527 1340 68561
rect 1133 67983 1167 68017
rect 1225 67983 1259 68017
rect 1317 67983 1340 68017
rect 1133 67439 1167 67473
rect 1225 67439 1259 67473
rect 1317 67439 1340 67473
rect 1133 66895 1167 66929
rect 1225 66895 1259 66929
rect 1317 66895 1340 66929
rect 1133 66351 1167 66385
rect 1225 66351 1259 66385
rect 1317 66351 1340 66385
rect 1133 65807 1167 65841
rect 1225 65807 1259 65841
rect 1317 65807 1340 65841
rect 1133 65263 1167 65297
rect 1225 65263 1259 65297
rect 1317 65263 1340 65297
rect 1133 64719 1167 64753
rect 1225 64719 1259 64753
rect 1317 64719 1340 64753
rect 1133 64175 1167 64209
rect 1225 64175 1259 64209
rect 1317 64175 1340 64209
rect 1133 63631 1167 63665
rect 1225 63631 1259 63665
rect 1317 63631 1340 63665
rect 1133 63087 1167 63121
rect 1225 63087 1259 63121
rect 1317 63087 1340 63121
rect 1133 62543 1167 62577
rect 1225 62543 1259 62577
rect 1317 62543 1340 62577
rect 1133 61999 1167 62033
rect 1225 61999 1259 62033
rect 1317 61999 1340 62033
rect 1133 61455 1167 61489
rect 1225 61455 1259 61489
rect 1317 61455 1340 61489
rect 1133 60911 1167 60945
rect 1225 60911 1259 60945
rect 1317 60911 1340 60945
rect 1133 60367 1167 60401
rect 1225 60367 1259 60401
rect 1317 60367 1340 60401
rect 1133 59823 1167 59857
rect 1225 59823 1259 59857
rect 1317 59823 1340 59857
rect 1133 59279 1167 59313
rect 1225 59279 1259 59313
rect 1317 59279 1340 59313
rect 1133 58735 1167 58769
rect 1225 58735 1259 58769
rect 1317 58735 1340 58769
rect 1133 58191 1167 58225
rect 1225 58191 1259 58225
rect 1317 58191 1340 58225
rect 1133 57647 1167 57681
rect 1225 57647 1259 57681
rect 1317 57647 1340 57681
rect 1133 57103 1167 57137
rect 1225 57103 1259 57137
rect 1317 57103 1340 57137
rect 1133 56559 1167 56593
rect 1225 56559 1259 56593
rect 1317 56559 1340 56593
rect 1133 56015 1167 56049
rect 1225 56015 1259 56049
rect 1317 56015 1340 56049
rect 1133 55471 1167 55505
rect 1225 55471 1259 55505
rect 1317 55471 1340 55505
rect 1133 54927 1167 54961
rect 1225 54927 1259 54961
rect 1317 54927 1340 54961
rect 1133 54383 1167 54417
rect 1225 54383 1259 54417
rect 1317 54383 1340 54417
rect 1133 53839 1167 53873
rect 1225 53839 1259 53873
rect 1317 53839 1340 53873
rect 1133 53295 1167 53329
rect 1225 53295 1259 53329
rect 1317 53295 1340 53329
rect 1133 52751 1167 52785
rect 1225 52751 1259 52785
rect 1317 52751 1340 52785
rect 1133 52207 1167 52241
rect 1225 52207 1259 52241
rect 1317 52207 1340 52241
rect 1133 51663 1167 51697
rect 1225 51663 1259 51697
rect 1317 51663 1340 51697
rect 1133 51119 1167 51153
rect 1225 51119 1259 51153
rect 1317 51119 1340 51153
rect 1133 50575 1167 50609
rect 1225 50575 1259 50609
rect 1317 50575 1340 50609
rect 1133 50031 1167 50065
rect 1225 50031 1259 50065
rect 1317 50031 1340 50065
rect 1133 49487 1167 49521
rect 1225 49487 1259 49521
rect 1317 49487 1340 49521
rect 1133 48943 1167 48977
rect 1225 48943 1259 48977
rect 1317 48943 1340 48977
rect 1133 48399 1167 48433
rect 1225 48399 1259 48433
rect 1317 48399 1340 48433
rect 1133 47855 1167 47889
rect 1225 47855 1259 47889
rect 1317 47855 1340 47889
rect 1133 47311 1167 47345
rect 1225 47311 1259 47345
rect 1317 47311 1340 47345
rect 1133 46767 1167 46801
rect 1225 46767 1259 46801
rect 1317 46767 1340 46801
rect 1133 46223 1167 46257
rect 1225 46223 1259 46257
rect 1317 46223 1340 46257
rect 1133 45679 1167 45713
rect 1225 45679 1259 45713
rect 1317 45679 1340 45713
rect 1133 45135 1167 45169
rect 1225 45135 1259 45169
rect 1317 45135 1340 45169
rect 1133 44591 1167 44625
rect 1225 44591 1259 44625
rect 1317 44591 1340 44625
rect 1133 44047 1167 44081
rect 1225 44047 1259 44081
rect 1317 44047 1340 44081
rect 1133 43503 1167 43537
rect 1225 43503 1259 43537
rect 1317 43503 1340 43537
rect 1133 42959 1167 42993
rect 1225 42959 1259 42993
rect 1317 42959 1340 42993
rect 1133 42415 1167 42449
rect 1225 42415 1259 42449
rect 1317 42415 1340 42449
rect 1133 41871 1167 41905
rect 1225 41871 1259 41905
rect 1317 41871 1340 41905
rect 1133 41327 1167 41361
rect 1225 41327 1259 41361
rect 1317 41327 1340 41361
rect 1133 40783 1167 40817
rect 1225 40783 1259 40817
rect 1317 40783 1340 40817
rect 1133 40239 1167 40273
rect 1225 40239 1259 40273
rect 1317 40239 1340 40273
rect 1133 39695 1167 39729
rect 1225 39695 1259 39729
rect 1317 39695 1340 39729
rect 1133 39151 1167 39185
rect 1225 39151 1259 39185
rect 1317 39151 1340 39185
rect 1133 38607 1167 38641
rect 1225 38607 1259 38641
rect 1317 38607 1340 38641
rect 1133 38063 1167 38097
rect 1225 38063 1259 38097
rect 1317 38063 1340 38097
rect 1133 37519 1167 37553
rect 1225 37519 1259 37553
rect 1317 37519 1340 37553
rect 1133 36975 1167 37009
rect 1225 36975 1259 37009
rect 1317 36975 1340 37009
rect 1133 36431 1167 36465
rect 1225 36431 1259 36465
rect 1317 36431 1340 36465
rect 1133 35887 1167 35921
rect 1225 35887 1259 35921
rect 1317 35887 1340 35921
rect 1133 35343 1167 35377
rect 1225 35343 1259 35377
rect 1317 35343 1340 35377
rect 1133 34799 1167 34833
rect 1225 34799 1259 34833
rect 1317 34799 1340 34833
rect 1133 34255 1167 34289
rect 1225 34255 1259 34289
rect 1317 34255 1340 34289
rect 1133 33711 1167 33745
rect 1225 33711 1259 33745
rect 1317 33711 1340 33745
rect 1133 33167 1167 33201
rect 1225 33167 1259 33201
rect 1317 33167 1340 33201
rect 1133 32623 1167 32657
rect 1225 32623 1259 32657
rect 1317 32623 1340 32657
rect 1133 32079 1167 32113
rect 1225 32079 1259 32113
rect 1317 32079 1340 32113
rect 1133 31535 1167 31569
rect 1225 31535 1259 31569
rect 1317 31535 1340 31569
rect 1133 30991 1167 31025
rect 1225 30991 1259 31025
rect 1317 30991 1340 31025
rect 1133 30447 1167 30481
rect 1225 30447 1259 30481
rect 1317 30447 1340 30481
rect 1133 29903 1167 29937
rect 1225 29903 1259 29937
rect 1317 29903 1340 29937
rect 1133 29359 1167 29393
rect 1225 29359 1259 29393
rect 1317 29359 1340 29393
rect 1133 28815 1167 28849
rect 1225 28815 1259 28849
rect 1317 28815 1340 28849
rect 1133 28271 1167 28305
rect 1225 28271 1259 28305
rect 1317 28271 1340 28305
rect 1133 27727 1167 27761
rect 1225 27727 1259 27761
rect 1317 27727 1340 27761
rect 1133 27183 1167 27217
rect 1225 27183 1259 27217
rect 1317 27183 1340 27217
rect 1133 26639 1167 26673
rect 1225 26639 1259 26673
rect 1317 26639 1340 26673
rect 1133 26095 1167 26129
rect 1225 26095 1259 26129
rect 1317 26095 1340 26129
rect 1133 25551 1167 25585
rect 1225 25551 1259 25585
rect 1317 25551 1340 25585
rect 1133 25007 1167 25041
rect 1225 25007 1259 25041
rect 1317 25007 1340 25041
rect 1133 24463 1167 24497
rect 1225 24463 1259 24497
rect 1317 24463 1340 24497
rect 1133 23919 1167 23953
rect 1225 23919 1259 23953
rect 1317 23919 1340 23953
rect 1133 23375 1167 23409
rect 1225 23375 1259 23409
rect 1317 23375 1340 23409
rect 1133 22831 1167 22865
rect 1225 22831 1259 22865
rect 1317 22831 1340 22865
rect 1133 22287 1167 22321
rect 1225 22287 1259 22321
rect 1317 22287 1340 22321
rect 1133 21743 1167 21777
rect 1225 21743 1259 21777
rect 1317 21743 1340 21777
rect 1133 21199 1167 21233
rect 1225 21199 1259 21233
rect 1317 21199 1340 21233
rect 1133 20655 1167 20689
rect 1225 20655 1259 20689
rect 1317 20655 1340 20689
rect 1133 20111 1167 20145
rect 1225 20111 1259 20145
rect 1317 20111 1340 20145
rect 1133 19567 1167 19601
rect 1225 19567 1259 19601
rect 1317 19567 1340 19601
rect 1133 19023 1167 19057
rect 1225 19023 1259 19057
rect 1317 19023 1340 19057
rect 1133 18479 1167 18513
rect 1225 18479 1259 18513
rect 1317 18479 1340 18513
rect 1133 17935 1167 17969
rect 1225 17935 1259 17969
rect 1317 17935 1340 17969
rect 1133 17391 1167 17425
rect 1225 17391 1259 17425
rect 1317 17391 1340 17425
rect 1133 16847 1167 16881
rect 1225 16847 1259 16881
rect 1317 16847 1340 16881
rect 1133 16303 1167 16337
rect 1225 16303 1259 16337
rect 1317 16303 1340 16337
rect 1133 15759 1167 15793
rect 1225 15759 1259 15793
rect 1317 15759 1340 15793
rect 1133 15215 1167 15249
rect 1225 15215 1259 15249
rect 1317 15215 1340 15249
rect 1133 14671 1167 14705
rect 1225 14671 1259 14705
rect 1317 14671 1340 14705
rect 1133 14127 1167 14161
rect 1225 14127 1259 14161
rect 1317 14127 1340 14161
rect 1133 13583 1167 13617
rect 1225 13583 1259 13617
rect 1317 13583 1340 13617
rect 1133 13039 1167 13073
rect 1225 13039 1259 13073
rect 1317 13039 1340 13073
rect 1133 12495 1167 12529
rect 1225 12495 1259 12529
rect 1317 12495 1340 12529
rect 1133 11951 1167 11985
rect 1225 11951 1259 11985
rect 1317 11951 1340 11985
rect 1133 11407 1167 11441
rect 1225 11407 1259 11441
rect 1317 11407 1340 11441
rect 1133 10863 1167 10897
rect 1225 10863 1259 10897
rect 1317 10863 1340 10897
rect 1133 10319 1167 10353
rect 1225 10319 1259 10353
rect 1317 10319 1340 10353
rect 1133 9775 1167 9809
rect 1225 9775 1259 9809
rect 1317 9775 1340 9809
rect 1133 9231 1167 9265
rect 1225 9231 1259 9265
rect 1317 9231 1340 9265
rect 1133 8687 1167 8721
rect 1225 8687 1259 8721
rect 1317 8687 1340 8721
rect 1133 8143 1167 8177
rect 1225 8143 1259 8177
rect 1317 8143 1340 8177
rect 1133 7599 1167 7633
rect 1225 7599 1259 7633
rect 1317 7599 1340 7633
rect 1133 7055 1167 7089
rect 1225 7055 1259 7089
rect 1317 7055 1340 7089
rect 1133 6511 1167 6545
rect 1225 6511 1259 6545
rect 1317 6511 1340 6545
rect 1133 5967 1167 6001
rect 1225 5967 1259 6001
rect 1317 5967 1340 6001
rect 1133 5423 1167 5457
rect 1225 5423 1259 5457
rect 1317 5423 1340 5457
rect 1133 4879 1167 4913
rect 1225 4879 1259 4913
rect 1317 4879 1340 4913
rect 1133 4335 1167 4369
rect 1225 4335 1259 4369
rect 1317 4335 1340 4369
rect 1133 3791 1167 3825
rect 1225 3791 1259 3825
rect 1317 3791 1340 3825
rect 1133 3247 1167 3281
rect 1225 3247 1259 3281
rect 1317 3247 1340 3281
rect 1133 2703 1167 2737
rect 1225 2703 1259 2737
rect 1317 2703 1340 2737
rect 1133 2159 1167 2193
rect 1225 2159 1259 2193
rect 1317 2159 1340 2193
rect 298661 297551 298695 297585
rect 298753 297551 298787 297585
rect 298661 297007 298695 297041
rect 298753 297007 298787 297041
rect 298661 296463 298695 296497
rect 298753 296463 298787 296497
rect 298661 295919 298695 295953
rect 298753 295919 298787 295953
rect 298661 295375 298695 295409
rect 298753 295375 298787 295409
rect 298661 294831 298695 294865
rect 298753 294831 298787 294865
rect 298661 294287 298695 294321
rect 298753 294287 298787 294321
rect 298661 293743 298695 293777
rect 298753 293743 298787 293777
rect 298661 293199 298695 293233
rect 298753 293199 298787 293233
rect 298661 292655 298695 292689
rect 298753 292655 298787 292689
rect 298661 292111 298695 292145
rect 298753 292111 298787 292145
rect 298661 291567 298695 291601
rect 298753 291567 298787 291601
rect 298661 291023 298695 291057
rect 298753 291023 298787 291057
rect 298661 290479 298695 290513
rect 298753 290479 298787 290513
rect 298661 289935 298695 289969
rect 298753 289935 298787 289969
rect 298661 289391 298695 289425
rect 298753 289391 298787 289425
rect 298661 288847 298695 288881
rect 298753 288847 298787 288881
rect 298661 288303 298695 288337
rect 298753 288303 298787 288337
rect 298661 287759 298695 287793
rect 298753 287759 298787 287793
rect 298661 287215 298695 287249
rect 298753 287215 298787 287249
rect 298661 286671 298695 286705
rect 298753 286671 298787 286705
rect 298661 286127 298695 286161
rect 298753 286127 298787 286161
rect 298661 285583 298695 285617
rect 298753 285583 298787 285617
rect 298661 285039 298695 285073
rect 298753 285039 298787 285073
rect 298661 284495 298695 284529
rect 298753 284495 298787 284529
rect 298661 283951 298695 283985
rect 298753 283951 298787 283985
rect 298661 283407 298695 283441
rect 298753 283407 298787 283441
rect 298661 282863 298695 282897
rect 298753 282863 298787 282897
rect 298661 282319 298695 282353
rect 298753 282319 298787 282353
rect 298661 281775 298695 281809
rect 298753 281775 298787 281809
rect 298661 281231 298695 281265
rect 298753 281231 298787 281265
rect 298661 280687 298695 280721
rect 298753 280687 298787 280721
rect 298661 280143 298695 280177
rect 298753 280143 298787 280177
rect 298661 279599 298695 279633
rect 298753 279599 298787 279633
rect 298661 279055 298695 279089
rect 298753 279055 298787 279089
rect 298661 278511 298695 278545
rect 298753 278511 298787 278545
rect 298661 277967 298695 278001
rect 298753 277967 298787 278001
rect 298661 277423 298695 277457
rect 298753 277423 298787 277457
rect 298661 276879 298695 276913
rect 298753 276879 298787 276913
rect 298661 276335 298695 276369
rect 298753 276335 298787 276369
rect 298661 275791 298695 275825
rect 298753 275791 298787 275825
rect 298661 275247 298695 275281
rect 298753 275247 298787 275281
rect 298661 274703 298695 274737
rect 298753 274703 298787 274737
rect 298661 274159 298695 274193
rect 298753 274159 298787 274193
rect 298661 273615 298695 273649
rect 298753 273615 298787 273649
rect 298661 273071 298695 273105
rect 298753 273071 298787 273105
rect 298661 272527 298695 272561
rect 298753 272527 298787 272561
rect 298661 271983 298695 272017
rect 298753 271983 298787 272017
rect 298661 271439 298695 271473
rect 298753 271439 298787 271473
rect 298661 270895 298695 270929
rect 298753 270895 298787 270929
rect 298661 270351 298695 270385
rect 298753 270351 298787 270385
rect 298661 269807 298695 269841
rect 298753 269807 298787 269841
rect 298661 269263 298695 269297
rect 298753 269263 298787 269297
rect 298661 268719 298695 268753
rect 298753 268719 298787 268753
rect 298661 268175 298695 268209
rect 298753 268175 298787 268209
rect 298661 267631 298695 267665
rect 298753 267631 298787 267665
rect 298661 267087 298695 267121
rect 298753 267087 298787 267121
rect 298661 266543 298695 266577
rect 298753 266543 298787 266577
rect 298661 265999 298695 266033
rect 298753 265999 298787 266033
rect 298661 265455 298695 265489
rect 298753 265455 298787 265489
rect 298661 264911 298695 264945
rect 298753 264911 298787 264945
rect 298661 264367 298695 264401
rect 298753 264367 298787 264401
rect 298661 263823 298695 263857
rect 298753 263823 298787 263857
rect 298661 263279 298695 263313
rect 298753 263279 298787 263313
rect 298661 262735 298695 262769
rect 298753 262735 298787 262769
rect 298661 262191 298695 262225
rect 298753 262191 298787 262225
rect 298661 261647 298695 261681
rect 298753 261647 298787 261681
rect 298661 261103 298695 261137
rect 298753 261103 298787 261137
rect 298661 260559 298695 260593
rect 298753 260559 298787 260593
rect 298661 260015 298695 260049
rect 298753 260015 298787 260049
rect 298661 259471 298695 259505
rect 298753 259471 298787 259505
rect 298661 258927 298695 258961
rect 298753 258927 298787 258961
rect 298661 258383 298695 258417
rect 298753 258383 298787 258417
rect 298661 257839 298695 257873
rect 298753 257839 298787 257873
rect 298661 257295 298695 257329
rect 298753 257295 298787 257329
rect 298661 256751 298695 256785
rect 298753 256751 298787 256785
rect 298661 256207 298695 256241
rect 298753 256207 298787 256241
rect 298661 255663 298695 255697
rect 298753 255663 298787 255697
rect 298661 255119 298695 255153
rect 298753 255119 298787 255153
rect 298661 254575 298695 254609
rect 298753 254575 298787 254609
rect 298661 254031 298695 254065
rect 298753 254031 298787 254065
rect 298661 253487 298695 253521
rect 298753 253487 298787 253521
rect 298661 252943 298695 252977
rect 298753 252943 298787 252977
rect 298661 252399 298695 252433
rect 298753 252399 298787 252433
rect 298661 251855 298695 251889
rect 298753 251855 298787 251889
rect 298661 251311 298695 251345
rect 298753 251311 298787 251345
rect 298661 250767 298695 250801
rect 298753 250767 298787 250801
rect 298661 250223 298695 250257
rect 298753 250223 298787 250257
rect 298661 249679 298695 249713
rect 298753 249679 298787 249713
rect 298661 249135 298695 249169
rect 298753 249135 298787 249169
rect 298661 248591 298695 248625
rect 298753 248591 298787 248625
rect 298661 248047 298695 248081
rect 298753 248047 298787 248081
rect 298661 247503 298695 247537
rect 298753 247503 298787 247537
rect 298661 246959 298695 246993
rect 298753 246959 298787 246993
rect 298661 246415 298695 246449
rect 298753 246415 298787 246449
rect 298661 245871 298695 245905
rect 298753 245871 298787 245905
rect 298661 245327 298695 245361
rect 298753 245327 298787 245361
rect 298661 244783 298695 244817
rect 298753 244783 298787 244817
rect 298661 244239 298695 244273
rect 298753 244239 298787 244273
rect 298661 243695 298695 243729
rect 298753 243695 298787 243729
rect 298661 243151 298695 243185
rect 298753 243151 298787 243185
rect 298661 242607 298695 242641
rect 298753 242607 298787 242641
rect 298661 242063 298695 242097
rect 298753 242063 298787 242097
rect 298661 241519 298695 241553
rect 298753 241519 298787 241553
rect 298661 240975 298695 241009
rect 298753 240975 298787 241009
rect 298661 240431 298695 240465
rect 298753 240431 298787 240465
rect 298661 239887 298695 239921
rect 298753 239887 298787 239921
rect 298661 239343 298695 239377
rect 298753 239343 298787 239377
rect 298661 238799 298695 238833
rect 298753 238799 298787 238833
rect 298661 238255 298695 238289
rect 298753 238255 298787 238289
rect 298661 237711 298695 237745
rect 298753 237711 298787 237745
rect 298661 237167 298695 237201
rect 298753 237167 298787 237201
rect 298661 236623 298695 236657
rect 298753 236623 298787 236657
rect 298661 236079 298695 236113
rect 298753 236079 298787 236113
rect 298661 235535 298695 235569
rect 298753 235535 298787 235569
rect 298661 234991 298695 235025
rect 298753 234991 298787 235025
rect 298661 234447 298695 234481
rect 298753 234447 298787 234481
rect 298661 233903 298695 233937
rect 298753 233903 298787 233937
rect 298661 233359 298695 233393
rect 298753 233359 298787 233393
rect 298661 232815 298695 232849
rect 298753 232815 298787 232849
rect 298661 232271 298695 232305
rect 298753 232271 298787 232305
rect 298661 231727 298695 231761
rect 298753 231727 298787 231761
rect 298661 231183 298695 231217
rect 298753 231183 298787 231217
rect 298661 230639 298695 230673
rect 298753 230639 298787 230673
rect 298661 230095 298695 230129
rect 298753 230095 298787 230129
rect 298661 229551 298695 229585
rect 298753 229551 298787 229585
rect 298661 229007 298695 229041
rect 298753 229007 298787 229041
rect 298661 228463 298695 228497
rect 298753 228463 298787 228497
rect 298661 227919 298695 227953
rect 298753 227919 298787 227953
rect 298661 227375 298695 227409
rect 298753 227375 298787 227409
rect 298661 226831 298695 226865
rect 298753 226831 298787 226865
rect 298661 226287 298695 226321
rect 298753 226287 298787 226321
rect 298661 225743 298695 225777
rect 298753 225743 298787 225777
rect 298661 225199 298695 225233
rect 298753 225199 298787 225233
rect 298661 224655 298695 224689
rect 298753 224655 298787 224689
rect 298661 224111 298695 224145
rect 298753 224111 298787 224145
rect 298661 223567 298695 223601
rect 298753 223567 298787 223601
rect 298661 223023 298695 223057
rect 298753 223023 298787 223057
rect 298661 222479 298695 222513
rect 298753 222479 298787 222513
rect 298661 221935 298695 221969
rect 298753 221935 298787 221969
rect 298661 221391 298695 221425
rect 298753 221391 298787 221425
rect 298661 220847 298695 220881
rect 298753 220847 298787 220881
rect 298661 220303 298695 220337
rect 298753 220303 298787 220337
rect 298661 219759 298695 219793
rect 298753 219759 298787 219793
rect 298661 219215 298695 219249
rect 298753 219215 298787 219249
rect 298661 218671 298695 218705
rect 298753 218671 298787 218705
rect 298661 218127 298695 218161
rect 298753 218127 298787 218161
rect 298661 217583 298695 217617
rect 298753 217583 298787 217617
rect 298661 217039 298695 217073
rect 298753 217039 298787 217073
rect 298661 216495 298695 216529
rect 298753 216495 298787 216529
rect 298661 215951 298695 215985
rect 298753 215951 298787 215985
rect 298661 215407 298695 215441
rect 298753 215407 298787 215441
rect 298661 214863 298695 214897
rect 298753 214863 298787 214897
rect 298661 214319 298695 214353
rect 298753 214319 298787 214353
rect 298661 213775 298695 213809
rect 298753 213775 298787 213809
rect 298661 213231 298695 213265
rect 298753 213231 298787 213265
rect 298661 212687 298695 212721
rect 298753 212687 298787 212721
rect 298661 212143 298695 212177
rect 298753 212143 298787 212177
rect 298661 211599 298695 211633
rect 298753 211599 298787 211633
rect 298661 211055 298695 211089
rect 298753 211055 298787 211089
rect 298661 210511 298695 210545
rect 298753 210511 298787 210545
rect 298661 209967 298695 210001
rect 298753 209967 298787 210001
rect 298661 209423 298695 209457
rect 298753 209423 298787 209457
rect 298661 208879 298695 208913
rect 298753 208879 298787 208913
rect 298661 208335 298695 208369
rect 298753 208335 298787 208369
rect 298661 207791 298695 207825
rect 298753 207791 298787 207825
rect 298661 207247 298695 207281
rect 298753 207247 298787 207281
rect 298661 206703 298695 206737
rect 298753 206703 298787 206737
rect 298661 206159 298695 206193
rect 298753 206159 298787 206193
rect 298661 205615 298695 205649
rect 298753 205615 298787 205649
rect 298661 205071 298695 205105
rect 298753 205071 298787 205105
rect 298661 204527 298695 204561
rect 298753 204527 298787 204561
rect 298661 203983 298695 204017
rect 298753 203983 298787 204017
rect 298661 203439 298695 203473
rect 298753 203439 298787 203473
rect 298661 202895 298695 202929
rect 298753 202895 298787 202929
rect 298661 202351 298695 202385
rect 298753 202351 298787 202385
rect 298661 201807 298695 201841
rect 298753 201807 298787 201841
rect 298661 201263 298695 201297
rect 298753 201263 298787 201297
rect 298661 200719 298695 200753
rect 298753 200719 298787 200753
rect 298661 200175 298695 200209
rect 298753 200175 298787 200209
rect 298661 199631 298695 199665
rect 298753 199631 298787 199665
rect 298661 199087 298695 199121
rect 298753 199087 298787 199121
rect 298661 198543 298695 198577
rect 298753 198543 298787 198577
rect 298661 197999 298695 198033
rect 298753 197999 298787 198033
rect 298661 197455 298695 197489
rect 298753 197455 298787 197489
rect 298661 196911 298695 196945
rect 298753 196911 298787 196945
rect 298661 196367 298695 196401
rect 298753 196367 298787 196401
rect 298661 195823 298695 195857
rect 298753 195823 298787 195857
rect 298661 195279 298695 195313
rect 298753 195279 298787 195313
rect 298661 194735 298695 194769
rect 298753 194735 298787 194769
rect 298661 194191 298695 194225
rect 298753 194191 298787 194225
rect 298661 193647 298695 193681
rect 298753 193647 298787 193681
rect 298661 193103 298695 193137
rect 298753 193103 298787 193137
rect 298661 192559 298695 192593
rect 298753 192559 298787 192593
rect 298661 192015 298695 192049
rect 298753 192015 298787 192049
rect 298661 191471 298695 191505
rect 298753 191471 298787 191505
rect 298661 190927 298695 190961
rect 298753 190927 298787 190961
rect 298661 190383 298695 190417
rect 298753 190383 298787 190417
rect 298661 189839 298695 189873
rect 298753 189839 298787 189873
rect 298661 189295 298695 189329
rect 298753 189295 298787 189329
rect 298661 188751 298695 188785
rect 298753 188751 298787 188785
rect 298661 188207 298695 188241
rect 298753 188207 298787 188241
rect 298661 187663 298695 187697
rect 298753 187663 298787 187697
rect 298661 187119 298695 187153
rect 298753 187119 298787 187153
rect 298661 186575 298695 186609
rect 298753 186575 298787 186609
rect 298661 186031 298695 186065
rect 298753 186031 298787 186065
rect 298661 185487 298695 185521
rect 298753 185487 298787 185521
rect 298661 184943 298695 184977
rect 298753 184943 298787 184977
rect 298661 184399 298695 184433
rect 298753 184399 298787 184433
rect 298661 183855 298695 183889
rect 298753 183855 298787 183889
rect 298661 183311 298695 183345
rect 298753 183311 298787 183345
rect 298661 182767 298695 182801
rect 298753 182767 298787 182801
rect 298661 182223 298695 182257
rect 298753 182223 298787 182257
rect 298661 181679 298695 181713
rect 298753 181679 298787 181713
rect 298661 181135 298695 181169
rect 298753 181135 298787 181169
rect 298661 180591 298695 180625
rect 298753 180591 298787 180625
rect 298661 180047 298695 180081
rect 298753 180047 298787 180081
rect 298661 179503 298695 179537
rect 298753 179503 298787 179537
rect 298661 178959 298695 178993
rect 298753 178959 298787 178993
rect 298661 178415 298695 178449
rect 298753 178415 298787 178449
rect 298661 177871 298695 177905
rect 298753 177871 298787 177905
rect 298661 177327 298695 177361
rect 298753 177327 298787 177361
rect 298661 176783 298695 176817
rect 298753 176783 298787 176817
rect 298661 176239 298695 176273
rect 298753 176239 298787 176273
rect 298661 175695 298695 175729
rect 298753 175695 298787 175729
rect 298661 175151 298695 175185
rect 298753 175151 298787 175185
rect 298661 174607 298695 174641
rect 298753 174607 298787 174641
rect 298661 174063 298695 174097
rect 298753 174063 298787 174097
rect 298661 173519 298695 173553
rect 298753 173519 298787 173553
rect 298661 172975 298695 173009
rect 298753 172975 298787 173009
rect 298661 172431 298695 172465
rect 298753 172431 298787 172465
rect 298661 171887 298695 171921
rect 298753 171887 298787 171921
rect 298661 171343 298695 171377
rect 298753 171343 298787 171377
rect 298661 170799 298695 170833
rect 298753 170799 298787 170833
rect 298661 170255 298695 170289
rect 298753 170255 298787 170289
rect 298661 169711 298695 169745
rect 298753 169711 298787 169745
rect 298661 169167 298695 169201
rect 298753 169167 298787 169201
rect 298661 168623 298695 168657
rect 298753 168623 298787 168657
rect 298661 168079 298695 168113
rect 298753 168079 298787 168113
rect 298661 167535 298695 167569
rect 298753 167535 298787 167569
rect 298661 166991 298695 167025
rect 298753 166991 298787 167025
rect 298661 166447 298695 166481
rect 298753 166447 298787 166481
rect 298661 165903 298695 165937
rect 298753 165903 298787 165937
rect 298661 165359 298695 165393
rect 298753 165359 298787 165393
rect 298661 164815 298695 164849
rect 298753 164815 298787 164849
rect 298661 164271 298695 164305
rect 298753 164271 298787 164305
rect 298661 163727 298695 163761
rect 298753 163727 298787 163761
rect 298661 163183 298695 163217
rect 298753 163183 298787 163217
rect 298661 162639 298695 162673
rect 298753 162639 298787 162673
rect 298661 162095 298695 162129
rect 298753 162095 298787 162129
rect 298661 161551 298695 161585
rect 298753 161551 298787 161585
rect 298661 161007 298695 161041
rect 298753 161007 298787 161041
rect 298661 160463 298695 160497
rect 298753 160463 298787 160497
rect 298661 159919 298695 159953
rect 298753 159919 298787 159953
rect 298661 159375 298695 159409
rect 298753 159375 298787 159409
rect 298661 158831 298695 158865
rect 298753 158831 298787 158865
rect 298661 158287 298695 158321
rect 298753 158287 298787 158321
rect 298661 157743 298695 157777
rect 298753 157743 298787 157777
rect 298661 157199 298695 157233
rect 298753 157199 298787 157233
rect 298661 156655 298695 156689
rect 298753 156655 298787 156689
rect 298661 156111 298695 156145
rect 298753 156111 298787 156145
rect 298661 155567 298695 155601
rect 298753 155567 298787 155601
rect 298661 155023 298695 155057
rect 298753 155023 298787 155057
rect 298661 154479 298695 154513
rect 298753 154479 298787 154513
rect 298661 153935 298695 153969
rect 298753 153935 298787 153969
rect 298661 153391 298695 153425
rect 298753 153391 298787 153425
rect 298661 152847 298695 152881
rect 298753 152847 298787 152881
rect 298661 152303 298695 152337
rect 298753 152303 298787 152337
rect 298661 151759 298695 151793
rect 298753 151759 298787 151793
rect 298661 151215 298695 151249
rect 298753 151215 298787 151249
rect 298661 150671 298695 150705
rect 298753 150671 298787 150705
rect 298661 150127 298695 150161
rect 298753 150127 298787 150161
rect 298661 149583 298695 149617
rect 298753 149583 298787 149617
rect 298661 149039 298695 149073
rect 298753 149039 298787 149073
rect 298661 148495 298695 148529
rect 298753 148495 298787 148529
rect 298661 147951 298695 147985
rect 298753 147951 298787 147985
rect 298661 147407 298695 147441
rect 298753 147407 298787 147441
rect 298661 146863 298695 146897
rect 298753 146863 298787 146897
rect 298661 146319 298695 146353
rect 298753 146319 298787 146353
rect 298661 145775 298695 145809
rect 298753 145775 298787 145809
rect 298661 145231 298695 145265
rect 298753 145231 298787 145265
rect 298661 144687 298695 144721
rect 298753 144687 298787 144721
rect 298661 144143 298695 144177
rect 298753 144143 298787 144177
rect 298661 143599 298695 143633
rect 298753 143599 298787 143633
rect 298661 143055 298695 143089
rect 298753 143055 298787 143089
rect 298661 142511 298695 142545
rect 298753 142511 298787 142545
rect 298661 141967 298695 142001
rect 298753 141967 298787 142001
rect 298661 141423 298695 141457
rect 298753 141423 298787 141457
rect 298661 140879 298695 140913
rect 298753 140879 298787 140913
rect 298661 140335 298695 140369
rect 298753 140335 298787 140369
rect 298661 139791 298695 139825
rect 298753 139791 298787 139825
rect 298661 139247 298695 139281
rect 298753 139247 298787 139281
rect 298661 138703 298695 138737
rect 298753 138703 298787 138737
rect 298661 138159 298695 138193
rect 298753 138159 298787 138193
rect 298661 137615 298695 137649
rect 298753 137615 298787 137649
rect 298661 137071 298695 137105
rect 298753 137071 298787 137105
rect 298661 136527 298695 136561
rect 298753 136527 298787 136561
rect 298661 135983 298695 136017
rect 298753 135983 298787 136017
rect 298661 135439 298695 135473
rect 298753 135439 298787 135473
rect 298661 134895 298695 134929
rect 298753 134895 298787 134929
rect 298661 134351 298695 134385
rect 298753 134351 298787 134385
rect 298661 133807 298695 133841
rect 298753 133807 298787 133841
rect 298661 133263 298695 133297
rect 298753 133263 298787 133297
rect 298661 132719 298695 132753
rect 298753 132719 298787 132753
rect 298661 132175 298695 132209
rect 298753 132175 298787 132209
rect 298661 131631 298695 131665
rect 298753 131631 298787 131665
rect 298661 131087 298695 131121
rect 298753 131087 298787 131121
rect 298661 130543 298695 130577
rect 298753 130543 298787 130577
rect 298661 129999 298695 130033
rect 298753 129999 298787 130033
rect 298661 129455 298695 129489
rect 298753 129455 298787 129489
rect 298661 128911 298695 128945
rect 298753 128911 298787 128945
rect 298661 128367 298695 128401
rect 298753 128367 298787 128401
rect 298661 127823 298695 127857
rect 298753 127823 298787 127857
rect 298661 127279 298695 127313
rect 298753 127279 298787 127313
rect 298661 126735 298695 126769
rect 298753 126735 298787 126769
rect 298661 126191 298695 126225
rect 298753 126191 298787 126225
rect 298661 125647 298695 125681
rect 298753 125647 298787 125681
rect 298661 125103 298695 125137
rect 298753 125103 298787 125137
rect 298661 124559 298695 124593
rect 298753 124559 298787 124593
rect 298661 124015 298695 124049
rect 298753 124015 298787 124049
rect 298661 123471 298695 123505
rect 298753 123471 298787 123505
rect 298661 122927 298695 122961
rect 298753 122927 298787 122961
rect 298661 122383 298695 122417
rect 298753 122383 298787 122417
rect 298661 121839 298695 121873
rect 298753 121839 298787 121873
rect 298661 121295 298695 121329
rect 298753 121295 298787 121329
rect 298661 120751 298695 120785
rect 298753 120751 298787 120785
rect 298661 120207 298695 120241
rect 298753 120207 298787 120241
rect 298661 119663 298695 119697
rect 298753 119663 298787 119697
rect 298661 119119 298695 119153
rect 298753 119119 298787 119153
rect 298661 118575 298695 118609
rect 298753 118575 298787 118609
rect 298661 118031 298695 118065
rect 298753 118031 298787 118065
rect 298661 117487 298695 117521
rect 298753 117487 298787 117521
rect 298661 116943 298695 116977
rect 298753 116943 298787 116977
rect 298661 116399 298695 116433
rect 298753 116399 298787 116433
rect 298661 115855 298695 115889
rect 298753 115855 298787 115889
rect 298661 115311 298695 115345
rect 298753 115311 298787 115345
rect 298661 114767 298695 114801
rect 298753 114767 298787 114801
rect 298661 114223 298695 114257
rect 298753 114223 298787 114257
rect 298661 113679 298695 113713
rect 298753 113679 298787 113713
rect 298661 113135 298695 113169
rect 298753 113135 298787 113169
rect 298661 112591 298695 112625
rect 298753 112591 298787 112625
rect 298661 112047 298695 112081
rect 298753 112047 298787 112081
rect 298661 111503 298695 111537
rect 298753 111503 298787 111537
rect 298661 110959 298695 110993
rect 298753 110959 298787 110993
rect 298661 110415 298695 110449
rect 298753 110415 298787 110449
rect 298661 109871 298695 109905
rect 298753 109871 298787 109905
rect 298661 109327 298695 109361
rect 298753 109327 298787 109361
rect 298661 108783 298695 108817
rect 298753 108783 298787 108817
rect 298661 108239 298695 108273
rect 298753 108239 298787 108273
rect 298661 107695 298695 107729
rect 298753 107695 298787 107729
rect 298661 107151 298695 107185
rect 298753 107151 298787 107185
rect 298661 106607 298695 106641
rect 298753 106607 298787 106641
rect 298661 106063 298695 106097
rect 298753 106063 298787 106097
rect 298661 105519 298695 105553
rect 298753 105519 298787 105553
rect 298661 104975 298695 105009
rect 298753 104975 298787 105009
rect 298661 104431 298695 104465
rect 298753 104431 298787 104465
rect 298661 103887 298695 103921
rect 298753 103887 298787 103921
rect 298661 103343 298695 103377
rect 298753 103343 298787 103377
rect 298661 102799 298695 102833
rect 298753 102799 298787 102833
rect 298661 102255 298695 102289
rect 298753 102255 298787 102289
rect 298661 101711 298695 101745
rect 298753 101711 298787 101745
rect 298661 101167 298695 101201
rect 298753 101167 298787 101201
rect 298661 100623 298695 100657
rect 298753 100623 298787 100657
rect 298661 100079 298695 100113
rect 298753 100079 298787 100113
rect 298661 99535 298695 99569
rect 298753 99535 298787 99569
rect 298661 98991 298695 99025
rect 298753 98991 298787 99025
rect 298661 98447 298695 98481
rect 298753 98447 298787 98481
rect 298661 97903 298695 97937
rect 298753 97903 298787 97937
rect 298661 97359 298695 97393
rect 298753 97359 298787 97393
rect 298661 96815 298695 96849
rect 298753 96815 298787 96849
rect 298661 96271 298695 96305
rect 298753 96271 298787 96305
rect 298661 95727 298695 95761
rect 298753 95727 298787 95761
rect 298661 95183 298695 95217
rect 298753 95183 298787 95217
rect 298661 94639 298695 94673
rect 298753 94639 298787 94673
rect 298661 94095 298695 94129
rect 298753 94095 298787 94129
rect 298661 93551 298695 93585
rect 298753 93551 298787 93585
rect 298661 93007 298695 93041
rect 298753 93007 298787 93041
rect 298661 92463 298695 92497
rect 298753 92463 298787 92497
rect 298661 91919 298695 91953
rect 298753 91919 298787 91953
rect 298661 91375 298695 91409
rect 298753 91375 298787 91409
rect 298661 90831 298695 90865
rect 298753 90831 298787 90865
rect 298661 90287 298695 90321
rect 298753 90287 298787 90321
rect 298661 89743 298695 89777
rect 298753 89743 298787 89777
rect 298661 89199 298695 89233
rect 298753 89199 298787 89233
rect 298661 88655 298695 88689
rect 298753 88655 298787 88689
rect 298661 88111 298695 88145
rect 298753 88111 298787 88145
rect 298661 87567 298695 87601
rect 298753 87567 298787 87601
rect 298661 87023 298695 87057
rect 298753 87023 298787 87057
rect 298661 86479 298695 86513
rect 298753 86479 298787 86513
rect 298661 85935 298695 85969
rect 298753 85935 298787 85969
rect 298661 85391 298695 85425
rect 298753 85391 298787 85425
rect 298661 84847 298695 84881
rect 298753 84847 298787 84881
rect 298661 84303 298695 84337
rect 298753 84303 298787 84337
rect 298661 83759 298695 83793
rect 298753 83759 298787 83793
rect 298661 83215 298695 83249
rect 298753 83215 298787 83249
rect 298661 82671 298695 82705
rect 298753 82671 298787 82705
rect 298661 82127 298695 82161
rect 298753 82127 298787 82161
rect 298661 81583 298695 81617
rect 298753 81583 298787 81617
rect 298661 81039 298695 81073
rect 298753 81039 298787 81073
rect 298661 80495 298695 80529
rect 298753 80495 298787 80529
rect 298661 79951 298695 79985
rect 298753 79951 298787 79985
rect 298661 79407 298695 79441
rect 298753 79407 298787 79441
rect 298661 78863 298695 78897
rect 298753 78863 298787 78897
rect 298661 78319 298695 78353
rect 298753 78319 298787 78353
rect 298661 77775 298695 77809
rect 298753 77775 298787 77809
rect 298661 77231 298695 77265
rect 298753 77231 298787 77265
rect 298661 76687 298695 76721
rect 298753 76687 298787 76721
rect 298661 76143 298695 76177
rect 298753 76143 298787 76177
rect 298661 75599 298695 75633
rect 298753 75599 298787 75633
rect 298661 75055 298695 75089
rect 298753 75055 298787 75089
rect 298661 74511 298695 74545
rect 298753 74511 298787 74545
rect 298661 73967 298695 74001
rect 298753 73967 298787 74001
rect 298661 73423 298695 73457
rect 298753 73423 298787 73457
rect 298661 72879 298695 72913
rect 298753 72879 298787 72913
rect 298661 72335 298695 72369
rect 298753 72335 298787 72369
rect 298661 71791 298695 71825
rect 298753 71791 298787 71825
rect 298661 71247 298695 71281
rect 298753 71247 298787 71281
rect 298661 70703 298695 70737
rect 298753 70703 298787 70737
rect 298661 70159 298695 70193
rect 298753 70159 298787 70193
rect 298661 69615 298695 69649
rect 298753 69615 298787 69649
rect 298661 69071 298695 69105
rect 298753 69071 298787 69105
rect 298661 68527 298695 68561
rect 298753 68527 298787 68561
rect 298661 67983 298695 68017
rect 298753 67983 298787 68017
rect 298661 67439 298695 67473
rect 298753 67439 298787 67473
rect 298661 66895 298695 66929
rect 298753 66895 298787 66929
rect 298661 66351 298695 66385
rect 298753 66351 298787 66385
rect 298661 65807 298695 65841
rect 298753 65807 298787 65841
rect 298661 65263 298695 65297
rect 298753 65263 298787 65297
rect 298661 64719 298695 64753
rect 298753 64719 298787 64753
rect 298661 64175 298695 64209
rect 298753 64175 298787 64209
rect 298661 63631 298695 63665
rect 298753 63631 298787 63665
rect 298661 63087 298695 63121
rect 298753 63087 298787 63121
rect 298661 62543 298695 62577
rect 298753 62543 298787 62577
rect 298661 61999 298695 62033
rect 298753 61999 298787 62033
rect 298661 61455 298695 61489
rect 298753 61455 298787 61489
rect 298661 60911 298695 60945
rect 298753 60911 298787 60945
rect 298661 60367 298695 60401
rect 298753 60367 298787 60401
rect 298661 59823 298695 59857
rect 298753 59823 298787 59857
rect 298661 59279 298695 59313
rect 298753 59279 298787 59313
rect 298661 58735 298695 58769
rect 298753 58735 298787 58769
rect 298661 58191 298695 58225
rect 298753 58191 298787 58225
rect 298661 57647 298695 57681
rect 298753 57647 298787 57681
rect 298661 57103 298695 57137
rect 298753 57103 298787 57137
rect 298661 56559 298695 56593
rect 298753 56559 298787 56593
rect 298661 56015 298695 56049
rect 298753 56015 298787 56049
rect 298661 55471 298695 55505
rect 298753 55471 298787 55505
rect 298661 54927 298695 54961
rect 298753 54927 298787 54961
rect 298661 54383 298695 54417
rect 298753 54383 298787 54417
rect 298661 53839 298695 53873
rect 298753 53839 298787 53873
rect 298661 53295 298695 53329
rect 298753 53295 298787 53329
rect 298661 52751 298695 52785
rect 298753 52751 298787 52785
rect 298661 52207 298695 52241
rect 298753 52207 298787 52241
rect 298661 51663 298695 51697
rect 298753 51663 298787 51697
rect 298661 51119 298695 51153
rect 298753 51119 298787 51153
rect 298661 50575 298695 50609
rect 298753 50575 298787 50609
rect 298661 50031 298695 50065
rect 298753 50031 298787 50065
rect 298661 49487 298695 49521
rect 298753 49487 298787 49521
rect 298661 48943 298695 48977
rect 298753 48943 298787 48977
rect 298661 48399 298695 48433
rect 298753 48399 298787 48433
rect 298661 47855 298695 47889
rect 298753 47855 298787 47889
rect 298661 47311 298695 47345
rect 298753 47311 298787 47345
rect 298661 46767 298695 46801
rect 298753 46767 298787 46801
rect 298661 46223 298695 46257
rect 298753 46223 298787 46257
rect 298661 45679 298695 45713
rect 298753 45679 298787 45713
rect 298661 45135 298695 45169
rect 298753 45135 298787 45169
rect 298661 44591 298695 44625
rect 298753 44591 298787 44625
rect 298661 44047 298695 44081
rect 298753 44047 298787 44081
rect 298661 43503 298695 43537
rect 298753 43503 298787 43537
rect 298661 42959 298695 42993
rect 298753 42959 298787 42993
rect 298661 42415 298695 42449
rect 298753 42415 298787 42449
rect 298661 41871 298695 41905
rect 298753 41871 298787 41905
rect 298661 41327 298695 41361
rect 298753 41327 298787 41361
rect 298661 40783 298695 40817
rect 298753 40783 298787 40817
rect 298661 40239 298695 40273
rect 298753 40239 298787 40273
rect 298661 39695 298695 39729
rect 298753 39695 298787 39729
rect 298661 39151 298695 39185
rect 298753 39151 298787 39185
rect 298661 38607 298695 38641
rect 298753 38607 298787 38641
rect 298661 38063 298695 38097
rect 298753 38063 298787 38097
rect 298661 37519 298695 37553
rect 298753 37519 298787 37553
rect 298661 36975 298695 37009
rect 298753 36975 298787 37009
rect 298661 36431 298695 36465
rect 298753 36431 298787 36465
rect 298661 35887 298695 35921
rect 298753 35887 298787 35921
rect 298661 35343 298695 35377
rect 298753 35343 298787 35377
rect 298661 34799 298695 34833
rect 298753 34799 298787 34833
rect 298661 34255 298695 34289
rect 298753 34255 298787 34289
rect 298661 33711 298695 33745
rect 298753 33711 298787 33745
rect 298661 33167 298695 33201
rect 298753 33167 298787 33201
rect 298661 32623 298695 32657
rect 298753 32623 298787 32657
rect 298661 32079 298695 32113
rect 298753 32079 298787 32113
rect 298661 31535 298695 31569
rect 298753 31535 298787 31569
rect 298661 30991 298695 31025
rect 298753 30991 298787 31025
rect 298661 30447 298695 30481
rect 298753 30447 298787 30481
rect 298661 29903 298695 29937
rect 298753 29903 298787 29937
rect 298661 29359 298695 29393
rect 298753 29359 298787 29393
rect 298661 28815 298695 28849
rect 298753 28815 298787 28849
rect 298661 28271 298695 28305
rect 298753 28271 298787 28305
rect 298661 27727 298695 27761
rect 298753 27727 298787 27761
rect 298661 27183 298695 27217
rect 298753 27183 298787 27217
rect 298661 26639 298695 26673
rect 298753 26639 298787 26673
rect 298661 26095 298695 26129
rect 298753 26095 298787 26129
rect 298661 25551 298695 25585
rect 298753 25551 298787 25585
rect 298661 25007 298695 25041
rect 298753 25007 298787 25041
rect 298661 24463 298695 24497
rect 298753 24463 298787 24497
rect 298661 23919 298695 23953
rect 298753 23919 298787 23953
rect 298661 23375 298695 23409
rect 298753 23375 298787 23409
rect 298661 22831 298695 22865
rect 298753 22831 298787 22865
rect 298661 22287 298695 22321
rect 298753 22287 298787 22321
rect 298661 21743 298695 21777
rect 298753 21743 298787 21777
rect 298661 21199 298695 21233
rect 298753 21199 298787 21233
rect 298661 20655 298695 20689
rect 298753 20655 298787 20689
rect 298661 20111 298695 20145
rect 298753 20111 298787 20145
rect 298661 19567 298695 19601
rect 298753 19567 298787 19601
rect 298661 19023 298695 19057
rect 298753 19023 298787 19057
rect 298661 18479 298695 18513
rect 298753 18479 298787 18513
rect 298661 17935 298695 17969
rect 298753 17935 298787 17969
rect 298661 17391 298695 17425
rect 298753 17391 298787 17425
rect 298661 16847 298695 16881
rect 298753 16847 298787 16881
rect 298661 16303 298695 16337
rect 298753 16303 298787 16337
rect 298661 15759 298695 15793
rect 298753 15759 298787 15793
rect 298661 15215 298695 15249
rect 298753 15215 298787 15249
rect 298661 14671 298695 14705
rect 298753 14671 298787 14705
rect 298661 14127 298695 14161
rect 298753 14127 298787 14161
rect 298661 13583 298695 13617
rect 298753 13583 298787 13617
rect 298661 13039 298695 13073
rect 298753 13039 298787 13073
rect 298661 12495 298695 12529
rect 298753 12495 298787 12529
rect 298661 11951 298695 11985
rect 298753 11951 298787 11985
rect 298661 11407 298695 11441
rect 298753 11407 298787 11441
rect 298661 10863 298695 10897
rect 298753 10863 298787 10897
rect 298661 10319 298695 10353
rect 298753 10319 298787 10353
rect 298661 9775 298695 9809
rect 298753 9775 298787 9809
rect 298661 9231 298695 9265
rect 298753 9231 298787 9265
rect 298661 8687 298695 8721
rect 298753 8687 298787 8721
rect 298661 8143 298695 8177
rect 298753 8143 298787 8177
rect 298661 7599 298695 7633
rect 298753 7599 298787 7633
rect 298661 7055 298695 7089
rect 298753 7055 298787 7089
rect 298661 6511 298695 6545
rect 298753 6511 298787 6545
rect 298661 5967 298695 6001
rect 298753 5967 298787 6001
rect 298661 5423 298695 5457
rect 298753 5423 298787 5457
rect 298661 4879 298695 4913
rect 298753 4879 298787 4913
rect 298661 4335 298695 4369
rect 298753 4335 298787 4369
rect 298661 3791 298695 3825
rect 298753 3791 298787 3825
rect 298661 3247 298695 3281
rect 298753 3247 298787 3281
rect 298661 2703 298695 2737
rect 298753 2703 298787 2737
rect 298661 2159 298695 2193
rect 298753 2159 298787 2193
<< obsli1 >>
rect 1340 2159 298660 297585
<< metal1 >>
rect 1104 297585 1340 297616
rect 1104 297551 1133 297585
rect 1167 297551 1225 297585
rect 1259 297551 1317 297585
rect 1104 297520 1340 297551
rect 1104 297041 1340 297072
rect 1104 297007 1133 297041
rect 1167 297007 1225 297041
rect 1259 297007 1317 297041
rect 1104 296976 1340 297007
rect 1104 296497 1340 296528
rect 1104 296463 1133 296497
rect 1167 296463 1225 296497
rect 1259 296463 1317 296497
rect 1104 296432 1340 296463
rect 1104 295953 1340 295984
rect 1104 295919 1133 295953
rect 1167 295919 1225 295953
rect 1259 295919 1317 295953
rect 1104 295888 1340 295919
rect 1104 295409 1340 295440
rect 1104 295375 1133 295409
rect 1167 295375 1225 295409
rect 1259 295375 1317 295409
rect 1104 295344 1340 295375
rect 1104 294865 1340 294896
rect 1104 294831 1133 294865
rect 1167 294831 1225 294865
rect 1259 294831 1317 294865
rect 1104 294800 1340 294831
rect 1104 294321 1340 294352
rect 1104 294287 1133 294321
rect 1167 294287 1225 294321
rect 1259 294287 1317 294321
rect 1104 294256 1340 294287
rect 1104 293777 1340 293808
rect 1104 293743 1133 293777
rect 1167 293743 1225 293777
rect 1259 293743 1317 293777
rect 1104 293712 1340 293743
rect 1104 293233 1340 293264
rect 1104 293199 1133 293233
rect 1167 293199 1225 293233
rect 1259 293199 1317 293233
rect 1104 293168 1340 293199
rect 1104 292689 1340 292720
rect 1104 292655 1133 292689
rect 1167 292655 1225 292689
rect 1259 292655 1317 292689
rect 1104 292624 1340 292655
rect 1104 292145 1340 292176
rect 1104 292111 1133 292145
rect 1167 292111 1225 292145
rect 1259 292111 1317 292145
rect 1104 292080 1340 292111
rect 1104 291601 1340 291632
rect 1104 291567 1133 291601
rect 1167 291567 1225 291601
rect 1259 291567 1317 291601
rect 1104 291536 1340 291567
rect 1104 291057 1340 291088
rect 1104 291023 1133 291057
rect 1167 291023 1225 291057
rect 1259 291023 1317 291057
rect 1104 290992 1340 291023
rect 1104 290513 1340 290544
rect 1104 290479 1133 290513
rect 1167 290479 1225 290513
rect 1259 290479 1317 290513
rect 1104 290448 1340 290479
rect 1104 289969 1340 290000
rect 1104 289935 1133 289969
rect 1167 289935 1225 289969
rect 1259 289935 1317 289969
rect 1104 289904 1340 289935
rect 1104 289425 1340 289456
rect 1104 289391 1133 289425
rect 1167 289391 1225 289425
rect 1259 289391 1317 289425
rect 1104 289360 1340 289391
rect 1104 288881 1340 288912
rect 1104 288847 1133 288881
rect 1167 288847 1225 288881
rect 1259 288847 1317 288881
rect 1104 288816 1340 288847
rect 1104 288337 1340 288368
rect 1104 288303 1133 288337
rect 1167 288303 1225 288337
rect 1259 288303 1317 288337
rect 1104 288272 1340 288303
rect 1104 287793 1340 287824
rect 1104 287759 1133 287793
rect 1167 287759 1225 287793
rect 1259 287759 1317 287793
rect 1104 287728 1340 287759
rect 1104 287249 1340 287280
rect 1104 287215 1133 287249
rect 1167 287215 1225 287249
rect 1259 287215 1317 287249
rect 1104 287184 1340 287215
rect 1104 286705 1340 286736
rect 1104 286671 1133 286705
rect 1167 286671 1225 286705
rect 1259 286671 1317 286705
rect 1104 286640 1340 286671
rect 1104 286161 1340 286192
rect 1104 286127 1133 286161
rect 1167 286127 1225 286161
rect 1259 286127 1317 286161
rect 1104 286096 1340 286127
rect 1104 285617 1340 285648
rect 1104 285583 1133 285617
rect 1167 285583 1225 285617
rect 1259 285583 1317 285617
rect 1104 285552 1340 285583
rect 1104 285073 1340 285104
rect 1104 285039 1133 285073
rect 1167 285039 1225 285073
rect 1259 285039 1317 285073
rect 1104 285008 1340 285039
rect 1104 284529 1340 284560
rect 1104 284495 1133 284529
rect 1167 284495 1225 284529
rect 1259 284495 1317 284529
rect 1104 284464 1340 284495
rect 1104 283985 1340 284016
rect 1104 283951 1133 283985
rect 1167 283951 1225 283985
rect 1259 283951 1317 283985
rect 1104 283920 1340 283951
rect 1104 283441 1340 283472
rect 1104 283407 1133 283441
rect 1167 283407 1225 283441
rect 1259 283407 1317 283441
rect 1104 283376 1340 283407
rect 1104 282897 1340 282928
rect 1104 282863 1133 282897
rect 1167 282863 1225 282897
rect 1259 282863 1317 282897
rect 1104 282832 1340 282863
rect 1104 282353 1340 282384
rect 1104 282319 1133 282353
rect 1167 282319 1225 282353
rect 1259 282319 1317 282353
rect 1104 282288 1340 282319
rect 1104 281809 1340 281840
rect 1104 281775 1133 281809
rect 1167 281775 1225 281809
rect 1259 281775 1317 281809
rect 1104 281744 1340 281775
rect 1104 281265 1340 281296
rect 1104 281231 1133 281265
rect 1167 281231 1225 281265
rect 1259 281231 1317 281265
rect 1104 281200 1340 281231
rect 1104 280721 1340 280752
rect 1104 280687 1133 280721
rect 1167 280687 1225 280721
rect 1259 280687 1317 280721
rect 1104 280656 1340 280687
rect 1104 280177 1340 280208
rect 1104 280143 1133 280177
rect 1167 280143 1225 280177
rect 1259 280143 1317 280177
rect 1104 280112 1340 280143
rect 1104 279633 1340 279664
rect 1104 279599 1133 279633
rect 1167 279599 1225 279633
rect 1259 279599 1317 279633
rect 1104 279568 1340 279599
rect 1104 279089 1340 279120
rect 1104 279055 1133 279089
rect 1167 279055 1225 279089
rect 1259 279055 1317 279089
rect 1104 279024 1340 279055
rect 1104 278545 1340 278576
rect 1104 278511 1133 278545
rect 1167 278511 1225 278545
rect 1259 278511 1317 278545
rect 1104 278480 1340 278511
rect 1104 278001 1340 278032
rect 1104 277967 1133 278001
rect 1167 277967 1225 278001
rect 1259 277967 1317 278001
rect 1104 277936 1340 277967
rect 1104 277457 1340 277488
rect 1104 277423 1133 277457
rect 1167 277423 1225 277457
rect 1259 277423 1317 277457
rect 1104 277392 1340 277423
rect 1104 276913 1340 276944
rect 1104 276879 1133 276913
rect 1167 276879 1225 276913
rect 1259 276879 1317 276913
rect 1104 276848 1340 276879
rect 1104 276369 1340 276400
rect 1104 276335 1133 276369
rect 1167 276335 1225 276369
rect 1259 276335 1317 276369
rect 1104 276304 1340 276335
rect 1104 275825 1340 275856
rect 1104 275791 1133 275825
rect 1167 275791 1225 275825
rect 1259 275791 1317 275825
rect 1104 275760 1340 275791
rect 1104 275281 1340 275312
rect 1104 275247 1133 275281
rect 1167 275247 1225 275281
rect 1259 275247 1317 275281
rect 1104 275216 1340 275247
rect 1104 274737 1340 274768
rect 1104 274703 1133 274737
rect 1167 274703 1225 274737
rect 1259 274703 1317 274737
rect 1104 274672 1340 274703
rect 1104 274193 1340 274224
rect 1104 274159 1133 274193
rect 1167 274159 1225 274193
rect 1259 274159 1317 274193
rect 1104 274128 1340 274159
rect 1104 273649 1340 273680
rect 1104 273615 1133 273649
rect 1167 273615 1225 273649
rect 1259 273615 1317 273649
rect 1104 273584 1340 273615
rect 1104 273105 1340 273136
rect 1104 273071 1133 273105
rect 1167 273071 1225 273105
rect 1259 273071 1317 273105
rect 1104 273040 1340 273071
rect 1104 272561 1340 272592
rect 1104 272527 1133 272561
rect 1167 272527 1225 272561
rect 1259 272527 1317 272561
rect 1104 272496 1340 272527
rect 1104 272017 1340 272048
rect 1104 271983 1133 272017
rect 1167 271983 1225 272017
rect 1259 271983 1317 272017
rect 1104 271952 1340 271983
rect 1104 271473 1340 271504
rect 1104 271439 1133 271473
rect 1167 271439 1225 271473
rect 1259 271439 1317 271473
rect 1104 271408 1340 271439
rect 1104 270929 1340 270960
rect 1104 270895 1133 270929
rect 1167 270895 1225 270929
rect 1259 270895 1317 270929
rect 1104 270864 1340 270895
rect 1104 270385 1340 270416
rect 1104 270351 1133 270385
rect 1167 270351 1225 270385
rect 1259 270351 1317 270385
rect 1104 270320 1340 270351
rect 1104 269841 1340 269872
rect 1104 269807 1133 269841
rect 1167 269807 1225 269841
rect 1259 269807 1317 269841
rect 1104 269776 1340 269807
rect 1104 269297 1340 269328
rect 1104 269263 1133 269297
rect 1167 269263 1225 269297
rect 1259 269263 1317 269297
rect 1104 269232 1340 269263
rect 1104 268753 1340 268784
rect 1104 268719 1133 268753
rect 1167 268719 1225 268753
rect 1259 268719 1317 268753
rect 1104 268688 1340 268719
rect 1104 268209 1340 268240
rect 1104 268175 1133 268209
rect 1167 268175 1225 268209
rect 1259 268175 1317 268209
rect 1104 268144 1340 268175
rect 1104 267665 1340 267696
rect 1104 267631 1133 267665
rect 1167 267631 1225 267665
rect 1259 267631 1317 267665
rect 1104 267600 1340 267631
rect 1104 267121 1340 267152
rect 1104 267087 1133 267121
rect 1167 267087 1225 267121
rect 1259 267087 1317 267121
rect 1104 267056 1340 267087
rect 1104 266577 1340 266608
rect 1104 266543 1133 266577
rect 1167 266543 1225 266577
rect 1259 266543 1317 266577
rect 1104 266512 1340 266543
rect 1104 266033 1340 266064
rect 1104 265999 1133 266033
rect 1167 265999 1225 266033
rect 1259 265999 1317 266033
rect 1104 265968 1340 265999
rect 1104 265489 1340 265520
rect 1104 265455 1133 265489
rect 1167 265455 1225 265489
rect 1259 265455 1317 265489
rect 1104 265424 1340 265455
rect 1104 264945 1340 264976
rect 1104 264911 1133 264945
rect 1167 264911 1225 264945
rect 1259 264911 1317 264945
rect 1104 264880 1340 264911
rect 1104 264401 1340 264432
rect 1104 264367 1133 264401
rect 1167 264367 1225 264401
rect 1259 264367 1317 264401
rect 1104 264336 1340 264367
rect 1104 263857 1340 263888
rect 1104 263823 1133 263857
rect 1167 263823 1225 263857
rect 1259 263823 1317 263857
rect 1104 263792 1340 263823
rect 1104 263313 1340 263344
rect 1104 263279 1133 263313
rect 1167 263279 1225 263313
rect 1259 263279 1317 263313
rect 1104 263248 1340 263279
rect 1104 262769 1340 262800
rect 1104 262735 1133 262769
rect 1167 262735 1225 262769
rect 1259 262735 1317 262769
rect 1104 262704 1340 262735
rect 1104 262225 1340 262256
rect 1104 262191 1133 262225
rect 1167 262191 1225 262225
rect 1259 262191 1317 262225
rect 1104 262160 1340 262191
rect 1104 261681 1340 261712
rect 1104 261647 1133 261681
rect 1167 261647 1225 261681
rect 1259 261647 1317 261681
rect 1104 261616 1340 261647
rect 1104 261137 1340 261168
rect 1104 261103 1133 261137
rect 1167 261103 1225 261137
rect 1259 261103 1317 261137
rect 1104 261072 1340 261103
rect 1104 260593 1340 260624
rect 1104 260559 1133 260593
rect 1167 260559 1225 260593
rect 1259 260559 1317 260593
rect 1104 260528 1340 260559
rect 1104 260049 1340 260080
rect 1104 260015 1133 260049
rect 1167 260015 1225 260049
rect 1259 260015 1317 260049
rect 1104 259984 1340 260015
rect 1104 259505 1340 259536
rect 1104 259471 1133 259505
rect 1167 259471 1225 259505
rect 1259 259471 1317 259505
rect 1104 259440 1340 259471
rect 1104 258961 1340 258992
rect 1104 258927 1133 258961
rect 1167 258927 1225 258961
rect 1259 258927 1317 258961
rect 1104 258896 1340 258927
rect 1104 258417 1340 258448
rect 1104 258383 1133 258417
rect 1167 258383 1225 258417
rect 1259 258383 1317 258417
rect 1104 258352 1340 258383
rect 1104 257873 1340 257904
rect 1104 257839 1133 257873
rect 1167 257839 1225 257873
rect 1259 257839 1317 257873
rect 1104 257808 1340 257839
rect 1104 257329 1340 257360
rect 1104 257295 1133 257329
rect 1167 257295 1225 257329
rect 1259 257295 1317 257329
rect 1104 257264 1340 257295
rect 1104 256785 1340 256816
rect 1104 256751 1133 256785
rect 1167 256751 1225 256785
rect 1259 256751 1317 256785
rect 1104 256720 1340 256751
rect 1104 256241 1340 256272
rect 1104 256207 1133 256241
rect 1167 256207 1225 256241
rect 1259 256207 1317 256241
rect 1104 256176 1340 256207
rect 1104 255697 1340 255728
rect 1104 255663 1133 255697
rect 1167 255663 1225 255697
rect 1259 255663 1317 255697
rect 1104 255632 1340 255663
rect 1104 255153 1340 255184
rect 1104 255119 1133 255153
rect 1167 255119 1225 255153
rect 1259 255119 1317 255153
rect 1104 255088 1340 255119
rect 1104 254609 1340 254640
rect 1104 254575 1133 254609
rect 1167 254575 1225 254609
rect 1259 254575 1317 254609
rect 1104 254544 1340 254575
rect 1104 254065 1340 254096
rect 1104 254031 1133 254065
rect 1167 254031 1225 254065
rect 1259 254031 1317 254065
rect 1104 254000 1340 254031
rect 1104 253521 1340 253552
rect 1104 253487 1133 253521
rect 1167 253487 1225 253521
rect 1259 253487 1317 253521
rect 1104 253456 1340 253487
rect 1104 252977 1340 253008
rect 1104 252943 1133 252977
rect 1167 252943 1225 252977
rect 1259 252943 1317 252977
rect 1104 252912 1340 252943
rect 1104 252433 1340 252464
rect 1104 252399 1133 252433
rect 1167 252399 1225 252433
rect 1259 252399 1317 252433
rect 1104 252368 1340 252399
rect 1104 251889 1340 251920
rect 1104 251855 1133 251889
rect 1167 251855 1225 251889
rect 1259 251855 1317 251889
rect 1104 251824 1340 251855
rect 1104 251345 1340 251376
rect 1104 251311 1133 251345
rect 1167 251311 1225 251345
rect 1259 251311 1317 251345
rect 1104 251280 1340 251311
rect 1104 250801 1340 250832
rect 1104 250767 1133 250801
rect 1167 250767 1225 250801
rect 1259 250767 1317 250801
rect 1104 250736 1340 250767
rect 1104 250257 1340 250288
rect 1104 250223 1133 250257
rect 1167 250223 1225 250257
rect 1259 250223 1317 250257
rect 1104 250192 1340 250223
rect 1104 249713 1340 249744
rect 1104 249679 1133 249713
rect 1167 249679 1225 249713
rect 1259 249679 1317 249713
rect 1104 249648 1340 249679
rect 1104 249169 1340 249200
rect 1104 249135 1133 249169
rect 1167 249135 1225 249169
rect 1259 249135 1317 249169
rect 1104 249104 1340 249135
rect 1104 248625 1340 248656
rect 1104 248591 1133 248625
rect 1167 248591 1225 248625
rect 1259 248591 1317 248625
rect 1104 248560 1340 248591
rect 1104 248081 1340 248112
rect 1104 248047 1133 248081
rect 1167 248047 1225 248081
rect 1259 248047 1317 248081
rect 1104 248016 1340 248047
rect 1104 247537 1340 247568
rect 1104 247503 1133 247537
rect 1167 247503 1225 247537
rect 1259 247503 1317 247537
rect 1104 247472 1340 247503
rect 1104 246993 1340 247024
rect 1104 246959 1133 246993
rect 1167 246959 1225 246993
rect 1259 246959 1317 246993
rect 1104 246928 1340 246959
rect 1104 246449 1340 246480
rect 1104 246415 1133 246449
rect 1167 246415 1225 246449
rect 1259 246415 1317 246449
rect 1104 246384 1340 246415
rect 1104 245905 1340 245936
rect 1104 245871 1133 245905
rect 1167 245871 1225 245905
rect 1259 245871 1317 245905
rect 1104 245840 1340 245871
rect 1104 245361 1340 245392
rect 1104 245327 1133 245361
rect 1167 245327 1225 245361
rect 1259 245327 1317 245361
rect 1104 245296 1340 245327
rect 1104 244817 1340 244848
rect 1104 244783 1133 244817
rect 1167 244783 1225 244817
rect 1259 244783 1317 244817
rect 1104 244752 1340 244783
rect 1104 244273 1340 244304
rect 1104 244239 1133 244273
rect 1167 244239 1225 244273
rect 1259 244239 1317 244273
rect 1104 244208 1340 244239
rect 1104 243729 1340 243760
rect 1104 243695 1133 243729
rect 1167 243695 1225 243729
rect 1259 243695 1317 243729
rect 1104 243664 1340 243695
rect 1104 243185 1340 243216
rect 1104 243151 1133 243185
rect 1167 243151 1225 243185
rect 1259 243151 1317 243185
rect 1104 243120 1340 243151
rect 1104 242641 1340 242672
rect 1104 242607 1133 242641
rect 1167 242607 1225 242641
rect 1259 242607 1317 242641
rect 1104 242576 1340 242607
rect 1104 242097 1340 242128
rect 1104 242063 1133 242097
rect 1167 242063 1225 242097
rect 1259 242063 1317 242097
rect 1104 242032 1340 242063
rect 1104 241553 1340 241584
rect 1104 241519 1133 241553
rect 1167 241519 1225 241553
rect 1259 241519 1317 241553
rect 1104 241488 1340 241519
rect 1104 241009 1340 241040
rect 1104 240975 1133 241009
rect 1167 240975 1225 241009
rect 1259 240975 1317 241009
rect 1104 240944 1340 240975
rect 1104 240465 1340 240496
rect 1104 240431 1133 240465
rect 1167 240431 1225 240465
rect 1259 240431 1317 240465
rect 1104 240400 1340 240431
rect 1104 239921 1340 239952
rect 1104 239887 1133 239921
rect 1167 239887 1225 239921
rect 1259 239887 1317 239921
rect 1104 239856 1340 239887
rect 1104 239377 1340 239408
rect 1104 239343 1133 239377
rect 1167 239343 1225 239377
rect 1259 239343 1317 239377
rect 1104 239312 1340 239343
rect 1104 238833 1340 238864
rect 1104 238799 1133 238833
rect 1167 238799 1225 238833
rect 1259 238799 1317 238833
rect 1104 238768 1340 238799
rect 1104 238289 1340 238320
rect 1104 238255 1133 238289
rect 1167 238255 1225 238289
rect 1259 238255 1317 238289
rect 1104 238224 1340 238255
rect 1104 237745 1340 237776
rect 1104 237711 1133 237745
rect 1167 237711 1225 237745
rect 1259 237711 1317 237745
rect 1104 237680 1340 237711
rect 1104 237201 1340 237232
rect 1104 237167 1133 237201
rect 1167 237167 1225 237201
rect 1259 237167 1317 237201
rect 1104 237136 1340 237167
rect 1104 236657 1340 236688
rect 1104 236623 1133 236657
rect 1167 236623 1225 236657
rect 1259 236623 1317 236657
rect 1104 236592 1340 236623
rect 1104 236113 1340 236144
rect 1104 236079 1133 236113
rect 1167 236079 1225 236113
rect 1259 236079 1317 236113
rect 1104 236048 1340 236079
rect 1104 235569 1340 235600
rect 1104 235535 1133 235569
rect 1167 235535 1225 235569
rect 1259 235535 1317 235569
rect 1104 235504 1340 235535
rect 1104 235025 1340 235056
rect 1104 234991 1133 235025
rect 1167 234991 1225 235025
rect 1259 234991 1317 235025
rect 1104 234960 1340 234991
rect 1104 234481 1340 234512
rect 1104 234447 1133 234481
rect 1167 234447 1225 234481
rect 1259 234447 1317 234481
rect 1104 234416 1340 234447
rect 1104 233937 1340 233968
rect 1104 233903 1133 233937
rect 1167 233903 1225 233937
rect 1259 233903 1317 233937
rect 1104 233872 1340 233903
rect 1104 233393 1340 233424
rect 1104 233359 1133 233393
rect 1167 233359 1225 233393
rect 1259 233359 1317 233393
rect 1104 233328 1340 233359
rect 1104 232849 1340 232880
rect 1104 232815 1133 232849
rect 1167 232815 1225 232849
rect 1259 232815 1317 232849
rect 1104 232784 1340 232815
rect 1104 232305 1340 232336
rect 1104 232271 1133 232305
rect 1167 232271 1225 232305
rect 1259 232271 1317 232305
rect 1104 232240 1340 232271
rect 1104 231761 1340 231792
rect 1104 231727 1133 231761
rect 1167 231727 1225 231761
rect 1259 231727 1317 231761
rect 1104 231696 1340 231727
rect 1104 231217 1340 231248
rect 1104 231183 1133 231217
rect 1167 231183 1225 231217
rect 1259 231183 1317 231217
rect 1104 231152 1340 231183
rect 1104 230673 1340 230704
rect 1104 230639 1133 230673
rect 1167 230639 1225 230673
rect 1259 230639 1317 230673
rect 1104 230608 1340 230639
rect 1104 230129 1340 230160
rect 1104 230095 1133 230129
rect 1167 230095 1225 230129
rect 1259 230095 1317 230129
rect 1104 230064 1340 230095
rect 1104 229585 1340 229616
rect 1104 229551 1133 229585
rect 1167 229551 1225 229585
rect 1259 229551 1317 229585
rect 1104 229520 1340 229551
rect 1104 229041 1340 229072
rect 1104 229007 1133 229041
rect 1167 229007 1225 229041
rect 1259 229007 1317 229041
rect 1104 228976 1340 229007
rect 1104 228497 1340 228528
rect 1104 228463 1133 228497
rect 1167 228463 1225 228497
rect 1259 228463 1317 228497
rect 1104 228432 1340 228463
rect 1104 227953 1340 227984
rect 1104 227919 1133 227953
rect 1167 227919 1225 227953
rect 1259 227919 1317 227953
rect 1104 227888 1340 227919
rect 1104 227409 1340 227440
rect 1104 227375 1133 227409
rect 1167 227375 1225 227409
rect 1259 227375 1317 227409
rect 1104 227344 1340 227375
rect 1104 226865 1340 226896
rect 1104 226831 1133 226865
rect 1167 226831 1225 226865
rect 1259 226831 1317 226865
rect 1104 226800 1340 226831
rect 1104 226321 1340 226352
rect 1104 226287 1133 226321
rect 1167 226287 1225 226321
rect 1259 226287 1317 226321
rect 1104 226256 1340 226287
rect 1104 225777 1340 225808
rect 1104 225743 1133 225777
rect 1167 225743 1225 225777
rect 1259 225743 1317 225777
rect 1104 225712 1340 225743
rect 1104 225233 1340 225264
rect 1104 225199 1133 225233
rect 1167 225199 1225 225233
rect 1259 225199 1317 225233
rect 1104 225168 1340 225199
rect 1104 224689 1340 224720
rect 1104 224655 1133 224689
rect 1167 224655 1225 224689
rect 1259 224655 1317 224689
rect 1104 224624 1340 224655
rect 1104 224145 1340 224176
rect 1104 224111 1133 224145
rect 1167 224111 1225 224145
rect 1259 224111 1317 224145
rect 1104 224080 1340 224111
rect 1104 223601 1340 223632
rect 1104 223567 1133 223601
rect 1167 223567 1225 223601
rect 1259 223567 1317 223601
rect 1104 223536 1340 223567
rect 1104 223057 1340 223088
rect 1104 223023 1133 223057
rect 1167 223023 1225 223057
rect 1259 223023 1317 223057
rect 1104 222992 1340 223023
rect 1104 222513 1340 222544
rect 1104 222479 1133 222513
rect 1167 222479 1225 222513
rect 1259 222479 1317 222513
rect 1104 222448 1340 222479
rect 1104 221969 1340 222000
rect 1104 221935 1133 221969
rect 1167 221935 1225 221969
rect 1259 221935 1317 221969
rect 1104 221904 1340 221935
rect 1104 221425 1340 221456
rect 1104 221391 1133 221425
rect 1167 221391 1225 221425
rect 1259 221391 1317 221425
rect 1104 221360 1340 221391
rect 1104 220881 1340 220912
rect 1104 220847 1133 220881
rect 1167 220847 1225 220881
rect 1259 220847 1317 220881
rect 1104 220816 1340 220847
rect 1104 220337 1340 220368
rect 1104 220303 1133 220337
rect 1167 220303 1225 220337
rect 1259 220303 1317 220337
rect 1104 220272 1340 220303
rect 1104 219793 1340 219824
rect 1104 219759 1133 219793
rect 1167 219759 1225 219793
rect 1259 219759 1317 219793
rect 1104 219728 1340 219759
rect 1104 219249 1340 219280
rect 1104 219215 1133 219249
rect 1167 219215 1225 219249
rect 1259 219215 1317 219249
rect 1104 219184 1340 219215
rect 1104 218705 1340 218736
rect 1104 218671 1133 218705
rect 1167 218671 1225 218705
rect 1259 218671 1317 218705
rect 1104 218640 1340 218671
rect 1104 218161 1340 218192
rect 1104 218127 1133 218161
rect 1167 218127 1225 218161
rect 1259 218127 1317 218161
rect 1104 218096 1340 218127
rect 1104 217617 1340 217648
rect 1104 217583 1133 217617
rect 1167 217583 1225 217617
rect 1259 217583 1317 217617
rect 1104 217552 1340 217583
rect 1104 217073 1340 217104
rect 1104 217039 1133 217073
rect 1167 217039 1225 217073
rect 1259 217039 1317 217073
rect 1104 217008 1340 217039
rect 1104 216529 1340 216560
rect 1104 216495 1133 216529
rect 1167 216495 1225 216529
rect 1259 216495 1317 216529
rect 1104 216464 1340 216495
rect 1104 215985 1340 216016
rect 1104 215951 1133 215985
rect 1167 215951 1225 215985
rect 1259 215951 1317 215985
rect 1104 215920 1340 215951
rect 1104 215441 1340 215472
rect 1104 215407 1133 215441
rect 1167 215407 1225 215441
rect 1259 215407 1317 215441
rect 1104 215376 1340 215407
rect 1104 214897 1340 214928
rect 1104 214863 1133 214897
rect 1167 214863 1225 214897
rect 1259 214863 1317 214897
rect 1104 214832 1340 214863
rect 1104 214353 1340 214384
rect 1104 214319 1133 214353
rect 1167 214319 1225 214353
rect 1259 214319 1317 214353
rect 1104 214288 1340 214319
rect 1104 213809 1340 213840
rect 1104 213775 1133 213809
rect 1167 213775 1225 213809
rect 1259 213775 1317 213809
rect 1104 213744 1340 213775
rect 1104 213265 1340 213296
rect 1104 213231 1133 213265
rect 1167 213231 1225 213265
rect 1259 213231 1317 213265
rect 1104 213200 1340 213231
rect 1104 212721 1340 212752
rect 1104 212687 1133 212721
rect 1167 212687 1225 212721
rect 1259 212687 1317 212721
rect 1104 212656 1340 212687
rect 1104 212177 1340 212208
rect 1104 212143 1133 212177
rect 1167 212143 1225 212177
rect 1259 212143 1317 212177
rect 1104 212112 1340 212143
rect 1104 211633 1340 211664
rect 1104 211599 1133 211633
rect 1167 211599 1225 211633
rect 1259 211599 1317 211633
rect 1104 211568 1340 211599
rect 1104 211089 1340 211120
rect 1104 211055 1133 211089
rect 1167 211055 1225 211089
rect 1259 211055 1317 211089
rect 1104 211024 1340 211055
rect 1104 210545 1340 210576
rect 1104 210511 1133 210545
rect 1167 210511 1225 210545
rect 1259 210511 1317 210545
rect 1104 210480 1340 210511
rect 1104 210001 1340 210032
rect 1104 209967 1133 210001
rect 1167 209967 1225 210001
rect 1259 209967 1317 210001
rect 1104 209936 1340 209967
rect 1104 209457 1340 209488
rect 1104 209423 1133 209457
rect 1167 209423 1225 209457
rect 1259 209423 1317 209457
rect 1104 209392 1340 209423
rect 1104 208913 1340 208944
rect 1104 208879 1133 208913
rect 1167 208879 1225 208913
rect 1259 208879 1317 208913
rect 1104 208848 1340 208879
rect 1104 208369 1340 208400
rect 1104 208335 1133 208369
rect 1167 208335 1225 208369
rect 1259 208335 1317 208369
rect 1104 208304 1340 208335
rect 1104 207825 1340 207856
rect 1104 207791 1133 207825
rect 1167 207791 1225 207825
rect 1259 207791 1317 207825
rect 1104 207760 1340 207791
rect 1104 207281 1340 207312
rect 1104 207247 1133 207281
rect 1167 207247 1225 207281
rect 1259 207247 1317 207281
rect 1104 207216 1340 207247
rect 1104 206737 1340 206768
rect 1104 206703 1133 206737
rect 1167 206703 1225 206737
rect 1259 206703 1317 206737
rect 1104 206672 1340 206703
rect 1104 206193 1340 206224
rect 1104 206159 1133 206193
rect 1167 206159 1225 206193
rect 1259 206159 1317 206193
rect 1104 206128 1340 206159
rect 1104 205649 1340 205680
rect 1104 205615 1133 205649
rect 1167 205615 1225 205649
rect 1259 205615 1317 205649
rect 1104 205584 1340 205615
rect 1104 205105 1340 205136
rect 1104 205071 1133 205105
rect 1167 205071 1225 205105
rect 1259 205071 1317 205105
rect 1104 205040 1340 205071
rect 1104 204561 1340 204592
rect 1104 204527 1133 204561
rect 1167 204527 1225 204561
rect 1259 204527 1317 204561
rect 1104 204496 1340 204527
rect 1104 204017 1340 204048
rect 1104 203983 1133 204017
rect 1167 203983 1225 204017
rect 1259 203983 1317 204017
rect 1104 203952 1340 203983
rect 1104 203473 1340 203504
rect 1104 203439 1133 203473
rect 1167 203439 1225 203473
rect 1259 203439 1317 203473
rect 1104 203408 1340 203439
rect 1104 202929 1340 202960
rect 1104 202895 1133 202929
rect 1167 202895 1225 202929
rect 1259 202895 1317 202929
rect 1104 202864 1340 202895
rect 1104 202385 1340 202416
rect 1104 202351 1133 202385
rect 1167 202351 1225 202385
rect 1259 202351 1317 202385
rect 1104 202320 1340 202351
rect 1104 201841 1340 201872
rect 1104 201807 1133 201841
rect 1167 201807 1225 201841
rect 1259 201807 1317 201841
rect 1104 201776 1340 201807
rect 1104 201297 1340 201328
rect 1104 201263 1133 201297
rect 1167 201263 1225 201297
rect 1259 201263 1317 201297
rect 1104 201232 1340 201263
rect 1104 200753 1340 200784
rect 1104 200719 1133 200753
rect 1167 200719 1225 200753
rect 1259 200719 1317 200753
rect 1104 200688 1340 200719
rect 1104 200209 1340 200240
rect 1104 200175 1133 200209
rect 1167 200175 1225 200209
rect 1259 200175 1317 200209
rect 1104 200144 1340 200175
rect 1104 199665 1340 199696
rect 1104 199631 1133 199665
rect 1167 199631 1225 199665
rect 1259 199631 1317 199665
rect 1104 199600 1340 199631
rect 1104 199121 1340 199152
rect 1104 199087 1133 199121
rect 1167 199087 1225 199121
rect 1259 199087 1317 199121
rect 1104 199056 1340 199087
rect 1104 198577 1340 198608
rect 1104 198543 1133 198577
rect 1167 198543 1225 198577
rect 1259 198543 1317 198577
rect 1104 198512 1340 198543
rect 1104 198033 1340 198064
rect 1104 197999 1133 198033
rect 1167 197999 1225 198033
rect 1259 197999 1317 198033
rect 1104 197968 1340 197999
rect 1104 197489 1340 197520
rect 1104 197455 1133 197489
rect 1167 197455 1225 197489
rect 1259 197455 1317 197489
rect 1104 197424 1340 197455
rect 1104 196945 1340 196976
rect 1104 196911 1133 196945
rect 1167 196911 1225 196945
rect 1259 196911 1317 196945
rect 1104 196880 1340 196911
rect 1104 196401 1340 196432
rect 1104 196367 1133 196401
rect 1167 196367 1225 196401
rect 1259 196367 1317 196401
rect 1104 196336 1340 196367
rect 1104 195857 1340 195888
rect 1104 195823 1133 195857
rect 1167 195823 1225 195857
rect 1259 195823 1317 195857
rect 1104 195792 1340 195823
rect 1104 195313 1340 195344
rect 1104 195279 1133 195313
rect 1167 195279 1225 195313
rect 1259 195279 1317 195313
rect 1104 195248 1340 195279
rect 1104 194769 1340 194800
rect 1104 194735 1133 194769
rect 1167 194735 1225 194769
rect 1259 194735 1317 194769
rect 1104 194704 1340 194735
rect 1104 194225 1340 194256
rect 1104 194191 1133 194225
rect 1167 194191 1225 194225
rect 1259 194191 1317 194225
rect 1104 194160 1340 194191
rect 1104 193681 1340 193712
rect 1104 193647 1133 193681
rect 1167 193647 1225 193681
rect 1259 193647 1317 193681
rect 1104 193616 1340 193647
rect 1104 193137 1340 193168
rect 1104 193103 1133 193137
rect 1167 193103 1225 193137
rect 1259 193103 1317 193137
rect 1104 193072 1340 193103
rect 1104 192593 1340 192624
rect 1104 192559 1133 192593
rect 1167 192559 1225 192593
rect 1259 192559 1317 192593
rect 1104 192528 1340 192559
rect 1104 192049 1340 192080
rect 1104 192015 1133 192049
rect 1167 192015 1225 192049
rect 1259 192015 1317 192049
rect 1104 191984 1340 192015
rect 1104 191505 1340 191536
rect 1104 191471 1133 191505
rect 1167 191471 1225 191505
rect 1259 191471 1317 191505
rect 1104 191440 1340 191471
rect 1104 190961 1340 190992
rect 1104 190927 1133 190961
rect 1167 190927 1225 190961
rect 1259 190927 1317 190961
rect 1104 190896 1340 190927
rect 1104 190417 1340 190448
rect 1104 190383 1133 190417
rect 1167 190383 1225 190417
rect 1259 190383 1317 190417
rect 1104 190352 1340 190383
rect 1104 189873 1340 189904
rect 1104 189839 1133 189873
rect 1167 189839 1225 189873
rect 1259 189839 1317 189873
rect 1104 189808 1340 189839
rect 1104 189329 1340 189360
rect 1104 189295 1133 189329
rect 1167 189295 1225 189329
rect 1259 189295 1317 189329
rect 1104 189264 1340 189295
rect 1104 188785 1340 188816
rect 1104 188751 1133 188785
rect 1167 188751 1225 188785
rect 1259 188751 1317 188785
rect 1104 188720 1340 188751
rect 1104 188241 1340 188272
rect 1104 188207 1133 188241
rect 1167 188207 1225 188241
rect 1259 188207 1317 188241
rect 1104 188176 1340 188207
rect 1104 187697 1340 187728
rect 1104 187663 1133 187697
rect 1167 187663 1225 187697
rect 1259 187663 1317 187697
rect 1104 187632 1340 187663
rect 1104 187153 1340 187184
rect 1104 187119 1133 187153
rect 1167 187119 1225 187153
rect 1259 187119 1317 187153
rect 1104 187088 1340 187119
rect 1104 186609 1340 186640
rect 1104 186575 1133 186609
rect 1167 186575 1225 186609
rect 1259 186575 1317 186609
rect 1104 186544 1340 186575
rect 1104 186065 1340 186096
rect 1104 186031 1133 186065
rect 1167 186031 1225 186065
rect 1259 186031 1317 186065
rect 1104 186000 1340 186031
rect 1104 185521 1340 185552
rect 1104 185487 1133 185521
rect 1167 185487 1225 185521
rect 1259 185487 1317 185521
rect 1104 185456 1340 185487
rect 1104 184977 1340 185008
rect 1104 184943 1133 184977
rect 1167 184943 1225 184977
rect 1259 184943 1317 184977
rect 1104 184912 1340 184943
rect 1104 184433 1340 184464
rect 1104 184399 1133 184433
rect 1167 184399 1225 184433
rect 1259 184399 1317 184433
rect 1104 184368 1340 184399
rect 1104 183889 1340 183920
rect 1104 183855 1133 183889
rect 1167 183855 1225 183889
rect 1259 183855 1317 183889
rect 1104 183824 1340 183855
rect 1104 183345 1340 183376
rect 1104 183311 1133 183345
rect 1167 183311 1225 183345
rect 1259 183311 1317 183345
rect 1104 183280 1340 183311
rect 1104 182801 1340 182832
rect 1104 182767 1133 182801
rect 1167 182767 1225 182801
rect 1259 182767 1317 182801
rect 1104 182736 1340 182767
rect 1104 182257 1340 182288
rect 1104 182223 1133 182257
rect 1167 182223 1225 182257
rect 1259 182223 1317 182257
rect 1104 182192 1340 182223
rect 1104 181713 1340 181744
rect 1104 181679 1133 181713
rect 1167 181679 1225 181713
rect 1259 181679 1317 181713
rect 1104 181648 1340 181679
rect 1104 181169 1340 181200
rect 1104 181135 1133 181169
rect 1167 181135 1225 181169
rect 1259 181135 1317 181169
rect 1104 181104 1340 181135
rect 1104 180625 1340 180656
rect 1104 180591 1133 180625
rect 1167 180591 1225 180625
rect 1259 180591 1317 180625
rect 1104 180560 1340 180591
rect 1104 180081 1340 180112
rect 1104 180047 1133 180081
rect 1167 180047 1225 180081
rect 1259 180047 1317 180081
rect 1104 180016 1340 180047
rect 1104 179537 1340 179568
rect 1104 179503 1133 179537
rect 1167 179503 1225 179537
rect 1259 179503 1317 179537
rect 1104 179472 1340 179503
rect 1104 178993 1340 179024
rect 1104 178959 1133 178993
rect 1167 178959 1225 178993
rect 1259 178959 1317 178993
rect 1104 178928 1340 178959
rect 1104 178449 1340 178480
rect 1104 178415 1133 178449
rect 1167 178415 1225 178449
rect 1259 178415 1317 178449
rect 1104 178384 1340 178415
rect 1104 177905 1340 177936
rect 1104 177871 1133 177905
rect 1167 177871 1225 177905
rect 1259 177871 1317 177905
rect 1104 177840 1340 177871
rect 1104 177361 1340 177392
rect 1104 177327 1133 177361
rect 1167 177327 1225 177361
rect 1259 177327 1317 177361
rect 1104 177296 1340 177327
rect 1104 176817 1340 176848
rect 1104 176783 1133 176817
rect 1167 176783 1225 176817
rect 1259 176783 1317 176817
rect 1104 176752 1340 176783
rect 1104 176273 1340 176304
rect 1104 176239 1133 176273
rect 1167 176239 1225 176273
rect 1259 176239 1317 176273
rect 1104 176208 1340 176239
rect 1104 175729 1340 175760
rect 1104 175695 1133 175729
rect 1167 175695 1225 175729
rect 1259 175695 1317 175729
rect 1104 175664 1340 175695
rect 1104 175185 1340 175216
rect 1104 175151 1133 175185
rect 1167 175151 1225 175185
rect 1259 175151 1317 175185
rect 1104 175120 1340 175151
rect 1104 174641 1340 174672
rect 1104 174607 1133 174641
rect 1167 174607 1225 174641
rect 1259 174607 1317 174641
rect 1104 174576 1340 174607
rect 1104 174097 1340 174128
rect 1104 174063 1133 174097
rect 1167 174063 1225 174097
rect 1259 174063 1317 174097
rect 1104 174032 1340 174063
rect 1104 173553 1340 173584
rect 1104 173519 1133 173553
rect 1167 173519 1225 173553
rect 1259 173519 1317 173553
rect 1104 173488 1340 173519
rect 1104 173009 1340 173040
rect 1104 172975 1133 173009
rect 1167 172975 1225 173009
rect 1259 172975 1317 173009
rect 1104 172944 1340 172975
rect 1104 172465 1340 172496
rect 1104 172431 1133 172465
rect 1167 172431 1225 172465
rect 1259 172431 1317 172465
rect 1104 172400 1340 172431
rect 1104 171921 1340 171952
rect 1104 171887 1133 171921
rect 1167 171887 1225 171921
rect 1259 171887 1317 171921
rect 1104 171856 1340 171887
rect 1104 171377 1340 171408
rect 1104 171343 1133 171377
rect 1167 171343 1225 171377
rect 1259 171343 1317 171377
rect 1104 171312 1340 171343
rect 1104 170833 1340 170864
rect 1104 170799 1133 170833
rect 1167 170799 1225 170833
rect 1259 170799 1317 170833
rect 1104 170768 1340 170799
rect 1104 170289 1340 170320
rect 1104 170255 1133 170289
rect 1167 170255 1225 170289
rect 1259 170255 1317 170289
rect 1104 170224 1340 170255
rect 1104 169745 1340 169776
rect 1104 169711 1133 169745
rect 1167 169711 1225 169745
rect 1259 169711 1317 169745
rect 1104 169680 1340 169711
rect 1104 169201 1340 169232
rect 1104 169167 1133 169201
rect 1167 169167 1225 169201
rect 1259 169167 1317 169201
rect 1104 169136 1340 169167
rect 1104 168657 1340 168688
rect 1104 168623 1133 168657
rect 1167 168623 1225 168657
rect 1259 168623 1317 168657
rect 1104 168592 1340 168623
rect 1104 168113 1340 168144
rect 1104 168079 1133 168113
rect 1167 168079 1225 168113
rect 1259 168079 1317 168113
rect 1104 168048 1340 168079
rect 1104 167569 1340 167600
rect 1104 167535 1133 167569
rect 1167 167535 1225 167569
rect 1259 167535 1317 167569
rect 1104 167504 1340 167535
rect 1104 167025 1340 167056
rect 1104 166991 1133 167025
rect 1167 166991 1225 167025
rect 1259 166991 1317 167025
rect 1104 166960 1340 166991
rect 1104 166481 1340 166512
rect 1104 166447 1133 166481
rect 1167 166447 1225 166481
rect 1259 166447 1317 166481
rect 1104 166416 1340 166447
rect 1104 165937 1340 165968
rect 1104 165903 1133 165937
rect 1167 165903 1225 165937
rect 1259 165903 1317 165937
rect 1104 165872 1340 165903
rect 1104 165393 1340 165424
rect 1104 165359 1133 165393
rect 1167 165359 1225 165393
rect 1259 165359 1317 165393
rect 1104 165328 1340 165359
rect 1104 164849 1340 164880
rect 1104 164815 1133 164849
rect 1167 164815 1225 164849
rect 1259 164815 1317 164849
rect 1104 164784 1340 164815
rect 1104 164305 1340 164336
rect 1104 164271 1133 164305
rect 1167 164271 1225 164305
rect 1259 164271 1317 164305
rect 1104 164240 1340 164271
rect 1104 163761 1340 163792
rect 1104 163727 1133 163761
rect 1167 163727 1225 163761
rect 1259 163727 1317 163761
rect 1104 163696 1340 163727
rect 1104 163217 1340 163248
rect 1104 163183 1133 163217
rect 1167 163183 1225 163217
rect 1259 163183 1317 163217
rect 1104 163152 1340 163183
rect 1104 162673 1340 162704
rect 1104 162639 1133 162673
rect 1167 162639 1225 162673
rect 1259 162639 1317 162673
rect 1104 162608 1340 162639
rect 1104 162129 1340 162160
rect 1104 162095 1133 162129
rect 1167 162095 1225 162129
rect 1259 162095 1317 162129
rect 1104 162064 1340 162095
rect 1104 161585 1340 161616
rect 1104 161551 1133 161585
rect 1167 161551 1225 161585
rect 1259 161551 1317 161585
rect 1104 161520 1340 161551
rect 1104 161041 1340 161072
rect 1104 161007 1133 161041
rect 1167 161007 1225 161041
rect 1259 161007 1317 161041
rect 1104 160976 1340 161007
rect 1104 160497 1340 160528
rect 1104 160463 1133 160497
rect 1167 160463 1225 160497
rect 1259 160463 1317 160497
rect 1104 160432 1340 160463
rect 1104 159953 1340 159984
rect 1104 159919 1133 159953
rect 1167 159919 1225 159953
rect 1259 159919 1317 159953
rect 1104 159888 1340 159919
rect 1104 159409 1340 159440
rect 1104 159375 1133 159409
rect 1167 159375 1225 159409
rect 1259 159375 1317 159409
rect 1104 159344 1340 159375
rect 1104 158865 1340 158896
rect 1104 158831 1133 158865
rect 1167 158831 1225 158865
rect 1259 158831 1317 158865
rect 1104 158800 1340 158831
rect 1104 158321 1340 158352
rect 1104 158287 1133 158321
rect 1167 158287 1225 158321
rect 1259 158287 1317 158321
rect 1104 158256 1340 158287
rect 1104 157777 1340 157808
rect 1104 157743 1133 157777
rect 1167 157743 1225 157777
rect 1259 157743 1317 157777
rect 1104 157712 1340 157743
rect 1104 157233 1340 157264
rect 1104 157199 1133 157233
rect 1167 157199 1225 157233
rect 1259 157199 1317 157233
rect 1104 157168 1340 157199
rect 1104 156689 1340 156720
rect 1104 156655 1133 156689
rect 1167 156655 1225 156689
rect 1259 156655 1317 156689
rect 1104 156624 1340 156655
rect 1104 156145 1340 156176
rect 1104 156111 1133 156145
rect 1167 156111 1225 156145
rect 1259 156111 1317 156145
rect 1104 156080 1340 156111
rect 1104 155601 1340 155632
rect 1104 155567 1133 155601
rect 1167 155567 1225 155601
rect 1259 155567 1317 155601
rect 1104 155536 1340 155567
rect 1104 155057 1340 155088
rect 1104 155023 1133 155057
rect 1167 155023 1225 155057
rect 1259 155023 1317 155057
rect 1104 154992 1340 155023
rect 1104 154513 1340 154544
rect 1104 154479 1133 154513
rect 1167 154479 1225 154513
rect 1259 154479 1317 154513
rect 1104 154448 1340 154479
rect 1104 153969 1340 154000
rect 1104 153935 1133 153969
rect 1167 153935 1225 153969
rect 1259 153935 1317 153969
rect 1104 153904 1340 153935
rect 1104 153425 1340 153456
rect 1104 153391 1133 153425
rect 1167 153391 1225 153425
rect 1259 153391 1317 153425
rect 1104 153360 1340 153391
rect 1104 152881 1340 152912
rect 1104 152847 1133 152881
rect 1167 152847 1225 152881
rect 1259 152847 1317 152881
rect 1104 152816 1340 152847
rect 1104 152337 1340 152368
rect 1104 152303 1133 152337
rect 1167 152303 1225 152337
rect 1259 152303 1317 152337
rect 1104 152272 1340 152303
rect 1104 151793 1340 151824
rect 1104 151759 1133 151793
rect 1167 151759 1225 151793
rect 1259 151759 1317 151793
rect 1104 151728 1340 151759
rect 1104 151249 1340 151280
rect 1104 151215 1133 151249
rect 1167 151215 1225 151249
rect 1259 151215 1317 151249
rect 1104 151184 1340 151215
rect 1104 150705 1340 150736
rect 1104 150671 1133 150705
rect 1167 150671 1225 150705
rect 1259 150671 1317 150705
rect 1104 150640 1340 150671
rect 1104 150161 1340 150192
rect 1104 150127 1133 150161
rect 1167 150127 1225 150161
rect 1259 150127 1317 150161
rect 1104 150096 1340 150127
rect 1104 149617 1340 149648
rect 1104 149583 1133 149617
rect 1167 149583 1225 149617
rect 1259 149583 1317 149617
rect 1104 149552 1340 149583
rect 1104 149073 1340 149104
rect 1104 149039 1133 149073
rect 1167 149039 1225 149073
rect 1259 149039 1317 149073
rect 1104 149008 1340 149039
rect 1104 148529 1340 148560
rect 1104 148495 1133 148529
rect 1167 148495 1225 148529
rect 1259 148495 1317 148529
rect 1104 148464 1340 148495
rect 1104 147985 1340 148016
rect 1104 147951 1133 147985
rect 1167 147951 1225 147985
rect 1259 147951 1317 147985
rect 1104 147920 1340 147951
rect 1104 147441 1340 147472
rect 1104 147407 1133 147441
rect 1167 147407 1225 147441
rect 1259 147407 1317 147441
rect 1104 147376 1340 147407
rect 1104 146897 1340 146928
rect 1104 146863 1133 146897
rect 1167 146863 1225 146897
rect 1259 146863 1317 146897
rect 1104 146832 1340 146863
rect 1104 146353 1340 146384
rect 1104 146319 1133 146353
rect 1167 146319 1225 146353
rect 1259 146319 1317 146353
rect 1104 146288 1340 146319
rect 1104 145809 1340 145840
rect 1104 145775 1133 145809
rect 1167 145775 1225 145809
rect 1259 145775 1317 145809
rect 1104 145744 1340 145775
rect 1104 145265 1340 145296
rect 1104 145231 1133 145265
rect 1167 145231 1225 145265
rect 1259 145231 1317 145265
rect 1104 145200 1340 145231
rect 1104 144721 1340 144752
rect 1104 144687 1133 144721
rect 1167 144687 1225 144721
rect 1259 144687 1317 144721
rect 1104 144656 1340 144687
rect 1104 144177 1340 144208
rect 1104 144143 1133 144177
rect 1167 144143 1225 144177
rect 1259 144143 1317 144177
rect 1104 144112 1340 144143
rect 1104 143633 1340 143664
rect 1104 143599 1133 143633
rect 1167 143599 1225 143633
rect 1259 143599 1317 143633
rect 1104 143568 1340 143599
rect 1104 143089 1340 143120
rect 1104 143055 1133 143089
rect 1167 143055 1225 143089
rect 1259 143055 1317 143089
rect 1104 143024 1340 143055
rect 1104 142545 1340 142576
rect 1104 142511 1133 142545
rect 1167 142511 1225 142545
rect 1259 142511 1317 142545
rect 1104 142480 1340 142511
rect 1104 142001 1340 142032
rect 1104 141967 1133 142001
rect 1167 141967 1225 142001
rect 1259 141967 1317 142001
rect 1104 141936 1340 141967
rect 1104 141457 1340 141488
rect 1104 141423 1133 141457
rect 1167 141423 1225 141457
rect 1259 141423 1317 141457
rect 1104 141392 1340 141423
rect 1104 140913 1340 140944
rect 1104 140879 1133 140913
rect 1167 140879 1225 140913
rect 1259 140879 1317 140913
rect 1104 140848 1340 140879
rect 1104 140369 1340 140400
rect 1104 140335 1133 140369
rect 1167 140335 1225 140369
rect 1259 140335 1317 140369
rect 1104 140304 1340 140335
rect 1104 139825 1340 139856
rect 1104 139791 1133 139825
rect 1167 139791 1225 139825
rect 1259 139791 1317 139825
rect 1104 139760 1340 139791
rect 1104 139281 1340 139312
rect 1104 139247 1133 139281
rect 1167 139247 1225 139281
rect 1259 139247 1317 139281
rect 1104 139216 1340 139247
rect 1104 138737 1340 138768
rect 1104 138703 1133 138737
rect 1167 138703 1225 138737
rect 1259 138703 1317 138737
rect 1104 138672 1340 138703
rect 1104 138193 1340 138224
rect 1104 138159 1133 138193
rect 1167 138159 1225 138193
rect 1259 138159 1317 138193
rect 1104 138128 1340 138159
rect 1104 137649 1340 137680
rect 1104 137615 1133 137649
rect 1167 137615 1225 137649
rect 1259 137615 1317 137649
rect 1104 137584 1340 137615
rect 1104 137105 1340 137136
rect 1104 137071 1133 137105
rect 1167 137071 1225 137105
rect 1259 137071 1317 137105
rect 1104 137040 1340 137071
rect 1104 136561 1340 136592
rect 1104 136527 1133 136561
rect 1167 136527 1225 136561
rect 1259 136527 1317 136561
rect 1104 136496 1340 136527
rect 1104 136017 1340 136048
rect 1104 135983 1133 136017
rect 1167 135983 1225 136017
rect 1259 135983 1317 136017
rect 1104 135952 1340 135983
rect 1104 135473 1340 135504
rect 1104 135439 1133 135473
rect 1167 135439 1225 135473
rect 1259 135439 1317 135473
rect 1104 135408 1340 135439
rect 1104 134929 1340 134960
rect 1104 134895 1133 134929
rect 1167 134895 1225 134929
rect 1259 134895 1317 134929
rect 1104 134864 1340 134895
rect 1104 134385 1340 134416
rect 1104 134351 1133 134385
rect 1167 134351 1225 134385
rect 1259 134351 1317 134385
rect 1104 134320 1340 134351
rect 1104 133841 1340 133872
rect 1104 133807 1133 133841
rect 1167 133807 1225 133841
rect 1259 133807 1317 133841
rect 1104 133776 1340 133807
rect 1104 133297 1340 133328
rect 1104 133263 1133 133297
rect 1167 133263 1225 133297
rect 1259 133263 1317 133297
rect 1104 133232 1340 133263
rect 1104 132753 1340 132784
rect 1104 132719 1133 132753
rect 1167 132719 1225 132753
rect 1259 132719 1317 132753
rect 1104 132688 1340 132719
rect 1104 132209 1340 132240
rect 1104 132175 1133 132209
rect 1167 132175 1225 132209
rect 1259 132175 1317 132209
rect 1104 132144 1340 132175
rect 1104 131665 1340 131696
rect 1104 131631 1133 131665
rect 1167 131631 1225 131665
rect 1259 131631 1317 131665
rect 1104 131600 1340 131631
rect 1104 131121 1340 131152
rect 1104 131087 1133 131121
rect 1167 131087 1225 131121
rect 1259 131087 1317 131121
rect 1104 131056 1340 131087
rect 1104 130577 1340 130608
rect 1104 130543 1133 130577
rect 1167 130543 1225 130577
rect 1259 130543 1317 130577
rect 1104 130512 1340 130543
rect 1104 130033 1340 130064
rect 1104 129999 1133 130033
rect 1167 129999 1225 130033
rect 1259 129999 1317 130033
rect 1104 129968 1340 129999
rect 1104 129489 1340 129520
rect 1104 129455 1133 129489
rect 1167 129455 1225 129489
rect 1259 129455 1317 129489
rect 1104 129424 1340 129455
rect 1104 128945 1340 128976
rect 1104 128911 1133 128945
rect 1167 128911 1225 128945
rect 1259 128911 1317 128945
rect 1104 128880 1340 128911
rect 1104 128401 1340 128432
rect 1104 128367 1133 128401
rect 1167 128367 1225 128401
rect 1259 128367 1317 128401
rect 1104 128336 1340 128367
rect 1104 127857 1340 127888
rect 1104 127823 1133 127857
rect 1167 127823 1225 127857
rect 1259 127823 1317 127857
rect 1104 127792 1340 127823
rect 1104 127313 1340 127344
rect 1104 127279 1133 127313
rect 1167 127279 1225 127313
rect 1259 127279 1317 127313
rect 1104 127248 1340 127279
rect 1104 126769 1340 126800
rect 1104 126735 1133 126769
rect 1167 126735 1225 126769
rect 1259 126735 1317 126769
rect 1104 126704 1340 126735
rect 1104 126225 1340 126256
rect 1104 126191 1133 126225
rect 1167 126191 1225 126225
rect 1259 126191 1317 126225
rect 1104 126160 1340 126191
rect 1104 125681 1340 125712
rect 1104 125647 1133 125681
rect 1167 125647 1225 125681
rect 1259 125647 1317 125681
rect 1104 125616 1340 125647
rect 1104 125137 1340 125168
rect 1104 125103 1133 125137
rect 1167 125103 1225 125137
rect 1259 125103 1317 125137
rect 1104 125072 1340 125103
rect 1104 124593 1340 124624
rect 1104 124559 1133 124593
rect 1167 124559 1225 124593
rect 1259 124559 1317 124593
rect 1104 124528 1340 124559
rect 1104 124049 1340 124080
rect 1104 124015 1133 124049
rect 1167 124015 1225 124049
rect 1259 124015 1317 124049
rect 1104 123984 1340 124015
rect 1104 123505 1340 123536
rect 1104 123471 1133 123505
rect 1167 123471 1225 123505
rect 1259 123471 1317 123505
rect 1104 123440 1340 123471
rect 1104 122961 1340 122992
rect 1104 122927 1133 122961
rect 1167 122927 1225 122961
rect 1259 122927 1317 122961
rect 1104 122896 1340 122927
rect 1104 122417 1340 122448
rect 1104 122383 1133 122417
rect 1167 122383 1225 122417
rect 1259 122383 1317 122417
rect 1104 122352 1340 122383
rect 1104 121873 1340 121904
rect 1104 121839 1133 121873
rect 1167 121839 1225 121873
rect 1259 121839 1317 121873
rect 1104 121808 1340 121839
rect 1104 121329 1340 121360
rect 1104 121295 1133 121329
rect 1167 121295 1225 121329
rect 1259 121295 1317 121329
rect 1104 121264 1340 121295
rect 1104 120785 1340 120816
rect 1104 120751 1133 120785
rect 1167 120751 1225 120785
rect 1259 120751 1317 120785
rect 1104 120720 1340 120751
rect 1104 120241 1340 120272
rect 1104 120207 1133 120241
rect 1167 120207 1225 120241
rect 1259 120207 1317 120241
rect 1104 120176 1340 120207
rect 1104 119697 1340 119728
rect 1104 119663 1133 119697
rect 1167 119663 1225 119697
rect 1259 119663 1317 119697
rect 1104 119632 1340 119663
rect 1104 119153 1340 119184
rect 1104 119119 1133 119153
rect 1167 119119 1225 119153
rect 1259 119119 1317 119153
rect 1104 119088 1340 119119
rect 1104 118609 1340 118640
rect 1104 118575 1133 118609
rect 1167 118575 1225 118609
rect 1259 118575 1317 118609
rect 1104 118544 1340 118575
rect 1104 118065 1340 118096
rect 1104 118031 1133 118065
rect 1167 118031 1225 118065
rect 1259 118031 1317 118065
rect 1104 118000 1340 118031
rect 1104 117521 1340 117552
rect 1104 117487 1133 117521
rect 1167 117487 1225 117521
rect 1259 117487 1317 117521
rect 1104 117456 1340 117487
rect 1104 116977 1340 117008
rect 1104 116943 1133 116977
rect 1167 116943 1225 116977
rect 1259 116943 1317 116977
rect 1104 116912 1340 116943
rect 1104 116433 1340 116464
rect 1104 116399 1133 116433
rect 1167 116399 1225 116433
rect 1259 116399 1317 116433
rect 1104 116368 1340 116399
rect 1104 115889 1340 115920
rect 1104 115855 1133 115889
rect 1167 115855 1225 115889
rect 1259 115855 1317 115889
rect 1104 115824 1340 115855
rect 1104 115345 1340 115376
rect 1104 115311 1133 115345
rect 1167 115311 1225 115345
rect 1259 115311 1317 115345
rect 1104 115280 1340 115311
rect 1104 114801 1340 114832
rect 1104 114767 1133 114801
rect 1167 114767 1225 114801
rect 1259 114767 1317 114801
rect 1104 114736 1340 114767
rect 1104 114257 1340 114288
rect 1104 114223 1133 114257
rect 1167 114223 1225 114257
rect 1259 114223 1317 114257
rect 1104 114192 1340 114223
rect 1104 113713 1340 113744
rect 1104 113679 1133 113713
rect 1167 113679 1225 113713
rect 1259 113679 1317 113713
rect 1104 113648 1340 113679
rect 1104 113169 1340 113200
rect 1104 113135 1133 113169
rect 1167 113135 1225 113169
rect 1259 113135 1317 113169
rect 1104 113104 1340 113135
rect 1104 112625 1340 112656
rect 1104 112591 1133 112625
rect 1167 112591 1225 112625
rect 1259 112591 1317 112625
rect 1104 112560 1340 112591
rect 1104 112081 1340 112112
rect 1104 112047 1133 112081
rect 1167 112047 1225 112081
rect 1259 112047 1317 112081
rect 1104 112016 1340 112047
rect 1104 111537 1340 111568
rect 1104 111503 1133 111537
rect 1167 111503 1225 111537
rect 1259 111503 1317 111537
rect 1104 111472 1340 111503
rect 1104 110993 1340 111024
rect 1104 110959 1133 110993
rect 1167 110959 1225 110993
rect 1259 110959 1317 110993
rect 1104 110928 1340 110959
rect 1104 110449 1340 110480
rect 1104 110415 1133 110449
rect 1167 110415 1225 110449
rect 1259 110415 1317 110449
rect 1104 110384 1340 110415
rect 1104 109905 1340 109936
rect 1104 109871 1133 109905
rect 1167 109871 1225 109905
rect 1259 109871 1317 109905
rect 1104 109840 1340 109871
rect 1104 109361 1340 109392
rect 1104 109327 1133 109361
rect 1167 109327 1225 109361
rect 1259 109327 1317 109361
rect 1104 109296 1340 109327
rect 1104 108817 1340 108848
rect 1104 108783 1133 108817
rect 1167 108783 1225 108817
rect 1259 108783 1317 108817
rect 1104 108752 1340 108783
rect 1104 108273 1340 108304
rect 1104 108239 1133 108273
rect 1167 108239 1225 108273
rect 1259 108239 1317 108273
rect 1104 108208 1340 108239
rect 1104 107729 1340 107760
rect 1104 107695 1133 107729
rect 1167 107695 1225 107729
rect 1259 107695 1317 107729
rect 1104 107664 1340 107695
rect 1104 107185 1340 107216
rect 1104 107151 1133 107185
rect 1167 107151 1225 107185
rect 1259 107151 1317 107185
rect 1104 107120 1340 107151
rect 1104 106641 1340 106672
rect 1104 106607 1133 106641
rect 1167 106607 1225 106641
rect 1259 106607 1317 106641
rect 1104 106576 1340 106607
rect 1104 106097 1340 106128
rect 1104 106063 1133 106097
rect 1167 106063 1225 106097
rect 1259 106063 1317 106097
rect 1104 106032 1340 106063
rect 1104 105553 1340 105584
rect 1104 105519 1133 105553
rect 1167 105519 1225 105553
rect 1259 105519 1317 105553
rect 1104 105488 1340 105519
rect 1104 105009 1340 105040
rect 1104 104975 1133 105009
rect 1167 104975 1225 105009
rect 1259 104975 1317 105009
rect 1104 104944 1340 104975
rect 1104 104465 1340 104496
rect 1104 104431 1133 104465
rect 1167 104431 1225 104465
rect 1259 104431 1317 104465
rect 1104 104400 1340 104431
rect 1104 103921 1340 103952
rect 1104 103887 1133 103921
rect 1167 103887 1225 103921
rect 1259 103887 1317 103921
rect 1104 103856 1340 103887
rect 1104 103377 1340 103408
rect 1104 103343 1133 103377
rect 1167 103343 1225 103377
rect 1259 103343 1317 103377
rect 1104 103312 1340 103343
rect 1104 102833 1340 102864
rect 1104 102799 1133 102833
rect 1167 102799 1225 102833
rect 1259 102799 1317 102833
rect 1104 102768 1340 102799
rect 1104 102289 1340 102320
rect 1104 102255 1133 102289
rect 1167 102255 1225 102289
rect 1259 102255 1317 102289
rect 1104 102224 1340 102255
rect 1104 101745 1340 101776
rect 1104 101711 1133 101745
rect 1167 101711 1225 101745
rect 1259 101711 1317 101745
rect 1104 101680 1340 101711
rect 1104 101201 1340 101232
rect 1104 101167 1133 101201
rect 1167 101167 1225 101201
rect 1259 101167 1317 101201
rect 1104 101136 1340 101167
rect 1104 100657 1340 100688
rect 1104 100623 1133 100657
rect 1167 100623 1225 100657
rect 1259 100623 1317 100657
rect 1104 100592 1340 100623
rect 1104 100113 1340 100144
rect 1104 100079 1133 100113
rect 1167 100079 1225 100113
rect 1259 100079 1317 100113
rect 1104 100048 1340 100079
rect 1104 99569 1340 99600
rect 1104 99535 1133 99569
rect 1167 99535 1225 99569
rect 1259 99535 1317 99569
rect 1104 99504 1340 99535
rect 1104 99025 1340 99056
rect 1104 98991 1133 99025
rect 1167 98991 1225 99025
rect 1259 98991 1317 99025
rect 1104 98960 1340 98991
rect 1104 98481 1340 98512
rect 1104 98447 1133 98481
rect 1167 98447 1225 98481
rect 1259 98447 1317 98481
rect 1104 98416 1340 98447
rect 1104 97937 1340 97968
rect 1104 97903 1133 97937
rect 1167 97903 1225 97937
rect 1259 97903 1317 97937
rect 1104 97872 1340 97903
rect 1104 97393 1340 97424
rect 1104 97359 1133 97393
rect 1167 97359 1225 97393
rect 1259 97359 1317 97393
rect 1104 97328 1340 97359
rect 1104 96849 1340 96880
rect 1104 96815 1133 96849
rect 1167 96815 1225 96849
rect 1259 96815 1317 96849
rect 1104 96784 1340 96815
rect 1104 96305 1340 96336
rect 1104 96271 1133 96305
rect 1167 96271 1225 96305
rect 1259 96271 1317 96305
rect 1104 96240 1340 96271
rect 1104 95761 1340 95792
rect 1104 95727 1133 95761
rect 1167 95727 1225 95761
rect 1259 95727 1317 95761
rect 1104 95696 1340 95727
rect 1104 95217 1340 95248
rect 1104 95183 1133 95217
rect 1167 95183 1225 95217
rect 1259 95183 1317 95217
rect 1104 95152 1340 95183
rect 1104 94673 1340 94704
rect 1104 94639 1133 94673
rect 1167 94639 1225 94673
rect 1259 94639 1317 94673
rect 1104 94608 1340 94639
rect 1104 94129 1340 94160
rect 1104 94095 1133 94129
rect 1167 94095 1225 94129
rect 1259 94095 1317 94129
rect 1104 94064 1340 94095
rect 1104 93585 1340 93616
rect 1104 93551 1133 93585
rect 1167 93551 1225 93585
rect 1259 93551 1317 93585
rect 1104 93520 1340 93551
rect 1104 93041 1340 93072
rect 1104 93007 1133 93041
rect 1167 93007 1225 93041
rect 1259 93007 1317 93041
rect 1104 92976 1340 93007
rect 1104 92497 1340 92528
rect 1104 92463 1133 92497
rect 1167 92463 1225 92497
rect 1259 92463 1317 92497
rect 1104 92432 1340 92463
rect 1104 91953 1340 91984
rect 1104 91919 1133 91953
rect 1167 91919 1225 91953
rect 1259 91919 1317 91953
rect 1104 91888 1340 91919
rect 1104 91409 1340 91440
rect 1104 91375 1133 91409
rect 1167 91375 1225 91409
rect 1259 91375 1317 91409
rect 1104 91344 1340 91375
rect 1104 90865 1340 90896
rect 1104 90831 1133 90865
rect 1167 90831 1225 90865
rect 1259 90831 1317 90865
rect 1104 90800 1340 90831
rect 1104 90321 1340 90352
rect 1104 90287 1133 90321
rect 1167 90287 1225 90321
rect 1259 90287 1317 90321
rect 1104 90256 1340 90287
rect 1104 89777 1340 89808
rect 1104 89743 1133 89777
rect 1167 89743 1225 89777
rect 1259 89743 1317 89777
rect 1104 89712 1340 89743
rect 1104 89233 1340 89264
rect 1104 89199 1133 89233
rect 1167 89199 1225 89233
rect 1259 89199 1317 89233
rect 1104 89168 1340 89199
rect 1104 88689 1340 88720
rect 1104 88655 1133 88689
rect 1167 88655 1225 88689
rect 1259 88655 1317 88689
rect 1104 88624 1340 88655
rect 1104 88145 1340 88176
rect 1104 88111 1133 88145
rect 1167 88111 1225 88145
rect 1259 88111 1317 88145
rect 1104 88080 1340 88111
rect 1104 87601 1340 87632
rect 1104 87567 1133 87601
rect 1167 87567 1225 87601
rect 1259 87567 1317 87601
rect 1104 87536 1340 87567
rect 1104 87057 1340 87088
rect 1104 87023 1133 87057
rect 1167 87023 1225 87057
rect 1259 87023 1317 87057
rect 1104 86992 1340 87023
rect 1104 86513 1340 86544
rect 1104 86479 1133 86513
rect 1167 86479 1225 86513
rect 1259 86479 1317 86513
rect 1104 86448 1340 86479
rect 1104 85969 1340 86000
rect 1104 85935 1133 85969
rect 1167 85935 1225 85969
rect 1259 85935 1317 85969
rect 1104 85904 1340 85935
rect 1104 85425 1340 85456
rect 1104 85391 1133 85425
rect 1167 85391 1225 85425
rect 1259 85391 1317 85425
rect 1104 85360 1340 85391
rect 1104 84881 1340 84912
rect 1104 84847 1133 84881
rect 1167 84847 1225 84881
rect 1259 84847 1317 84881
rect 1104 84816 1340 84847
rect 1104 84337 1340 84368
rect 1104 84303 1133 84337
rect 1167 84303 1225 84337
rect 1259 84303 1317 84337
rect 1104 84272 1340 84303
rect 1104 83793 1340 83824
rect 1104 83759 1133 83793
rect 1167 83759 1225 83793
rect 1259 83759 1317 83793
rect 1104 83728 1340 83759
rect 1104 83249 1340 83280
rect 1104 83215 1133 83249
rect 1167 83215 1225 83249
rect 1259 83215 1317 83249
rect 1104 83184 1340 83215
rect 1104 82705 1340 82736
rect 1104 82671 1133 82705
rect 1167 82671 1225 82705
rect 1259 82671 1317 82705
rect 1104 82640 1340 82671
rect 1104 82161 1340 82192
rect 1104 82127 1133 82161
rect 1167 82127 1225 82161
rect 1259 82127 1317 82161
rect 1104 82096 1340 82127
rect 1104 81617 1340 81648
rect 1104 81583 1133 81617
rect 1167 81583 1225 81617
rect 1259 81583 1317 81617
rect 1104 81552 1340 81583
rect 1104 81073 1340 81104
rect 1104 81039 1133 81073
rect 1167 81039 1225 81073
rect 1259 81039 1317 81073
rect 1104 81008 1340 81039
rect 1104 80529 1340 80560
rect 1104 80495 1133 80529
rect 1167 80495 1225 80529
rect 1259 80495 1317 80529
rect 1104 80464 1340 80495
rect 1104 79985 1340 80016
rect 1104 79951 1133 79985
rect 1167 79951 1225 79985
rect 1259 79951 1317 79985
rect 1104 79920 1340 79951
rect 1104 79441 1340 79472
rect 1104 79407 1133 79441
rect 1167 79407 1225 79441
rect 1259 79407 1317 79441
rect 1104 79376 1340 79407
rect 1104 78897 1340 78928
rect 1104 78863 1133 78897
rect 1167 78863 1225 78897
rect 1259 78863 1317 78897
rect 1104 78832 1340 78863
rect 1104 78353 1340 78384
rect 1104 78319 1133 78353
rect 1167 78319 1225 78353
rect 1259 78319 1317 78353
rect 1104 78288 1340 78319
rect 1104 77809 1340 77840
rect 1104 77775 1133 77809
rect 1167 77775 1225 77809
rect 1259 77775 1317 77809
rect 1104 77744 1340 77775
rect 1104 77265 1340 77296
rect 1104 77231 1133 77265
rect 1167 77231 1225 77265
rect 1259 77231 1317 77265
rect 1104 77200 1340 77231
rect 1104 76721 1340 76752
rect 1104 76687 1133 76721
rect 1167 76687 1225 76721
rect 1259 76687 1317 76721
rect 1104 76656 1340 76687
rect 1104 76177 1340 76208
rect 1104 76143 1133 76177
rect 1167 76143 1225 76177
rect 1259 76143 1317 76177
rect 1104 76112 1340 76143
rect 1104 75633 1340 75664
rect 1104 75599 1133 75633
rect 1167 75599 1225 75633
rect 1259 75599 1317 75633
rect 1104 75568 1340 75599
rect 1104 75089 1340 75120
rect 1104 75055 1133 75089
rect 1167 75055 1225 75089
rect 1259 75055 1317 75089
rect 1104 75024 1340 75055
rect 1104 74545 1340 74576
rect 1104 74511 1133 74545
rect 1167 74511 1225 74545
rect 1259 74511 1317 74545
rect 1104 74480 1340 74511
rect 1104 74001 1340 74032
rect 1104 73967 1133 74001
rect 1167 73967 1225 74001
rect 1259 73967 1317 74001
rect 1104 73936 1340 73967
rect 1104 73457 1340 73488
rect 1104 73423 1133 73457
rect 1167 73423 1225 73457
rect 1259 73423 1317 73457
rect 1104 73392 1340 73423
rect 1104 72913 1340 72944
rect 1104 72879 1133 72913
rect 1167 72879 1225 72913
rect 1259 72879 1317 72913
rect 1104 72848 1340 72879
rect 1104 72369 1340 72400
rect 1104 72335 1133 72369
rect 1167 72335 1225 72369
rect 1259 72335 1317 72369
rect 1104 72304 1340 72335
rect 1104 71825 1340 71856
rect 1104 71791 1133 71825
rect 1167 71791 1225 71825
rect 1259 71791 1317 71825
rect 1104 71760 1340 71791
rect 1104 71281 1340 71312
rect 1104 71247 1133 71281
rect 1167 71247 1225 71281
rect 1259 71247 1317 71281
rect 1104 71216 1340 71247
rect 1104 70737 1340 70768
rect 1104 70703 1133 70737
rect 1167 70703 1225 70737
rect 1259 70703 1317 70737
rect 1104 70672 1340 70703
rect 1104 70193 1340 70224
rect 1104 70159 1133 70193
rect 1167 70159 1225 70193
rect 1259 70159 1317 70193
rect 1104 70128 1340 70159
rect 1104 69649 1340 69680
rect 1104 69615 1133 69649
rect 1167 69615 1225 69649
rect 1259 69615 1317 69649
rect 1104 69584 1340 69615
rect 1104 69105 1340 69136
rect 1104 69071 1133 69105
rect 1167 69071 1225 69105
rect 1259 69071 1317 69105
rect 1104 69040 1340 69071
rect 1104 68561 1340 68592
rect 1104 68527 1133 68561
rect 1167 68527 1225 68561
rect 1259 68527 1317 68561
rect 1104 68496 1340 68527
rect 1104 68017 1340 68048
rect 1104 67983 1133 68017
rect 1167 67983 1225 68017
rect 1259 67983 1317 68017
rect 1104 67952 1340 67983
rect 1104 67473 1340 67504
rect 1104 67439 1133 67473
rect 1167 67439 1225 67473
rect 1259 67439 1317 67473
rect 1104 67408 1340 67439
rect 1104 66929 1340 66960
rect 1104 66895 1133 66929
rect 1167 66895 1225 66929
rect 1259 66895 1317 66929
rect 1104 66864 1340 66895
rect 1104 66385 1340 66416
rect 1104 66351 1133 66385
rect 1167 66351 1225 66385
rect 1259 66351 1317 66385
rect 1104 66320 1340 66351
rect 1104 65841 1340 65872
rect 1104 65807 1133 65841
rect 1167 65807 1225 65841
rect 1259 65807 1317 65841
rect 1104 65776 1340 65807
rect 1104 65297 1340 65328
rect 1104 65263 1133 65297
rect 1167 65263 1225 65297
rect 1259 65263 1317 65297
rect 1104 65232 1340 65263
rect 1104 64753 1340 64784
rect 1104 64719 1133 64753
rect 1167 64719 1225 64753
rect 1259 64719 1317 64753
rect 1104 64688 1340 64719
rect 1104 64209 1340 64240
rect 1104 64175 1133 64209
rect 1167 64175 1225 64209
rect 1259 64175 1317 64209
rect 1104 64144 1340 64175
rect 1104 63665 1340 63696
rect 1104 63631 1133 63665
rect 1167 63631 1225 63665
rect 1259 63631 1317 63665
rect 1104 63600 1340 63631
rect 1104 63121 1340 63152
rect 1104 63087 1133 63121
rect 1167 63087 1225 63121
rect 1259 63087 1317 63121
rect 1104 63056 1340 63087
rect 1104 62577 1340 62608
rect 1104 62543 1133 62577
rect 1167 62543 1225 62577
rect 1259 62543 1317 62577
rect 1104 62512 1340 62543
rect 1104 62033 1340 62064
rect 1104 61999 1133 62033
rect 1167 61999 1225 62033
rect 1259 61999 1317 62033
rect 1104 61968 1340 61999
rect 1104 61489 1340 61520
rect 1104 61455 1133 61489
rect 1167 61455 1225 61489
rect 1259 61455 1317 61489
rect 1104 61424 1340 61455
rect 1104 60945 1340 60976
rect 1104 60911 1133 60945
rect 1167 60911 1225 60945
rect 1259 60911 1317 60945
rect 1104 60880 1340 60911
rect 1104 60401 1340 60432
rect 1104 60367 1133 60401
rect 1167 60367 1225 60401
rect 1259 60367 1317 60401
rect 1104 60336 1340 60367
rect 1104 59857 1340 59888
rect 1104 59823 1133 59857
rect 1167 59823 1225 59857
rect 1259 59823 1317 59857
rect 1104 59792 1340 59823
rect 1104 59313 1340 59344
rect 1104 59279 1133 59313
rect 1167 59279 1225 59313
rect 1259 59279 1317 59313
rect 1104 59248 1340 59279
rect 1104 58769 1340 58800
rect 1104 58735 1133 58769
rect 1167 58735 1225 58769
rect 1259 58735 1317 58769
rect 1104 58704 1340 58735
rect 1104 58225 1340 58256
rect 1104 58191 1133 58225
rect 1167 58191 1225 58225
rect 1259 58191 1317 58225
rect 1104 58160 1340 58191
rect 1104 57681 1340 57712
rect 1104 57647 1133 57681
rect 1167 57647 1225 57681
rect 1259 57647 1317 57681
rect 1104 57616 1340 57647
rect 1104 57137 1340 57168
rect 1104 57103 1133 57137
rect 1167 57103 1225 57137
rect 1259 57103 1317 57137
rect 1104 57072 1340 57103
rect 1104 56593 1340 56624
rect 1104 56559 1133 56593
rect 1167 56559 1225 56593
rect 1259 56559 1317 56593
rect 1104 56528 1340 56559
rect 1104 56049 1340 56080
rect 1104 56015 1133 56049
rect 1167 56015 1225 56049
rect 1259 56015 1317 56049
rect 1104 55984 1340 56015
rect 1104 55505 1340 55536
rect 1104 55471 1133 55505
rect 1167 55471 1225 55505
rect 1259 55471 1317 55505
rect 1104 55440 1340 55471
rect 1104 54961 1340 54992
rect 1104 54927 1133 54961
rect 1167 54927 1225 54961
rect 1259 54927 1317 54961
rect 1104 54896 1340 54927
rect 1104 54417 1340 54448
rect 1104 54383 1133 54417
rect 1167 54383 1225 54417
rect 1259 54383 1317 54417
rect 1104 54352 1340 54383
rect 1104 53873 1340 53904
rect 1104 53839 1133 53873
rect 1167 53839 1225 53873
rect 1259 53839 1317 53873
rect 1104 53808 1340 53839
rect 1104 53329 1340 53360
rect 1104 53295 1133 53329
rect 1167 53295 1225 53329
rect 1259 53295 1317 53329
rect 1104 53264 1340 53295
rect 1104 52785 1340 52816
rect 1104 52751 1133 52785
rect 1167 52751 1225 52785
rect 1259 52751 1317 52785
rect 1104 52720 1340 52751
rect 1104 52241 1340 52272
rect 1104 52207 1133 52241
rect 1167 52207 1225 52241
rect 1259 52207 1317 52241
rect 1104 52176 1340 52207
rect 1104 51697 1340 51728
rect 1104 51663 1133 51697
rect 1167 51663 1225 51697
rect 1259 51663 1317 51697
rect 1104 51632 1340 51663
rect 1104 51153 1340 51184
rect 1104 51119 1133 51153
rect 1167 51119 1225 51153
rect 1259 51119 1317 51153
rect 1104 51088 1340 51119
rect 1104 50609 1340 50640
rect 1104 50575 1133 50609
rect 1167 50575 1225 50609
rect 1259 50575 1317 50609
rect 1104 50544 1340 50575
rect 1104 50065 1340 50096
rect 1104 50031 1133 50065
rect 1167 50031 1225 50065
rect 1259 50031 1317 50065
rect 1104 50000 1340 50031
rect 1104 49521 1340 49552
rect 1104 49487 1133 49521
rect 1167 49487 1225 49521
rect 1259 49487 1317 49521
rect 1104 49456 1340 49487
rect 1104 48977 1340 49008
rect 1104 48943 1133 48977
rect 1167 48943 1225 48977
rect 1259 48943 1317 48977
rect 1104 48912 1340 48943
rect 1104 48433 1340 48464
rect 1104 48399 1133 48433
rect 1167 48399 1225 48433
rect 1259 48399 1317 48433
rect 1104 48368 1340 48399
rect 1104 47889 1340 47920
rect 1104 47855 1133 47889
rect 1167 47855 1225 47889
rect 1259 47855 1317 47889
rect 1104 47824 1340 47855
rect 1104 47345 1340 47376
rect 1104 47311 1133 47345
rect 1167 47311 1225 47345
rect 1259 47311 1317 47345
rect 1104 47280 1340 47311
rect 1104 46801 1340 46832
rect 1104 46767 1133 46801
rect 1167 46767 1225 46801
rect 1259 46767 1317 46801
rect 1104 46736 1340 46767
rect 1104 46257 1340 46288
rect 1104 46223 1133 46257
rect 1167 46223 1225 46257
rect 1259 46223 1317 46257
rect 1104 46192 1340 46223
rect 1104 45713 1340 45744
rect 1104 45679 1133 45713
rect 1167 45679 1225 45713
rect 1259 45679 1317 45713
rect 1104 45648 1340 45679
rect 1104 45169 1340 45200
rect 1104 45135 1133 45169
rect 1167 45135 1225 45169
rect 1259 45135 1317 45169
rect 1104 45104 1340 45135
rect 1104 44625 1340 44656
rect 1104 44591 1133 44625
rect 1167 44591 1225 44625
rect 1259 44591 1317 44625
rect 1104 44560 1340 44591
rect 1104 44081 1340 44112
rect 1104 44047 1133 44081
rect 1167 44047 1225 44081
rect 1259 44047 1317 44081
rect 1104 44016 1340 44047
rect 1104 43537 1340 43568
rect 1104 43503 1133 43537
rect 1167 43503 1225 43537
rect 1259 43503 1317 43537
rect 1104 43472 1340 43503
rect 1104 42993 1340 43024
rect 1104 42959 1133 42993
rect 1167 42959 1225 42993
rect 1259 42959 1317 42993
rect 1104 42928 1340 42959
rect 1104 42449 1340 42480
rect 1104 42415 1133 42449
rect 1167 42415 1225 42449
rect 1259 42415 1317 42449
rect 1104 42384 1340 42415
rect 1104 41905 1340 41936
rect 1104 41871 1133 41905
rect 1167 41871 1225 41905
rect 1259 41871 1317 41905
rect 1104 41840 1340 41871
rect 1104 41361 1340 41392
rect 1104 41327 1133 41361
rect 1167 41327 1225 41361
rect 1259 41327 1317 41361
rect 1104 41296 1340 41327
rect 1104 40817 1340 40848
rect 1104 40783 1133 40817
rect 1167 40783 1225 40817
rect 1259 40783 1317 40817
rect 1104 40752 1340 40783
rect 1104 40273 1340 40304
rect 1104 40239 1133 40273
rect 1167 40239 1225 40273
rect 1259 40239 1317 40273
rect 1104 40208 1340 40239
rect 1104 39729 1340 39760
rect 1104 39695 1133 39729
rect 1167 39695 1225 39729
rect 1259 39695 1317 39729
rect 1104 39664 1340 39695
rect 1104 39185 1340 39216
rect 1104 39151 1133 39185
rect 1167 39151 1225 39185
rect 1259 39151 1317 39185
rect 1104 39120 1340 39151
rect 1104 38641 1340 38672
rect 1104 38607 1133 38641
rect 1167 38607 1225 38641
rect 1259 38607 1317 38641
rect 1104 38576 1340 38607
rect 1104 38097 1340 38128
rect 1104 38063 1133 38097
rect 1167 38063 1225 38097
rect 1259 38063 1317 38097
rect 1104 38032 1340 38063
rect 1104 37553 1340 37584
rect 1104 37519 1133 37553
rect 1167 37519 1225 37553
rect 1259 37519 1317 37553
rect 1104 37488 1340 37519
rect 1104 37009 1340 37040
rect 1104 36975 1133 37009
rect 1167 36975 1225 37009
rect 1259 36975 1317 37009
rect 1104 36944 1340 36975
rect 1104 36465 1340 36496
rect 1104 36431 1133 36465
rect 1167 36431 1225 36465
rect 1259 36431 1317 36465
rect 1104 36400 1340 36431
rect 1104 35921 1340 35952
rect 1104 35887 1133 35921
rect 1167 35887 1225 35921
rect 1259 35887 1317 35921
rect 1104 35856 1340 35887
rect 1104 35377 1340 35408
rect 1104 35343 1133 35377
rect 1167 35343 1225 35377
rect 1259 35343 1317 35377
rect 1104 35312 1340 35343
rect 1104 34833 1340 34864
rect 1104 34799 1133 34833
rect 1167 34799 1225 34833
rect 1259 34799 1317 34833
rect 1104 34768 1340 34799
rect 1104 34289 1340 34320
rect 1104 34255 1133 34289
rect 1167 34255 1225 34289
rect 1259 34255 1317 34289
rect 1104 34224 1340 34255
rect 1104 33745 1340 33776
rect 1104 33711 1133 33745
rect 1167 33711 1225 33745
rect 1259 33711 1317 33745
rect 1104 33680 1340 33711
rect 1104 33201 1340 33232
rect 1104 33167 1133 33201
rect 1167 33167 1225 33201
rect 1259 33167 1317 33201
rect 1104 33136 1340 33167
rect 1104 32657 1340 32688
rect 1104 32623 1133 32657
rect 1167 32623 1225 32657
rect 1259 32623 1317 32657
rect 1104 32592 1340 32623
rect 1104 32113 1340 32144
rect 1104 32079 1133 32113
rect 1167 32079 1225 32113
rect 1259 32079 1317 32113
rect 1104 32048 1340 32079
rect 1104 31569 1340 31600
rect 1104 31535 1133 31569
rect 1167 31535 1225 31569
rect 1259 31535 1317 31569
rect 1104 31504 1340 31535
rect 1104 31025 1340 31056
rect 1104 30991 1133 31025
rect 1167 30991 1225 31025
rect 1259 30991 1317 31025
rect 1104 30960 1340 30991
rect 1104 30481 1340 30512
rect 1104 30447 1133 30481
rect 1167 30447 1225 30481
rect 1259 30447 1317 30481
rect 1104 30416 1340 30447
rect 1104 29937 1340 29968
rect 1104 29903 1133 29937
rect 1167 29903 1225 29937
rect 1259 29903 1317 29937
rect 1104 29872 1340 29903
rect 1104 29393 1340 29424
rect 1104 29359 1133 29393
rect 1167 29359 1225 29393
rect 1259 29359 1317 29393
rect 1104 29328 1340 29359
rect 1104 28849 1340 28880
rect 1104 28815 1133 28849
rect 1167 28815 1225 28849
rect 1259 28815 1317 28849
rect 1104 28784 1340 28815
rect 1104 28305 1340 28336
rect 1104 28271 1133 28305
rect 1167 28271 1225 28305
rect 1259 28271 1317 28305
rect 1104 28240 1340 28271
rect 1104 27761 1340 27792
rect 1104 27727 1133 27761
rect 1167 27727 1225 27761
rect 1259 27727 1317 27761
rect 1104 27696 1340 27727
rect 1104 27217 1340 27248
rect 1104 27183 1133 27217
rect 1167 27183 1225 27217
rect 1259 27183 1317 27217
rect 1104 27152 1340 27183
rect 1104 26673 1340 26704
rect 1104 26639 1133 26673
rect 1167 26639 1225 26673
rect 1259 26639 1317 26673
rect 1104 26608 1340 26639
rect 1104 26129 1340 26160
rect 1104 26095 1133 26129
rect 1167 26095 1225 26129
rect 1259 26095 1317 26129
rect 1104 26064 1340 26095
rect 1104 25585 1340 25616
rect 1104 25551 1133 25585
rect 1167 25551 1225 25585
rect 1259 25551 1317 25585
rect 1104 25520 1340 25551
rect 1104 25041 1340 25072
rect 1104 25007 1133 25041
rect 1167 25007 1225 25041
rect 1259 25007 1317 25041
rect 1104 24976 1340 25007
rect 1104 24497 1340 24528
rect 1104 24463 1133 24497
rect 1167 24463 1225 24497
rect 1259 24463 1317 24497
rect 1104 24432 1340 24463
rect 1104 23953 1340 23984
rect 1104 23919 1133 23953
rect 1167 23919 1225 23953
rect 1259 23919 1317 23953
rect 1104 23888 1340 23919
rect 1104 23409 1340 23440
rect 1104 23375 1133 23409
rect 1167 23375 1225 23409
rect 1259 23375 1317 23409
rect 1104 23344 1340 23375
rect 1104 22865 1340 22896
rect 1104 22831 1133 22865
rect 1167 22831 1225 22865
rect 1259 22831 1317 22865
rect 1104 22800 1340 22831
rect 1104 22321 1340 22352
rect 1104 22287 1133 22321
rect 1167 22287 1225 22321
rect 1259 22287 1317 22321
rect 1104 22256 1340 22287
rect 1104 21777 1340 21808
rect 1104 21743 1133 21777
rect 1167 21743 1225 21777
rect 1259 21743 1317 21777
rect 1104 21712 1340 21743
rect 1104 21233 1340 21264
rect 1104 21199 1133 21233
rect 1167 21199 1225 21233
rect 1259 21199 1317 21233
rect 1104 21168 1340 21199
rect 1104 20689 1340 20720
rect 1104 20655 1133 20689
rect 1167 20655 1225 20689
rect 1259 20655 1317 20689
rect 1104 20624 1340 20655
rect 1104 20145 1340 20176
rect 1104 20111 1133 20145
rect 1167 20111 1225 20145
rect 1259 20111 1317 20145
rect 1104 20080 1340 20111
rect 1104 19601 1340 19632
rect 1104 19567 1133 19601
rect 1167 19567 1225 19601
rect 1259 19567 1317 19601
rect 1104 19536 1340 19567
rect 1104 19057 1340 19088
rect 1104 19023 1133 19057
rect 1167 19023 1225 19057
rect 1259 19023 1317 19057
rect 1104 18992 1340 19023
rect 1104 18513 1340 18544
rect 1104 18479 1133 18513
rect 1167 18479 1225 18513
rect 1259 18479 1317 18513
rect 1104 18448 1340 18479
rect 1104 17969 1340 18000
rect 1104 17935 1133 17969
rect 1167 17935 1225 17969
rect 1259 17935 1317 17969
rect 1104 17904 1340 17935
rect 1104 17425 1340 17456
rect 1104 17391 1133 17425
rect 1167 17391 1225 17425
rect 1259 17391 1317 17425
rect 1104 17360 1340 17391
rect 1104 16881 1340 16912
rect 1104 16847 1133 16881
rect 1167 16847 1225 16881
rect 1259 16847 1317 16881
rect 1104 16816 1340 16847
rect 1104 16337 1340 16368
rect 1104 16303 1133 16337
rect 1167 16303 1225 16337
rect 1259 16303 1317 16337
rect 1104 16272 1340 16303
rect 1104 15793 1340 15824
rect 1104 15759 1133 15793
rect 1167 15759 1225 15793
rect 1259 15759 1317 15793
rect 1104 15728 1340 15759
rect 1104 15249 1340 15280
rect 1104 15215 1133 15249
rect 1167 15215 1225 15249
rect 1259 15215 1317 15249
rect 1104 15184 1340 15215
rect 1104 14705 1340 14736
rect 1104 14671 1133 14705
rect 1167 14671 1225 14705
rect 1259 14671 1317 14705
rect 1104 14640 1340 14671
rect 1104 14161 1340 14192
rect 1104 14127 1133 14161
rect 1167 14127 1225 14161
rect 1259 14127 1317 14161
rect 1104 14096 1340 14127
rect 1104 13617 1340 13648
rect 1104 13583 1133 13617
rect 1167 13583 1225 13617
rect 1259 13583 1317 13617
rect 1104 13552 1340 13583
rect 1104 13073 1340 13104
rect 1104 13039 1133 13073
rect 1167 13039 1225 13073
rect 1259 13039 1317 13073
rect 1104 13008 1340 13039
rect 1104 12529 1340 12560
rect 1104 12495 1133 12529
rect 1167 12495 1225 12529
rect 1259 12495 1317 12529
rect 1104 12464 1340 12495
rect 1104 11985 1340 12016
rect 1104 11951 1133 11985
rect 1167 11951 1225 11985
rect 1259 11951 1317 11985
rect 1104 11920 1340 11951
rect 1104 11441 1340 11472
rect 1104 11407 1133 11441
rect 1167 11407 1225 11441
rect 1259 11407 1317 11441
rect 1104 11376 1340 11407
rect 1104 10897 1340 10928
rect 1104 10863 1133 10897
rect 1167 10863 1225 10897
rect 1259 10863 1317 10897
rect 1104 10832 1340 10863
rect 1104 10353 1340 10384
rect 1104 10319 1133 10353
rect 1167 10319 1225 10353
rect 1259 10319 1317 10353
rect 1104 10288 1340 10319
rect 1104 9809 1340 9840
rect 1104 9775 1133 9809
rect 1167 9775 1225 9809
rect 1259 9775 1317 9809
rect 1104 9744 1340 9775
rect 1104 9265 1340 9296
rect 1104 9231 1133 9265
rect 1167 9231 1225 9265
rect 1259 9231 1317 9265
rect 1104 9200 1340 9231
rect 1104 8721 1340 8752
rect 1104 8687 1133 8721
rect 1167 8687 1225 8721
rect 1259 8687 1317 8721
rect 1104 8656 1340 8687
rect 1104 8177 1340 8208
rect 1104 8143 1133 8177
rect 1167 8143 1225 8177
rect 1259 8143 1317 8177
rect 1104 8112 1340 8143
rect 1104 7633 1340 7664
rect 1104 7599 1133 7633
rect 1167 7599 1225 7633
rect 1259 7599 1317 7633
rect 1104 7568 1340 7599
rect 1104 7089 1340 7120
rect 1104 7055 1133 7089
rect 1167 7055 1225 7089
rect 1259 7055 1317 7089
rect 1104 7024 1340 7055
rect 1104 6545 1340 6576
rect 1104 6511 1133 6545
rect 1167 6511 1225 6545
rect 1259 6511 1317 6545
rect 1104 6480 1340 6511
rect 1104 6001 1340 6032
rect 1104 5967 1133 6001
rect 1167 5967 1225 6001
rect 1259 5967 1317 6001
rect 1104 5936 1340 5967
rect 1104 5457 1340 5488
rect 1104 5423 1133 5457
rect 1167 5423 1225 5457
rect 1259 5423 1317 5457
rect 1104 5392 1340 5423
rect 1104 4913 1340 4944
rect 1104 4879 1133 4913
rect 1167 4879 1225 4913
rect 1259 4879 1317 4913
rect 1104 4848 1340 4879
rect 1104 4369 1340 4400
rect 1104 4335 1133 4369
rect 1167 4335 1225 4369
rect 1259 4335 1317 4369
rect 1104 4304 1340 4335
rect 290 4088 296 4140
rect 348 4128 354 4140
rect 348 4100 1340 4128
rect 348 4088 354 4100
rect 1104 3825 1340 3856
rect 1104 3791 1133 3825
rect 1167 3791 1225 3825
rect 1259 3791 1317 3825
rect 1104 3760 1340 3791
rect 842 3408 848 3460
rect 900 3448 906 3460
rect 900 3420 1340 3448
rect 900 3408 906 3420
rect 1104 3281 1340 3312
rect 1104 3247 1133 3281
rect 1167 3247 1225 3281
rect 1259 3247 1317 3281
rect 1104 3216 1340 3247
rect 1104 2737 1340 2768
rect 1104 2703 1133 2737
rect 1167 2703 1225 2737
rect 1259 2703 1317 2737
rect 1104 2672 1340 2703
rect 1104 2193 1340 2224
rect 1104 2159 1133 2193
rect 1167 2159 1225 2193
rect 1259 2159 1317 2193
rect 1104 2128 1340 2159
rect 298660 297585 298816 297616
rect 298660 297551 298661 297585
rect 298695 297551 298753 297585
rect 298787 297551 298816 297585
rect 298660 297520 298816 297551
rect 298660 297041 298816 297072
rect 298660 297007 298661 297041
rect 298695 297007 298753 297041
rect 298787 297007 298816 297041
rect 298660 296976 298816 297007
rect 298660 296497 298816 296528
rect 298660 296463 298661 296497
rect 298695 296463 298753 296497
rect 298787 296463 298816 296497
rect 298660 296432 298816 296463
rect 298660 295953 298816 295984
rect 298660 295919 298661 295953
rect 298695 295919 298753 295953
rect 298787 295919 298816 295953
rect 298660 295888 298816 295919
rect 298660 295409 298816 295440
rect 298660 295375 298661 295409
rect 298695 295375 298753 295409
rect 298787 295375 298816 295409
rect 298660 295344 298816 295375
rect 298660 294865 298816 294896
rect 298660 294831 298661 294865
rect 298695 294831 298753 294865
rect 298787 294831 298816 294865
rect 298660 294800 298816 294831
rect 298660 294321 298816 294352
rect 298660 294287 298661 294321
rect 298695 294287 298753 294321
rect 298787 294287 298816 294321
rect 298660 294256 298816 294287
rect 298660 293777 298816 293808
rect 298660 293743 298661 293777
rect 298695 293743 298753 293777
rect 298787 293743 298816 293777
rect 298660 293712 298816 293743
rect 298660 293233 298816 293264
rect 298660 293199 298661 293233
rect 298695 293199 298753 293233
rect 298787 293199 298816 293233
rect 298660 293168 298816 293199
rect 298660 292689 298816 292720
rect 298660 292655 298661 292689
rect 298695 292655 298753 292689
rect 298787 292655 298816 292689
rect 298660 292624 298816 292655
rect 298660 292145 298816 292176
rect 298660 292111 298661 292145
rect 298695 292111 298753 292145
rect 298787 292111 298816 292145
rect 298660 292080 298816 292111
rect 298660 291601 298816 291632
rect 298660 291567 298661 291601
rect 298695 291567 298753 291601
rect 298787 291567 298816 291601
rect 298660 291536 298816 291567
rect 298660 291057 298816 291088
rect 298660 291023 298661 291057
rect 298695 291023 298753 291057
rect 298787 291023 298816 291057
rect 298660 290992 298816 291023
rect 298660 290513 298816 290544
rect 298660 290479 298661 290513
rect 298695 290479 298753 290513
rect 298787 290479 298816 290513
rect 298660 290448 298816 290479
rect 298660 289969 298816 290000
rect 298660 289935 298661 289969
rect 298695 289935 298753 289969
rect 298787 289935 298816 289969
rect 298660 289904 298816 289935
rect 298660 289425 298816 289456
rect 298660 289391 298661 289425
rect 298695 289391 298753 289425
rect 298787 289391 298816 289425
rect 298660 289360 298816 289391
rect 298660 288881 298816 288912
rect 298660 288847 298661 288881
rect 298695 288847 298753 288881
rect 298787 288847 298816 288881
rect 298660 288816 298816 288847
rect 298660 288337 298816 288368
rect 298660 288303 298661 288337
rect 298695 288303 298753 288337
rect 298787 288303 298816 288337
rect 298660 288272 298816 288303
rect 298660 287793 298816 287824
rect 298660 287759 298661 287793
rect 298695 287759 298753 287793
rect 298787 287759 298816 287793
rect 298660 287728 298816 287759
rect 298660 287249 298816 287280
rect 298660 287215 298661 287249
rect 298695 287215 298753 287249
rect 298787 287215 298816 287249
rect 298660 287184 298816 287215
rect 298660 286705 298816 286736
rect 298660 286671 298661 286705
rect 298695 286671 298753 286705
rect 298787 286671 298816 286705
rect 298660 286640 298816 286671
rect 298660 286161 298816 286192
rect 298660 286127 298661 286161
rect 298695 286127 298753 286161
rect 298787 286127 298816 286161
rect 298660 286096 298816 286127
rect 298660 285617 298816 285648
rect 298660 285583 298661 285617
rect 298695 285583 298753 285617
rect 298787 285583 298816 285617
rect 298660 285552 298816 285583
rect 298660 285073 298816 285104
rect 298660 285039 298661 285073
rect 298695 285039 298753 285073
rect 298787 285039 298816 285073
rect 298660 285008 298816 285039
rect 298660 284529 298816 284560
rect 298660 284495 298661 284529
rect 298695 284495 298753 284529
rect 298787 284495 298816 284529
rect 298660 284464 298816 284495
rect 298660 283985 298816 284016
rect 298660 283951 298661 283985
rect 298695 283951 298753 283985
rect 298787 283951 298816 283985
rect 298660 283920 298816 283951
rect 298660 283441 298816 283472
rect 298660 283407 298661 283441
rect 298695 283407 298753 283441
rect 298787 283407 298816 283441
rect 298660 283376 298816 283407
rect 298660 282897 298816 282928
rect 298660 282863 298661 282897
rect 298695 282863 298753 282897
rect 298787 282863 298816 282897
rect 298660 282832 298816 282863
rect 298660 282353 298816 282384
rect 298660 282319 298661 282353
rect 298695 282319 298753 282353
rect 298787 282319 298816 282353
rect 298660 282288 298816 282319
rect 298660 281809 298816 281840
rect 298660 281775 298661 281809
rect 298695 281775 298753 281809
rect 298787 281775 298816 281809
rect 298660 281744 298816 281775
rect 298660 281265 298816 281296
rect 298660 281231 298661 281265
rect 298695 281231 298753 281265
rect 298787 281231 298816 281265
rect 298660 281200 298816 281231
rect 298660 280721 298816 280752
rect 298660 280687 298661 280721
rect 298695 280687 298753 280721
rect 298787 280687 298816 280721
rect 298660 280656 298816 280687
rect 298660 280177 298816 280208
rect 298660 280143 298661 280177
rect 298695 280143 298753 280177
rect 298787 280143 298816 280177
rect 298660 280112 298816 280143
rect 298660 279633 298816 279664
rect 298660 279599 298661 279633
rect 298695 279599 298753 279633
rect 298787 279599 298816 279633
rect 298660 279568 298816 279599
rect 298660 279089 298816 279120
rect 298660 279055 298661 279089
rect 298695 279055 298753 279089
rect 298787 279055 298816 279089
rect 298660 279024 298816 279055
rect 298660 278545 298816 278576
rect 298660 278511 298661 278545
rect 298695 278511 298753 278545
rect 298787 278511 298816 278545
rect 298660 278480 298816 278511
rect 298660 278001 298816 278032
rect 298660 277967 298661 278001
rect 298695 277967 298753 278001
rect 298787 277967 298816 278001
rect 298660 277936 298816 277967
rect 298660 277457 298816 277488
rect 298660 277423 298661 277457
rect 298695 277423 298753 277457
rect 298787 277423 298816 277457
rect 298660 277392 298816 277423
rect 298660 276913 298816 276944
rect 298660 276879 298661 276913
rect 298695 276879 298753 276913
rect 298787 276879 298816 276913
rect 298660 276848 298816 276879
rect 298660 276369 298816 276400
rect 298660 276335 298661 276369
rect 298695 276335 298753 276369
rect 298787 276335 298816 276369
rect 298660 276304 298816 276335
rect 298660 275825 298816 275856
rect 298660 275791 298661 275825
rect 298695 275791 298753 275825
rect 298787 275791 298816 275825
rect 298660 275760 298816 275791
rect 298660 275281 298816 275312
rect 298660 275247 298661 275281
rect 298695 275247 298753 275281
rect 298787 275247 298816 275281
rect 298660 275216 298816 275247
rect 298660 274737 298816 274768
rect 298660 274703 298661 274737
rect 298695 274703 298753 274737
rect 298787 274703 298816 274737
rect 298660 274672 298816 274703
rect 298660 274193 298816 274224
rect 298660 274159 298661 274193
rect 298695 274159 298753 274193
rect 298787 274159 298816 274193
rect 298660 274128 298816 274159
rect 298660 273649 298816 273680
rect 298660 273615 298661 273649
rect 298695 273615 298753 273649
rect 298787 273615 298816 273649
rect 298660 273584 298816 273615
rect 298660 273105 298816 273136
rect 298660 273071 298661 273105
rect 298695 273071 298753 273105
rect 298787 273071 298816 273105
rect 298660 273040 298816 273071
rect 298660 272561 298816 272592
rect 298660 272527 298661 272561
rect 298695 272527 298753 272561
rect 298787 272527 298816 272561
rect 298660 272496 298816 272527
rect 298660 272017 298816 272048
rect 298660 271983 298661 272017
rect 298695 271983 298753 272017
rect 298787 271983 298816 272017
rect 298660 271952 298816 271983
rect 298660 271473 298816 271504
rect 298660 271439 298661 271473
rect 298695 271439 298753 271473
rect 298787 271439 298816 271473
rect 298660 271408 298816 271439
rect 298660 270929 298816 270960
rect 298660 270895 298661 270929
rect 298695 270895 298753 270929
rect 298787 270895 298816 270929
rect 298660 270864 298816 270895
rect 298660 270385 298816 270416
rect 298660 270351 298661 270385
rect 298695 270351 298753 270385
rect 298787 270351 298816 270385
rect 298660 270320 298816 270351
rect 298660 269841 298816 269872
rect 298660 269807 298661 269841
rect 298695 269807 298753 269841
rect 298787 269807 298816 269841
rect 298660 269776 298816 269807
rect 298660 269297 298816 269328
rect 298660 269263 298661 269297
rect 298695 269263 298753 269297
rect 298787 269263 298816 269297
rect 298660 269232 298816 269263
rect 298660 268753 298816 268784
rect 298660 268719 298661 268753
rect 298695 268719 298753 268753
rect 298787 268719 298816 268753
rect 298660 268688 298816 268719
rect 298660 268209 298816 268240
rect 298660 268175 298661 268209
rect 298695 268175 298753 268209
rect 298787 268175 298816 268209
rect 298660 268144 298816 268175
rect 298660 267665 298816 267696
rect 298660 267631 298661 267665
rect 298695 267631 298753 267665
rect 298787 267631 298816 267665
rect 298660 267600 298816 267631
rect 298660 267121 298816 267152
rect 298660 267087 298661 267121
rect 298695 267087 298753 267121
rect 298787 267087 298816 267121
rect 298660 267056 298816 267087
rect 298660 266577 298816 266608
rect 298660 266543 298661 266577
rect 298695 266543 298753 266577
rect 298787 266543 298816 266577
rect 298660 266512 298816 266543
rect 298660 266033 298816 266064
rect 298660 265999 298661 266033
rect 298695 265999 298753 266033
rect 298787 265999 298816 266033
rect 298660 265968 298816 265999
rect 298660 265489 298816 265520
rect 298660 265455 298661 265489
rect 298695 265455 298753 265489
rect 298787 265455 298816 265489
rect 298660 265424 298816 265455
rect 298660 264945 298816 264976
rect 298660 264911 298661 264945
rect 298695 264911 298753 264945
rect 298787 264911 298816 264945
rect 298660 264880 298816 264911
rect 298660 264401 298816 264432
rect 298660 264367 298661 264401
rect 298695 264367 298753 264401
rect 298787 264367 298816 264401
rect 298660 264336 298816 264367
rect 298660 263857 298816 263888
rect 298660 263823 298661 263857
rect 298695 263823 298753 263857
rect 298787 263823 298816 263857
rect 298660 263792 298816 263823
rect 298660 263313 298816 263344
rect 298660 263279 298661 263313
rect 298695 263279 298753 263313
rect 298787 263279 298816 263313
rect 298660 263248 298816 263279
rect 298660 262769 298816 262800
rect 298660 262735 298661 262769
rect 298695 262735 298753 262769
rect 298787 262735 298816 262769
rect 298660 262704 298816 262735
rect 298660 262225 298816 262256
rect 298660 262191 298661 262225
rect 298695 262191 298753 262225
rect 298787 262191 298816 262225
rect 298660 262160 298816 262191
rect 298660 261681 298816 261712
rect 298660 261647 298661 261681
rect 298695 261647 298753 261681
rect 298787 261647 298816 261681
rect 298660 261616 298816 261647
rect 298660 261137 298816 261168
rect 298660 261103 298661 261137
rect 298695 261103 298753 261137
rect 298787 261103 298816 261137
rect 298660 261072 298816 261103
rect 298660 260593 298816 260624
rect 298660 260559 298661 260593
rect 298695 260559 298753 260593
rect 298787 260559 298816 260593
rect 298660 260528 298816 260559
rect 298660 260049 298816 260080
rect 298660 260015 298661 260049
rect 298695 260015 298753 260049
rect 298787 260015 298816 260049
rect 298660 259984 298816 260015
rect 298660 259505 298816 259536
rect 298660 259471 298661 259505
rect 298695 259471 298753 259505
rect 298787 259471 298816 259505
rect 298660 259440 298816 259471
rect 298660 258961 298816 258992
rect 298660 258927 298661 258961
rect 298695 258927 298753 258961
rect 298787 258927 298816 258961
rect 298660 258896 298816 258927
rect 298660 258417 298816 258448
rect 298660 258383 298661 258417
rect 298695 258383 298753 258417
rect 298787 258383 298816 258417
rect 298660 258352 298816 258383
rect 298660 257873 298816 257904
rect 298660 257839 298661 257873
rect 298695 257839 298753 257873
rect 298787 257839 298816 257873
rect 298660 257808 298816 257839
rect 298660 257329 298816 257360
rect 298660 257295 298661 257329
rect 298695 257295 298753 257329
rect 298787 257295 298816 257329
rect 298660 257264 298816 257295
rect 298660 256785 298816 256816
rect 298660 256751 298661 256785
rect 298695 256751 298753 256785
rect 298787 256751 298816 256785
rect 298660 256720 298816 256751
rect 298660 256241 298816 256272
rect 298660 256207 298661 256241
rect 298695 256207 298753 256241
rect 298787 256207 298816 256241
rect 298660 256176 298816 256207
rect 298660 255697 298816 255728
rect 298660 255663 298661 255697
rect 298695 255663 298753 255697
rect 298787 255663 298816 255697
rect 298660 255632 298816 255663
rect 298660 255153 298816 255184
rect 298660 255119 298661 255153
rect 298695 255119 298753 255153
rect 298787 255119 298816 255153
rect 298660 255088 298816 255119
rect 298660 254609 298816 254640
rect 298660 254575 298661 254609
rect 298695 254575 298753 254609
rect 298787 254575 298816 254609
rect 298660 254544 298816 254575
rect 298660 254065 298816 254096
rect 298660 254031 298661 254065
rect 298695 254031 298753 254065
rect 298787 254031 298816 254065
rect 298660 254000 298816 254031
rect 298660 253521 298816 253552
rect 298660 253487 298661 253521
rect 298695 253487 298753 253521
rect 298787 253487 298816 253521
rect 298660 253456 298816 253487
rect 298660 252977 298816 253008
rect 298660 252943 298661 252977
rect 298695 252943 298753 252977
rect 298787 252943 298816 252977
rect 298660 252912 298816 252943
rect 298660 252433 298816 252464
rect 298660 252399 298661 252433
rect 298695 252399 298753 252433
rect 298787 252399 298816 252433
rect 298660 252368 298816 252399
rect 298660 251889 298816 251920
rect 298660 251855 298661 251889
rect 298695 251855 298753 251889
rect 298787 251855 298816 251889
rect 298660 251824 298816 251855
rect 298660 251345 298816 251376
rect 298660 251311 298661 251345
rect 298695 251311 298753 251345
rect 298787 251311 298816 251345
rect 298660 251280 298816 251311
rect 298660 250801 298816 250832
rect 298660 250767 298661 250801
rect 298695 250767 298753 250801
rect 298787 250767 298816 250801
rect 298660 250736 298816 250767
rect 298660 250257 298816 250288
rect 298660 250223 298661 250257
rect 298695 250223 298753 250257
rect 298787 250223 298816 250257
rect 298660 250192 298816 250223
rect 298660 249713 298816 249744
rect 298660 249679 298661 249713
rect 298695 249679 298753 249713
rect 298787 249679 298816 249713
rect 298660 249648 298816 249679
rect 298660 249169 298816 249200
rect 298660 249135 298661 249169
rect 298695 249135 298753 249169
rect 298787 249135 298816 249169
rect 298660 249104 298816 249135
rect 298660 248625 298816 248656
rect 298660 248591 298661 248625
rect 298695 248591 298753 248625
rect 298787 248591 298816 248625
rect 298660 248560 298816 248591
rect 298660 248081 298816 248112
rect 298660 248047 298661 248081
rect 298695 248047 298753 248081
rect 298787 248047 298816 248081
rect 298660 248016 298816 248047
rect 298660 247537 298816 247568
rect 298660 247503 298661 247537
rect 298695 247503 298753 247537
rect 298787 247503 298816 247537
rect 298660 247472 298816 247503
rect 298660 246993 298816 247024
rect 298660 246959 298661 246993
rect 298695 246959 298753 246993
rect 298787 246959 298816 246993
rect 298660 246928 298816 246959
rect 298660 246449 298816 246480
rect 298660 246415 298661 246449
rect 298695 246415 298753 246449
rect 298787 246415 298816 246449
rect 298660 246384 298816 246415
rect 298660 245905 298816 245936
rect 298660 245871 298661 245905
rect 298695 245871 298753 245905
rect 298787 245871 298816 245905
rect 298660 245840 298816 245871
rect 298660 245361 298816 245392
rect 298660 245327 298661 245361
rect 298695 245327 298753 245361
rect 298787 245327 298816 245361
rect 298660 245296 298816 245327
rect 298660 244817 298816 244848
rect 298660 244783 298661 244817
rect 298695 244783 298753 244817
rect 298787 244783 298816 244817
rect 298660 244752 298816 244783
rect 298660 244273 298816 244304
rect 298660 244239 298661 244273
rect 298695 244239 298753 244273
rect 298787 244239 298816 244273
rect 298660 244208 298816 244239
rect 298660 243729 298816 243760
rect 298660 243695 298661 243729
rect 298695 243695 298753 243729
rect 298787 243695 298816 243729
rect 298660 243664 298816 243695
rect 298660 243185 298816 243216
rect 298660 243151 298661 243185
rect 298695 243151 298753 243185
rect 298787 243151 298816 243185
rect 298660 243120 298816 243151
rect 298660 242641 298816 242672
rect 298660 242607 298661 242641
rect 298695 242607 298753 242641
rect 298787 242607 298816 242641
rect 298660 242576 298816 242607
rect 298660 242097 298816 242128
rect 298660 242063 298661 242097
rect 298695 242063 298753 242097
rect 298787 242063 298816 242097
rect 298660 242032 298816 242063
rect 298660 241553 298816 241584
rect 298660 241519 298661 241553
rect 298695 241519 298753 241553
rect 298787 241519 298816 241553
rect 298660 241488 298816 241519
rect 298660 241009 298816 241040
rect 298660 240975 298661 241009
rect 298695 240975 298753 241009
rect 298787 240975 298816 241009
rect 298660 240944 298816 240975
rect 298660 240465 298816 240496
rect 298660 240431 298661 240465
rect 298695 240431 298753 240465
rect 298787 240431 298816 240465
rect 298660 240400 298816 240431
rect 298660 239921 298816 239952
rect 298660 239887 298661 239921
rect 298695 239887 298753 239921
rect 298787 239887 298816 239921
rect 298660 239856 298816 239887
rect 298660 239377 298816 239408
rect 298660 239343 298661 239377
rect 298695 239343 298753 239377
rect 298787 239343 298816 239377
rect 298660 239312 298816 239343
rect 298660 238833 298816 238864
rect 298660 238799 298661 238833
rect 298695 238799 298753 238833
rect 298787 238799 298816 238833
rect 298660 238768 298816 238799
rect 298660 238289 298816 238320
rect 298660 238255 298661 238289
rect 298695 238255 298753 238289
rect 298787 238255 298816 238289
rect 298660 238224 298816 238255
rect 298660 237745 298816 237776
rect 298660 237711 298661 237745
rect 298695 237711 298753 237745
rect 298787 237711 298816 237745
rect 298660 237680 298816 237711
rect 298660 237201 298816 237232
rect 298660 237167 298661 237201
rect 298695 237167 298753 237201
rect 298787 237167 298816 237201
rect 298660 237136 298816 237167
rect 298660 236657 298816 236688
rect 298660 236623 298661 236657
rect 298695 236623 298753 236657
rect 298787 236623 298816 236657
rect 298660 236592 298816 236623
rect 298660 236113 298816 236144
rect 298660 236079 298661 236113
rect 298695 236079 298753 236113
rect 298787 236079 298816 236113
rect 298660 236048 298816 236079
rect 298660 235569 298816 235600
rect 298660 235535 298661 235569
rect 298695 235535 298753 235569
rect 298787 235535 298816 235569
rect 298660 235504 298816 235535
rect 298660 235025 298816 235056
rect 298660 234991 298661 235025
rect 298695 234991 298753 235025
rect 298787 234991 298816 235025
rect 298660 234960 298816 234991
rect 298660 234481 298816 234512
rect 298660 234447 298661 234481
rect 298695 234447 298753 234481
rect 298787 234447 298816 234481
rect 298660 234416 298816 234447
rect 298660 233937 298816 233968
rect 298660 233903 298661 233937
rect 298695 233903 298753 233937
rect 298787 233903 298816 233937
rect 298660 233872 298816 233903
rect 298660 233393 298816 233424
rect 298660 233359 298661 233393
rect 298695 233359 298753 233393
rect 298787 233359 298816 233393
rect 298660 233328 298816 233359
rect 298660 232849 298816 232880
rect 298660 232815 298661 232849
rect 298695 232815 298753 232849
rect 298787 232815 298816 232849
rect 298660 232784 298816 232815
rect 298660 232305 298816 232336
rect 298660 232271 298661 232305
rect 298695 232271 298753 232305
rect 298787 232271 298816 232305
rect 298660 232240 298816 232271
rect 298660 231761 298816 231792
rect 298660 231727 298661 231761
rect 298695 231727 298753 231761
rect 298787 231727 298816 231761
rect 298660 231696 298816 231727
rect 298660 231217 298816 231248
rect 298660 231183 298661 231217
rect 298695 231183 298753 231217
rect 298787 231183 298816 231217
rect 298660 231152 298816 231183
rect 298660 230673 298816 230704
rect 298660 230639 298661 230673
rect 298695 230639 298753 230673
rect 298787 230639 298816 230673
rect 298660 230608 298816 230639
rect 298660 230129 298816 230160
rect 298660 230095 298661 230129
rect 298695 230095 298753 230129
rect 298787 230095 298816 230129
rect 298660 230064 298816 230095
rect 298660 229585 298816 229616
rect 298660 229551 298661 229585
rect 298695 229551 298753 229585
rect 298787 229551 298816 229585
rect 298660 229520 298816 229551
rect 298660 229041 298816 229072
rect 298660 229007 298661 229041
rect 298695 229007 298753 229041
rect 298787 229007 298816 229041
rect 298660 228976 298816 229007
rect 298660 228497 298816 228528
rect 298660 228463 298661 228497
rect 298695 228463 298753 228497
rect 298787 228463 298816 228497
rect 298660 228432 298816 228463
rect 298660 227953 298816 227984
rect 298660 227919 298661 227953
rect 298695 227919 298753 227953
rect 298787 227919 298816 227953
rect 298660 227888 298816 227919
rect 298660 227409 298816 227440
rect 298660 227375 298661 227409
rect 298695 227375 298753 227409
rect 298787 227375 298816 227409
rect 298660 227344 298816 227375
rect 298660 226865 298816 226896
rect 298660 226831 298661 226865
rect 298695 226831 298753 226865
rect 298787 226831 298816 226865
rect 298660 226800 298816 226831
rect 298660 226321 298816 226352
rect 298660 226287 298661 226321
rect 298695 226287 298753 226321
rect 298787 226287 298816 226321
rect 298660 226256 298816 226287
rect 298660 225777 298816 225808
rect 298660 225743 298661 225777
rect 298695 225743 298753 225777
rect 298787 225743 298816 225777
rect 298660 225712 298816 225743
rect 298660 225233 298816 225264
rect 298660 225199 298661 225233
rect 298695 225199 298753 225233
rect 298787 225199 298816 225233
rect 298660 225168 298816 225199
rect 298660 224689 298816 224720
rect 298660 224655 298661 224689
rect 298695 224655 298753 224689
rect 298787 224655 298816 224689
rect 298660 224624 298816 224655
rect 298660 224145 298816 224176
rect 298660 224111 298661 224145
rect 298695 224111 298753 224145
rect 298787 224111 298816 224145
rect 298660 224080 298816 224111
rect 298660 223601 298816 223632
rect 298660 223567 298661 223601
rect 298695 223567 298753 223601
rect 298787 223567 298816 223601
rect 298660 223536 298816 223567
rect 298660 223057 298816 223088
rect 298660 223023 298661 223057
rect 298695 223023 298753 223057
rect 298787 223023 298816 223057
rect 298660 222992 298816 223023
rect 298660 222513 298816 222544
rect 298660 222479 298661 222513
rect 298695 222479 298753 222513
rect 298787 222479 298816 222513
rect 298660 222448 298816 222479
rect 298660 221969 298816 222000
rect 298660 221935 298661 221969
rect 298695 221935 298753 221969
rect 298787 221935 298816 221969
rect 298660 221904 298816 221935
rect 298660 221425 298816 221456
rect 298660 221391 298661 221425
rect 298695 221391 298753 221425
rect 298787 221391 298816 221425
rect 298660 221360 298816 221391
rect 298660 220881 298816 220912
rect 298660 220847 298661 220881
rect 298695 220847 298753 220881
rect 298787 220847 298816 220881
rect 298660 220816 298816 220847
rect 298660 220337 298816 220368
rect 298660 220303 298661 220337
rect 298695 220303 298753 220337
rect 298787 220303 298816 220337
rect 298660 220272 298816 220303
rect 298660 219793 298816 219824
rect 298660 219759 298661 219793
rect 298695 219759 298753 219793
rect 298787 219759 298816 219793
rect 298660 219728 298816 219759
rect 298660 219249 298816 219280
rect 298660 219215 298661 219249
rect 298695 219215 298753 219249
rect 298787 219215 298816 219249
rect 298660 219184 298816 219215
rect 298660 218705 298816 218736
rect 298660 218671 298661 218705
rect 298695 218671 298753 218705
rect 298787 218671 298816 218705
rect 298660 218640 298816 218671
rect 298660 218161 298816 218192
rect 298660 218127 298661 218161
rect 298695 218127 298753 218161
rect 298787 218127 298816 218161
rect 298660 218096 298816 218127
rect 298660 217617 298816 217648
rect 298660 217583 298661 217617
rect 298695 217583 298753 217617
rect 298787 217583 298816 217617
rect 298660 217552 298816 217583
rect 298660 217073 298816 217104
rect 298660 217039 298661 217073
rect 298695 217039 298753 217073
rect 298787 217039 298816 217073
rect 298660 217008 298816 217039
rect 298660 216529 298816 216560
rect 298660 216495 298661 216529
rect 298695 216495 298753 216529
rect 298787 216495 298816 216529
rect 298660 216464 298816 216495
rect 298660 215985 298816 216016
rect 298660 215951 298661 215985
rect 298695 215951 298753 215985
rect 298787 215951 298816 215985
rect 298660 215920 298816 215951
rect 298660 215441 298816 215472
rect 298660 215407 298661 215441
rect 298695 215407 298753 215441
rect 298787 215407 298816 215441
rect 298660 215376 298816 215407
rect 298660 214897 298816 214928
rect 298660 214863 298661 214897
rect 298695 214863 298753 214897
rect 298787 214863 298816 214897
rect 298660 214832 298816 214863
rect 298660 214353 298816 214384
rect 298660 214319 298661 214353
rect 298695 214319 298753 214353
rect 298787 214319 298816 214353
rect 298660 214288 298816 214319
rect 298660 213809 298816 213840
rect 298660 213775 298661 213809
rect 298695 213775 298753 213809
rect 298787 213775 298816 213809
rect 298660 213744 298816 213775
rect 298660 213265 298816 213296
rect 298660 213231 298661 213265
rect 298695 213231 298753 213265
rect 298787 213231 298816 213265
rect 298660 213200 298816 213231
rect 298660 212721 298816 212752
rect 298660 212687 298661 212721
rect 298695 212687 298753 212721
rect 298787 212687 298816 212721
rect 298660 212656 298816 212687
rect 298660 212177 298816 212208
rect 298660 212143 298661 212177
rect 298695 212143 298753 212177
rect 298787 212143 298816 212177
rect 298660 212112 298816 212143
rect 298660 211633 298816 211664
rect 298660 211599 298661 211633
rect 298695 211599 298753 211633
rect 298787 211599 298816 211633
rect 298660 211568 298816 211599
rect 298660 211089 298816 211120
rect 298660 211055 298661 211089
rect 298695 211055 298753 211089
rect 298787 211055 298816 211089
rect 298660 211024 298816 211055
rect 298660 210545 298816 210576
rect 298660 210511 298661 210545
rect 298695 210511 298753 210545
rect 298787 210511 298816 210545
rect 298660 210480 298816 210511
rect 298660 210001 298816 210032
rect 298660 209967 298661 210001
rect 298695 209967 298753 210001
rect 298787 209967 298816 210001
rect 298660 209936 298816 209967
rect 298660 209457 298816 209488
rect 298660 209423 298661 209457
rect 298695 209423 298753 209457
rect 298787 209423 298816 209457
rect 298660 209392 298816 209423
rect 298660 208913 298816 208944
rect 298660 208879 298661 208913
rect 298695 208879 298753 208913
rect 298787 208879 298816 208913
rect 298660 208848 298816 208879
rect 298660 208369 298816 208400
rect 298660 208335 298661 208369
rect 298695 208335 298753 208369
rect 298787 208335 298816 208369
rect 298660 208304 298816 208335
rect 298660 207825 298816 207856
rect 298660 207791 298661 207825
rect 298695 207791 298753 207825
rect 298787 207791 298816 207825
rect 298660 207760 298816 207791
rect 298660 207281 298816 207312
rect 298660 207247 298661 207281
rect 298695 207247 298753 207281
rect 298787 207247 298816 207281
rect 298660 207216 298816 207247
rect 298660 206737 298816 206768
rect 298660 206703 298661 206737
rect 298695 206703 298753 206737
rect 298787 206703 298816 206737
rect 298660 206672 298816 206703
rect 298660 206193 298816 206224
rect 298660 206159 298661 206193
rect 298695 206159 298753 206193
rect 298787 206159 298816 206193
rect 298660 206128 298816 206159
rect 298660 205649 298816 205680
rect 298660 205615 298661 205649
rect 298695 205615 298753 205649
rect 298787 205615 298816 205649
rect 298660 205584 298816 205615
rect 298660 205105 298816 205136
rect 298660 205071 298661 205105
rect 298695 205071 298753 205105
rect 298787 205071 298816 205105
rect 298660 205040 298816 205071
rect 298660 204561 298816 204592
rect 298660 204527 298661 204561
rect 298695 204527 298753 204561
rect 298787 204527 298816 204561
rect 298660 204496 298816 204527
rect 298660 204017 298816 204048
rect 298660 203983 298661 204017
rect 298695 203983 298753 204017
rect 298787 203983 298816 204017
rect 298660 203952 298816 203983
rect 298660 203473 298816 203504
rect 298660 203439 298661 203473
rect 298695 203439 298753 203473
rect 298787 203439 298816 203473
rect 298660 203408 298816 203439
rect 298660 202929 298816 202960
rect 298660 202895 298661 202929
rect 298695 202895 298753 202929
rect 298787 202895 298816 202929
rect 298660 202864 298816 202895
rect 298660 202385 298816 202416
rect 298660 202351 298661 202385
rect 298695 202351 298753 202385
rect 298787 202351 298816 202385
rect 298660 202320 298816 202351
rect 298660 201841 298816 201872
rect 298660 201807 298661 201841
rect 298695 201807 298753 201841
rect 298787 201807 298816 201841
rect 298660 201776 298816 201807
rect 298660 201297 298816 201328
rect 298660 201263 298661 201297
rect 298695 201263 298753 201297
rect 298787 201263 298816 201297
rect 298660 201232 298816 201263
rect 298660 200753 298816 200784
rect 298660 200719 298661 200753
rect 298695 200719 298753 200753
rect 298787 200719 298816 200753
rect 298660 200688 298816 200719
rect 298660 200209 298816 200240
rect 298660 200175 298661 200209
rect 298695 200175 298753 200209
rect 298787 200175 298816 200209
rect 298660 200144 298816 200175
rect 298660 199665 298816 199696
rect 298660 199631 298661 199665
rect 298695 199631 298753 199665
rect 298787 199631 298816 199665
rect 298660 199600 298816 199631
rect 298660 199121 298816 199152
rect 298660 199087 298661 199121
rect 298695 199087 298753 199121
rect 298787 199087 298816 199121
rect 298660 199056 298816 199087
rect 298660 198577 298816 198608
rect 298660 198543 298661 198577
rect 298695 198543 298753 198577
rect 298787 198543 298816 198577
rect 298660 198512 298816 198543
rect 298660 198033 298816 198064
rect 298660 197999 298661 198033
rect 298695 197999 298753 198033
rect 298787 197999 298816 198033
rect 298660 197968 298816 197999
rect 298660 197489 298816 197520
rect 298660 197455 298661 197489
rect 298695 197455 298753 197489
rect 298787 197455 298816 197489
rect 298660 197424 298816 197455
rect 298660 196945 298816 196976
rect 298660 196911 298661 196945
rect 298695 196911 298753 196945
rect 298787 196911 298816 196945
rect 298660 196880 298816 196911
rect 298660 196401 298816 196432
rect 298660 196367 298661 196401
rect 298695 196367 298753 196401
rect 298787 196367 298816 196401
rect 298660 196336 298816 196367
rect 298660 195857 298816 195888
rect 298660 195823 298661 195857
rect 298695 195823 298753 195857
rect 298787 195823 298816 195857
rect 298660 195792 298816 195823
rect 298660 195313 298816 195344
rect 298660 195279 298661 195313
rect 298695 195279 298753 195313
rect 298787 195279 298816 195313
rect 298660 195248 298816 195279
rect 298660 194769 298816 194800
rect 298660 194735 298661 194769
rect 298695 194735 298753 194769
rect 298787 194735 298816 194769
rect 298660 194704 298816 194735
rect 298660 194225 298816 194256
rect 298660 194191 298661 194225
rect 298695 194191 298753 194225
rect 298787 194191 298816 194225
rect 298660 194160 298816 194191
rect 298660 193681 298816 193712
rect 298660 193647 298661 193681
rect 298695 193647 298753 193681
rect 298787 193647 298816 193681
rect 298660 193616 298816 193647
rect 298660 193137 298816 193168
rect 298660 193103 298661 193137
rect 298695 193103 298753 193137
rect 298787 193103 298816 193137
rect 298660 193072 298816 193103
rect 298660 192593 298816 192624
rect 298660 192559 298661 192593
rect 298695 192559 298753 192593
rect 298787 192559 298816 192593
rect 298660 192528 298816 192559
rect 298660 192049 298816 192080
rect 298660 192015 298661 192049
rect 298695 192015 298753 192049
rect 298787 192015 298816 192049
rect 298660 191984 298816 192015
rect 298660 191505 298816 191536
rect 298660 191471 298661 191505
rect 298695 191471 298753 191505
rect 298787 191471 298816 191505
rect 298660 191440 298816 191471
rect 298660 190961 298816 190992
rect 298660 190927 298661 190961
rect 298695 190927 298753 190961
rect 298787 190927 298816 190961
rect 298660 190896 298816 190927
rect 298660 190417 298816 190448
rect 298660 190383 298661 190417
rect 298695 190383 298753 190417
rect 298787 190383 298816 190417
rect 298660 190352 298816 190383
rect 298660 189873 298816 189904
rect 298660 189839 298661 189873
rect 298695 189839 298753 189873
rect 298787 189839 298816 189873
rect 298660 189808 298816 189839
rect 298660 189329 298816 189360
rect 298660 189295 298661 189329
rect 298695 189295 298753 189329
rect 298787 189295 298816 189329
rect 298660 189264 298816 189295
rect 298660 188785 298816 188816
rect 298660 188751 298661 188785
rect 298695 188751 298753 188785
rect 298787 188751 298816 188785
rect 298660 188720 298816 188751
rect 298660 188241 298816 188272
rect 298660 188207 298661 188241
rect 298695 188207 298753 188241
rect 298787 188207 298816 188241
rect 298660 188176 298816 188207
rect 298660 187697 298816 187728
rect 298660 187663 298661 187697
rect 298695 187663 298753 187697
rect 298787 187663 298816 187697
rect 298660 187632 298816 187663
rect 298660 187153 298816 187184
rect 298660 187119 298661 187153
rect 298695 187119 298753 187153
rect 298787 187119 298816 187153
rect 298660 187088 298816 187119
rect 298660 186609 298816 186640
rect 298660 186575 298661 186609
rect 298695 186575 298753 186609
rect 298787 186575 298816 186609
rect 298660 186544 298816 186575
rect 298660 186065 298816 186096
rect 298660 186031 298661 186065
rect 298695 186031 298753 186065
rect 298787 186031 298816 186065
rect 298660 186000 298816 186031
rect 298660 185521 298816 185552
rect 298660 185487 298661 185521
rect 298695 185487 298753 185521
rect 298787 185487 298816 185521
rect 298660 185456 298816 185487
rect 298660 184977 298816 185008
rect 298660 184943 298661 184977
rect 298695 184943 298753 184977
rect 298787 184943 298816 184977
rect 298660 184912 298816 184943
rect 298660 184433 298816 184464
rect 298660 184399 298661 184433
rect 298695 184399 298753 184433
rect 298787 184399 298816 184433
rect 298660 184368 298816 184399
rect 298660 183889 298816 183920
rect 298660 183855 298661 183889
rect 298695 183855 298753 183889
rect 298787 183855 298816 183889
rect 298660 183824 298816 183855
rect 298660 183345 298816 183376
rect 298660 183311 298661 183345
rect 298695 183311 298753 183345
rect 298787 183311 298816 183345
rect 298660 183280 298816 183311
rect 298660 182801 298816 182832
rect 298660 182767 298661 182801
rect 298695 182767 298753 182801
rect 298787 182767 298816 182801
rect 298660 182736 298816 182767
rect 298660 182257 298816 182288
rect 298660 182223 298661 182257
rect 298695 182223 298753 182257
rect 298787 182223 298816 182257
rect 298660 182192 298816 182223
rect 298660 181713 298816 181744
rect 298660 181679 298661 181713
rect 298695 181679 298753 181713
rect 298787 181679 298816 181713
rect 298660 181648 298816 181679
rect 298660 181169 298816 181200
rect 298660 181135 298661 181169
rect 298695 181135 298753 181169
rect 298787 181135 298816 181169
rect 298660 181104 298816 181135
rect 298660 180625 298816 180656
rect 298660 180591 298661 180625
rect 298695 180591 298753 180625
rect 298787 180591 298816 180625
rect 298660 180560 298816 180591
rect 298660 180081 298816 180112
rect 298660 180047 298661 180081
rect 298695 180047 298753 180081
rect 298787 180047 298816 180081
rect 298660 180016 298816 180047
rect 298660 179537 298816 179568
rect 298660 179503 298661 179537
rect 298695 179503 298753 179537
rect 298787 179503 298816 179537
rect 298660 179472 298816 179503
rect 298660 178993 298816 179024
rect 298660 178959 298661 178993
rect 298695 178959 298753 178993
rect 298787 178959 298816 178993
rect 298660 178928 298816 178959
rect 298660 178449 298816 178480
rect 298660 178415 298661 178449
rect 298695 178415 298753 178449
rect 298787 178415 298816 178449
rect 298660 178384 298816 178415
rect 298660 177905 298816 177936
rect 298660 177871 298661 177905
rect 298695 177871 298753 177905
rect 298787 177871 298816 177905
rect 298660 177840 298816 177871
rect 298660 177361 298816 177392
rect 298660 177327 298661 177361
rect 298695 177327 298753 177361
rect 298787 177327 298816 177361
rect 298660 177296 298816 177327
rect 298660 176817 298816 176848
rect 298660 176783 298661 176817
rect 298695 176783 298753 176817
rect 298787 176783 298816 176817
rect 298660 176752 298816 176783
rect 298660 176273 298816 176304
rect 298660 176239 298661 176273
rect 298695 176239 298753 176273
rect 298787 176239 298816 176273
rect 298660 176208 298816 176239
rect 298660 175729 298816 175760
rect 298660 175695 298661 175729
rect 298695 175695 298753 175729
rect 298787 175695 298816 175729
rect 298660 175664 298816 175695
rect 298660 175185 298816 175216
rect 298660 175151 298661 175185
rect 298695 175151 298753 175185
rect 298787 175151 298816 175185
rect 298660 175120 298816 175151
rect 298660 174641 298816 174672
rect 298660 174607 298661 174641
rect 298695 174607 298753 174641
rect 298787 174607 298816 174641
rect 298660 174576 298816 174607
rect 298660 174097 298816 174128
rect 298660 174063 298661 174097
rect 298695 174063 298753 174097
rect 298787 174063 298816 174097
rect 298660 174032 298816 174063
rect 298660 173553 298816 173584
rect 298660 173519 298661 173553
rect 298695 173519 298753 173553
rect 298787 173519 298816 173553
rect 298660 173488 298816 173519
rect 298660 173009 298816 173040
rect 298660 172975 298661 173009
rect 298695 172975 298753 173009
rect 298787 172975 298816 173009
rect 298660 172944 298816 172975
rect 298660 172465 298816 172496
rect 298660 172431 298661 172465
rect 298695 172431 298753 172465
rect 298787 172431 298816 172465
rect 298660 172400 298816 172431
rect 298660 171921 298816 171952
rect 298660 171887 298661 171921
rect 298695 171887 298753 171921
rect 298787 171887 298816 171921
rect 298660 171856 298816 171887
rect 298660 171377 298816 171408
rect 298660 171343 298661 171377
rect 298695 171343 298753 171377
rect 298787 171343 298816 171377
rect 298660 171312 298816 171343
rect 298660 170833 298816 170864
rect 298660 170799 298661 170833
rect 298695 170799 298753 170833
rect 298787 170799 298816 170833
rect 298660 170768 298816 170799
rect 298660 170289 298816 170320
rect 298660 170255 298661 170289
rect 298695 170255 298753 170289
rect 298787 170255 298816 170289
rect 298660 170224 298816 170255
rect 298660 169745 298816 169776
rect 298660 169711 298661 169745
rect 298695 169711 298753 169745
rect 298787 169711 298816 169745
rect 298660 169680 298816 169711
rect 298660 169201 298816 169232
rect 298660 169167 298661 169201
rect 298695 169167 298753 169201
rect 298787 169167 298816 169201
rect 298660 169136 298816 169167
rect 298660 168657 298816 168688
rect 298660 168623 298661 168657
rect 298695 168623 298753 168657
rect 298787 168623 298816 168657
rect 298660 168592 298816 168623
rect 298660 168113 298816 168144
rect 298660 168079 298661 168113
rect 298695 168079 298753 168113
rect 298787 168079 298816 168113
rect 298660 168048 298816 168079
rect 298660 167569 298816 167600
rect 298660 167535 298661 167569
rect 298695 167535 298753 167569
rect 298787 167535 298816 167569
rect 298660 167504 298816 167535
rect 298660 167025 298816 167056
rect 298660 166991 298661 167025
rect 298695 166991 298753 167025
rect 298787 166991 298816 167025
rect 298660 166960 298816 166991
rect 298660 166481 298816 166512
rect 298660 166447 298661 166481
rect 298695 166447 298753 166481
rect 298787 166447 298816 166481
rect 298660 166416 298816 166447
rect 298660 165937 298816 165968
rect 298660 165903 298661 165937
rect 298695 165903 298753 165937
rect 298787 165903 298816 165937
rect 298660 165872 298816 165903
rect 298660 165393 298816 165424
rect 298660 165359 298661 165393
rect 298695 165359 298753 165393
rect 298787 165359 298816 165393
rect 298660 165328 298816 165359
rect 298660 164849 298816 164880
rect 298660 164815 298661 164849
rect 298695 164815 298753 164849
rect 298787 164815 298816 164849
rect 298660 164784 298816 164815
rect 298660 164305 298816 164336
rect 298660 164271 298661 164305
rect 298695 164271 298753 164305
rect 298787 164271 298816 164305
rect 298660 164240 298816 164271
rect 298660 163761 298816 163792
rect 298660 163727 298661 163761
rect 298695 163727 298753 163761
rect 298787 163727 298816 163761
rect 298660 163696 298816 163727
rect 298660 163217 298816 163248
rect 298660 163183 298661 163217
rect 298695 163183 298753 163217
rect 298787 163183 298816 163217
rect 298660 163152 298816 163183
rect 298660 162673 298816 162704
rect 298660 162639 298661 162673
rect 298695 162639 298753 162673
rect 298787 162639 298816 162673
rect 298660 162608 298816 162639
rect 298660 162129 298816 162160
rect 298660 162095 298661 162129
rect 298695 162095 298753 162129
rect 298787 162095 298816 162129
rect 298660 162064 298816 162095
rect 298660 161585 298816 161616
rect 298660 161551 298661 161585
rect 298695 161551 298753 161585
rect 298787 161551 298816 161585
rect 298660 161520 298816 161551
rect 298660 161041 298816 161072
rect 298660 161007 298661 161041
rect 298695 161007 298753 161041
rect 298787 161007 298816 161041
rect 298660 160976 298816 161007
rect 298660 160497 298816 160528
rect 298660 160463 298661 160497
rect 298695 160463 298753 160497
rect 298787 160463 298816 160497
rect 298660 160432 298816 160463
rect 298660 159953 298816 159984
rect 298660 159919 298661 159953
rect 298695 159919 298753 159953
rect 298787 159919 298816 159953
rect 298660 159888 298816 159919
rect 298660 159409 298816 159440
rect 298660 159375 298661 159409
rect 298695 159375 298753 159409
rect 298787 159375 298816 159409
rect 298660 159344 298816 159375
rect 298660 158865 298816 158896
rect 298660 158831 298661 158865
rect 298695 158831 298753 158865
rect 298787 158831 298816 158865
rect 298660 158800 298816 158831
rect 298660 158321 298816 158352
rect 298660 158287 298661 158321
rect 298695 158287 298753 158321
rect 298787 158287 298816 158321
rect 298660 158256 298816 158287
rect 298660 157777 298816 157808
rect 298660 157743 298661 157777
rect 298695 157743 298753 157777
rect 298787 157743 298816 157777
rect 298660 157712 298816 157743
rect 298660 157233 298816 157264
rect 298660 157199 298661 157233
rect 298695 157199 298753 157233
rect 298787 157199 298816 157233
rect 298660 157168 298816 157199
rect 298660 156689 298816 156720
rect 298660 156655 298661 156689
rect 298695 156655 298753 156689
rect 298787 156655 298816 156689
rect 298660 156624 298816 156655
rect 298660 156145 298816 156176
rect 298660 156111 298661 156145
rect 298695 156111 298753 156145
rect 298787 156111 298816 156145
rect 298660 156080 298816 156111
rect 298660 155601 298816 155632
rect 298660 155567 298661 155601
rect 298695 155567 298753 155601
rect 298787 155567 298816 155601
rect 298660 155536 298816 155567
rect 298660 155057 298816 155088
rect 298660 155023 298661 155057
rect 298695 155023 298753 155057
rect 298787 155023 298816 155057
rect 298660 154992 298816 155023
rect 298660 154513 298816 154544
rect 298660 154479 298661 154513
rect 298695 154479 298753 154513
rect 298787 154479 298816 154513
rect 298660 154448 298816 154479
rect 298660 153969 298816 154000
rect 298660 153935 298661 153969
rect 298695 153935 298753 153969
rect 298787 153935 298816 153969
rect 298660 153904 298816 153935
rect 298660 153425 298816 153456
rect 298660 153391 298661 153425
rect 298695 153391 298753 153425
rect 298787 153391 298816 153425
rect 298660 153360 298816 153391
rect 298660 152881 298816 152912
rect 298660 152847 298661 152881
rect 298695 152847 298753 152881
rect 298787 152847 298816 152881
rect 298660 152816 298816 152847
rect 298660 152337 298816 152368
rect 298660 152303 298661 152337
rect 298695 152303 298753 152337
rect 298787 152303 298816 152337
rect 298660 152272 298816 152303
rect 298660 151793 298816 151824
rect 298660 151759 298661 151793
rect 298695 151759 298753 151793
rect 298787 151759 298816 151793
rect 298660 151728 298816 151759
rect 298660 151249 298816 151280
rect 298660 151215 298661 151249
rect 298695 151215 298753 151249
rect 298787 151215 298816 151249
rect 298660 151184 298816 151215
rect 298660 150705 298816 150736
rect 298660 150671 298661 150705
rect 298695 150671 298753 150705
rect 298787 150671 298816 150705
rect 298660 150640 298816 150671
rect 298660 150161 298816 150192
rect 298660 150127 298661 150161
rect 298695 150127 298753 150161
rect 298787 150127 298816 150161
rect 298660 150096 298816 150127
rect 298660 149617 298816 149648
rect 298660 149583 298661 149617
rect 298695 149583 298753 149617
rect 298787 149583 298816 149617
rect 298660 149552 298816 149583
rect 298660 149073 298816 149104
rect 298660 149039 298661 149073
rect 298695 149039 298753 149073
rect 298787 149039 298816 149073
rect 298660 149008 298816 149039
rect 298660 148529 298816 148560
rect 298660 148495 298661 148529
rect 298695 148495 298753 148529
rect 298787 148495 298816 148529
rect 298660 148464 298816 148495
rect 298660 147985 298816 148016
rect 298660 147951 298661 147985
rect 298695 147951 298753 147985
rect 298787 147951 298816 147985
rect 298660 147920 298816 147951
rect 298660 147441 298816 147472
rect 298660 147407 298661 147441
rect 298695 147407 298753 147441
rect 298787 147407 298816 147441
rect 298660 147376 298816 147407
rect 298660 146897 298816 146928
rect 298660 146863 298661 146897
rect 298695 146863 298753 146897
rect 298787 146863 298816 146897
rect 298660 146832 298816 146863
rect 298660 146353 298816 146384
rect 298660 146319 298661 146353
rect 298695 146319 298753 146353
rect 298787 146319 298816 146353
rect 298660 146288 298816 146319
rect 298660 145809 298816 145840
rect 298660 145775 298661 145809
rect 298695 145775 298753 145809
rect 298787 145775 298816 145809
rect 298660 145744 298816 145775
rect 298660 145265 298816 145296
rect 298660 145231 298661 145265
rect 298695 145231 298753 145265
rect 298787 145231 298816 145265
rect 298660 145200 298816 145231
rect 298660 144721 298816 144752
rect 298660 144687 298661 144721
rect 298695 144687 298753 144721
rect 298787 144687 298816 144721
rect 298660 144656 298816 144687
rect 298660 144177 298816 144208
rect 298660 144143 298661 144177
rect 298695 144143 298753 144177
rect 298787 144143 298816 144177
rect 298660 144112 298816 144143
rect 298660 143633 298816 143664
rect 298660 143599 298661 143633
rect 298695 143599 298753 143633
rect 298787 143599 298816 143633
rect 298660 143568 298816 143599
rect 298660 143089 298816 143120
rect 298660 143055 298661 143089
rect 298695 143055 298753 143089
rect 298787 143055 298816 143089
rect 298660 143024 298816 143055
rect 298660 142545 298816 142576
rect 298660 142511 298661 142545
rect 298695 142511 298753 142545
rect 298787 142511 298816 142545
rect 298660 142480 298816 142511
rect 298660 142001 298816 142032
rect 298660 141967 298661 142001
rect 298695 141967 298753 142001
rect 298787 141967 298816 142001
rect 298660 141936 298816 141967
rect 298660 141457 298816 141488
rect 298660 141423 298661 141457
rect 298695 141423 298753 141457
rect 298787 141423 298816 141457
rect 298660 141392 298816 141423
rect 298660 140913 298816 140944
rect 298660 140879 298661 140913
rect 298695 140879 298753 140913
rect 298787 140879 298816 140913
rect 298660 140848 298816 140879
rect 298660 140369 298816 140400
rect 298660 140335 298661 140369
rect 298695 140335 298753 140369
rect 298787 140335 298816 140369
rect 298660 140304 298816 140335
rect 298660 139825 298816 139856
rect 298660 139791 298661 139825
rect 298695 139791 298753 139825
rect 298787 139791 298816 139825
rect 298660 139760 298816 139791
rect 298660 139281 298816 139312
rect 298660 139247 298661 139281
rect 298695 139247 298753 139281
rect 298787 139247 298816 139281
rect 298660 139216 298816 139247
rect 298660 138737 298816 138768
rect 298660 138703 298661 138737
rect 298695 138703 298753 138737
rect 298787 138703 298816 138737
rect 298660 138672 298816 138703
rect 298660 138193 298816 138224
rect 298660 138159 298661 138193
rect 298695 138159 298753 138193
rect 298787 138159 298816 138193
rect 298660 138128 298816 138159
rect 298660 137649 298816 137680
rect 298660 137615 298661 137649
rect 298695 137615 298753 137649
rect 298787 137615 298816 137649
rect 298660 137584 298816 137615
rect 298660 137105 298816 137136
rect 298660 137071 298661 137105
rect 298695 137071 298753 137105
rect 298787 137071 298816 137105
rect 298660 137040 298816 137071
rect 298660 136561 298816 136592
rect 298660 136527 298661 136561
rect 298695 136527 298753 136561
rect 298787 136527 298816 136561
rect 298660 136496 298816 136527
rect 298660 136017 298816 136048
rect 298660 135983 298661 136017
rect 298695 135983 298753 136017
rect 298787 135983 298816 136017
rect 298660 135952 298816 135983
rect 298660 135473 298816 135504
rect 298660 135439 298661 135473
rect 298695 135439 298753 135473
rect 298787 135439 298816 135473
rect 298660 135408 298816 135439
rect 298660 134929 298816 134960
rect 298660 134895 298661 134929
rect 298695 134895 298753 134929
rect 298787 134895 298816 134929
rect 298660 134864 298816 134895
rect 298660 134385 298816 134416
rect 298660 134351 298661 134385
rect 298695 134351 298753 134385
rect 298787 134351 298816 134385
rect 298660 134320 298816 134351
rect 298660 133841 298816 133872
rect 298660 133807 298661 133841
rect 298695 133807 298753 133841
rect 298787 133807 298816 133841
rect 298660 133776 298816 133807
rect 298660 133297 298816 133328
rect 298660 133263 298661 133297
rect 298695 133263 298753 133297
rect 298787 133263 298816 133297
rect 298660 133232 298816 133263
rect 298660 132753 298816 132784
rect 298660 132719 298661 132753
rect 298695 132719 298753 132753
rect 298787 132719 298816 132753
rect 298660 132688 298816 132719
rect 298660 132209 298816 132240
rect 298660 132175 298661 132209
rect 298695 132175 298753 132209
rect 298787 132175 298816 132209
rect 298660 132144 298816 132175
rect 298660 131665 298816 131696
rect 298660 131631 298661 131665
rect 298695 131631 298753 131665
rect 298787 131631 298816 131665
rect 298660 131600 298816 131631
rect 298660 131121 298816 131152
rect 298660 131087 298661 131121
rect 298695 131087 298753 131121
rect 298787 131087 298816 131121
rect 298660 131056 298816 131087
rect 298660 130577 298816 130608
rect 298660 130543 298661 130577
rect 298695 130543 298753 130577
rect 298787 130543 298816 130577
rect 298660 130512 298816 130543
rect 298660 130033 298816 130064
rect 298660 129999 298661 130033
rect 298695 129999 298753 130033
rect 298787 129999 298816 130033
rect 298660 129968 298816 129999
rect 298660 129489 298816 129520
rect 298660 129455 298661 129489
rect 298695 129455 298753 129489
rect 298787 129455 298816 129489
rect 298660 129424 298816 129455
rect 298660 128945 298816 128976
rect 298660 128911 298661 128945
rect 298695 128911 298753 128945
rect 298787 128911 298816 128945
rect 298660 128880 298816 128911
rect 298660 128401 298816 128432
rect 298660 128367 298661 128401
rect 298695 128367 298753 128401
rect 298787 128367 298816 128401
rect 298660 128336 298816 128367
rect 298660 127857 298816 127888
rect 298660 127823 298661 127857
rect 298695 127823 298753 127857
rect 298787 127823 298816 127857
rect 298660 127792 298816 127823
rect 298660 127313 298816 127344
rect 298660 127279 298661 127313
rect 298695 127279 298753 127313
rect 298787 127279 298816 127313
rect 298660 127248 298816 127279
rect 298660 126769 298816 126800
rect 298660 126735 298661 126769
rect 298695 126735 298753 126769
rect 298787 126735 298816 126769
rect 298660 126704 298816 126735
rect 298660 126225 298816 126256
rect 298660 126191 298661 126225
rect 298695 126191 298753 126225
rect 298787 126191 298816 126225
rect 298660 126160 298816 126191
rect 298660 125681 298816 125712
rect 298660 125647 298661 125681
rect 298695 125647 298753 125681
rect 298787 125647 298816 125681
rect 298660 125616 298816 125647
rect 298660 125137 298816 125168
rect 298660 125103 298661 125137
rect 298695 125103 298753 125137
rect 298787 125103 298816 125137
rect 298660 125072 298816 125103
rect 298660 124593 298816 124624
rect 298660 124559 298661 124593
rect 298695 124559 298753 124593
rect 298787 124559 298816 124593
rect 298660 124528 298816 124559
rect 298660 124049 298816 124080
rect 298660 124015 298661 124049
rect 298695 124015 298753 124049
rect 298787 124015 298816 124049
rect 298660 123984 298816 124015
rect 298660 123505 298816 123536
rect 298660 123471 298661 123505
rect 298695 123471 298753 123505
rect 298787 123471 298816 123505
rect 298660 123440 298816 123471
rect 298660 122961 298816 122992
rect 298660 122927 298661 122961
rect 298695 122927 298753 122961
rect 298787 122927 298816 122961
rect 298660 122896 298816 122927
rect 298660 122417 298816 122448
rect 298660 122383 298661 122417
rect 298695 122383 298753 122417
rect 298787 122383 298816 122417
rect 298660 122352 298816 122383
rect 298660 121873 298816 121904
rect 298660 121839 298661 121873
rect 298695 121839 298753 121873
rect 298787 121839 298816 121873
rect 298660 121808 298816 121839
rect 298660 121329 298816 121360
rect 298660 121295 298661 121329
rect 298695 121295 298753 121329
rect 298787 121295 298816 121329
rect 298660 121264 298816 121295
rect 298660 120785 298816 120816
rect 298660 120751 298661 120785
rect 298695 120751 298753 120785
rect 298787 120751 298816 120785
rect 298660 120720 298816 120751
rect 298660 120241 298816 120272
rect 298660 120207 298661 120241
rect 298695 120207 298753 120241
rect 298787 120207 298816 120241
rect 298660 120176 298816 120207
rect 298660 119697 298816 119728
rect 298660 119663 298661 119697
rect 298695 119663 298753 119697
rect 298787 119663 298816 119697
rect 298660 119632 298816 119663
rect 298660 119153 298816 119184
rect 298660 119119 298661 119153
rect 298695 119119 298753 119153
rect 298787 119119 298816 119153
rect 298660 119088 298816 119119
rect 298660 118609 298816 118640
rect 298660 118575 298661 118609
rect 298695 118575 298753 118609
rect 298787 118575 298816 118609
rect 298660 118544 298816 118575
rect 298660 118065 298816 118096
rect 298660 118031 298661 118065
rect 298695 118031 298753 118065
rect 298787 118031 298816 118065
rect 298660 118000 298816 118031
rect 298660 117521 298816 117552
rect 298660 117487 298661 117521
rect 298695 117487 298753 117521
rect 298787 117487 298816 117521
rect 298660 117456 298816 117487
rect 298660 116977 298816 117008
rect 298660 116943 298661 116977
rect 298695 116943 298753 116977
rect 298787 116943 298816 116977
rect 298660 116912 298816 116943
rect 298660 116433 298816 116464
rect 298660 116399 298661 116433
rect 298695 116399 298753 116433
rect 298787 116399 298816 116433
rect 298660 116368 298816 116399
rect 298660 115889 298816 115920
rect 298660 115855 298661 115889
rect 298695 115855 298753 115889
rect 298787 115855 298816 115889
rect 298660 115824 298816 115855
rect 298660 115345 298816 115376
rect 298660 115311 298661 115345
rect 298695 115311 298753 115345
rect 298787 115311 298816 115345
rect 298660 115280 298816 115311
rect 298660 114801 298816 114832
rect 298660 114767 298661 114801
rect 298695 114767 298753 114801
rect 298787 114767 298816 114801
rect 298660 114736 298816 114767
rect 298660 114257 298816 114288
rect 298660 114223 298661 114257
rect 298695 114223 298753 114257
rect 298787 114223 298816 114257
rect 298660 114192 298816 114223
rect 298660 113713 298816 113744
rect 298660 113679 298661 113713
rect 298695 113679 298753 113713
rect 298787 113679 298816 113713
rect 298660 113648 298816 113679
rect 298660 113169 298816 113200
rect 298660 113135 298661 113169
rect 298695 113135 298753 113169
rect 298787 113135 298816 113169
rect 298660 113104 298816 113135
rect 298660 112625 298816 112656
rect 298660 112591 298661 112625
rect 298695 112591 298753 112625
rect 298787 112591 298816 112625
rect 298660 112560 298816 112591
rect 298660 112081 298816 112112
rect 298660 112047 298661 112081
rect 298695 112047 298753 112081
rect 298787 112047 298816 112081
rect 298660 112016 298816 112047
rect 298660 111537 298816 111568
rect 298660 111503 298661 111537
rect 298695 111503 298753 111537
rect 298787 111503 298816 111537
rect 298660 111472 298816 111503
rect 298660 110993 298816 111024
rect 298660 110959 298661 110993
rect 298695 110959 298753 110993
rect 298787 110959 298816 110993
rect 298660 110928 298816 110959
rect 298660 110449 298816 110480
rect 298660 110415 298661 110449
rect 298695 110415 298753 110449
rect 298787 110415 298816 110449
rect 298660 110384 298816 110415
rect 298660 109905 298816 109936
rect 298660 109871 298661 109905
rect 298695 109871 298753 109905
rect 298787 109871 298816 109905
rect 298660 109840 298816 109871
rect 298660 109361 298816 109392
rect 298660 109327 298661 109361
rect 298695 109327 298753 109361
rect 298787 109327 298816 109361
rect 298660 109296 298816 109327
rect 298660 108817 298816 108848
rect 298660 108783 298661 108817
rect 298695 108783 298753 108817
rect 298787 108783 298816 108817
rect 298660 108752 298816 108783
rect 298660 108273 298816 108304
rect 298660 108239 298661 108273
rect 298695 108239 298753 108273
rect 298787 108239 298816 108273
rect 298660 108208 298816 108239
rect 298660 107729 298816 107760
rect 298660 107695 298661 107729
rect 298695 107695 298753 107729
rect 298787 107695 298816 107729
rect 298660 107664 298816 107695
rect 298660 107185 298816 107216
rect 298660 107151 298661 107185
rect 298695 107151 298753 107185
rect 298787 107151 298816 107185
rect 298660 107120 298816 107151
rect 298660 106641 298816 106672
rect 298660 106607 298661 106641
rect 298695 106607 298753 106641
rect 298787 106607 298816 106641
rect 298660 106576 298816 106607
rect 298660 106097 298816 106128
rect 298660 106063 298661 106097
rect 298695 106063 298753 106097
rect 298787 106063 298816 106097
rect 298660 106032 298816 106063
rect 298660 105553 298816 105584
rect 298660 105519 298661 105553
rect 298695 105519 298753 105553
rect 298787 105519 298816 105553
rect 298660 105488 298816 105519
rect 298660 105009 298816 105040
rect 298660 104975 298661 105009
rect 298695 104975 298753 105009
rect 298787 104975 298816 105009
rect 298660 104944 298816 104975
rect 298660 104465 298816 104496
rect 298660 104431 298661 104465
rect 298695 104431 298753 104465
rect 298787 104431 298816 104465
rect 298660 104400 298816 104431
rect 298660 103921 298816 103952
rect 298660 103887 298661 103921
rect 298695 103887 298753 103921
rect 298787 103887 298816 103921
rect 298660 103856 298816 103887
rect 298660 103377 298816 103408
rect 298660 103343 298661 103377
rect 298695 103343 298753 103377
rect 298787 103343 298816 103377
rect 298660 103312 298816 103343
rect 298660 102833 298816 102864
rect 298660 102799 298661 102833
rect 298695 102799 298753 102833
rect 298787 102799 298816 102833
rect 298660 102768 298816 102799
rect 298660 102289 298816 102320
rect 298660 102255 298661 102289
rect 298695 102255 298753 102289
rect 298787 102255 298816 102289
rect 298660 102224 298816 102255
rect 298660 101745 298816 101776
rect 298660 101711 298661 101745
rect 298695 101711 298753 101745
rect 298787 101711 298816 101745
rect 298660 101680 298816 101711
rect 298660 101201 298816 101232
rect 298660 101167 298661 101201
rect 298695 101167 298753 101201
rect 298787 101167 298816 101201
rect 298660 101136 298816 101167
rect 298660 100657 298816 100688
rect 298660 100623 298661 100657
rect 298695 100623 298753 100657
rect 298787 100623 298816 100657
rect 298660 100592 298816 100623
rect 298660 100113 298816 100144
rect 298660 100079 298661 100113
rect 298695 100079 298753 100113
rect 298787 100079 298816 100113
rect 298660 100048 298816 100079
rect 298660 99569 298816 99600
rect 298660 99535 298661 99569
rect 298695 99535 298753 99569
rect 298787 99535 298816 99569
rect 298660 99504 298816 99535
rect 298660 99025 298816 99056
rect 298660 98991 298661 99025
rect 298695 98991 298753 99025
rect 298787 98991 298816 99025
rect 298660 98960 298816 98991
rect 298660 98481 298816 98512
rect 298660 98447 298661 98481
rect 298695 98447 298753 98481
rect 298787 98447 298816 98481
rect 298660 98416 298816 98447
rect 298660 97937 298816 97968
rect 298660 97903 298661 97937
rect 298695 97903 298753 97937
rect 298787 97903 298816 97937
rect 298660 97872 298816 97903
rect 298660 97393 298816 97424
rect 298660 97359 298661 97393
rect 298695 97359 298753 97393
rect 298787 97359 298816 97393
rect 298660 97328 298816 97359
rect 298660 96849 298816 96880
rect 298660 96815 298661 96849
rect 298695 96815 298753 96849
rect 298787 96815 298816 96849
rect 298660 96784 298816 96815
rect 298660 96305 298816 96336
rect 298660 96271 298661 96305
rect 298695 96271 298753 96305
rect 298787 96271 298816 96305
rect 298660 96240 298816 96271
rect 298660 95761 298816 95792
rect 298660 95727 298661 95761
rect 298695 95727 298753 95761
rect 298787 95727 298816 95761
rect 298660 95696 298816 95727
rect 298660 95217 298816 95248
rect 298660 95183 298661 95217
rect 298695 95183 298753 95217
rect 298787 95183 298816 95217
rect 298660 95152 298816 95183
rect 298660 94673 298816 94704
rect 298660 94639 298661 94673
rect 298695 94639 298753 94673
rect 298787 94639 298816 94673
rect 298660 94608 298816 94639
rect 298660 94129 298816 94160
rect 298660 94095 298661 94129
rect 298695 94095 298753 94129
rect 298787 94095 298816 94129
rect 298660 94064 298816 94095
rect 298660 93585 298816 93616
rect 298660 93551 298661 93585
rect 298695 93551 298753 93585
rect 298787 93551 298816 93585
rect 298660 93520 298816 93551
rect 298660 93041 298816 93072
rect 298660 93007 298661 93041
rect 298695 93007 298753 93041
rect 298787 93007 298816 93041
rect 298660 92976 298816 93007
rect 298660 92497 298816 92528
rect 298660 92463 298661 92497
rect 298695 92463 298753 92497
rect 298787 92463 298816 92497
rect 298660 92432 298816 92463
rect 298660 91953 298816 91984
rect 298660 91919 298661 91953
rect 298695 91919 298753 91953
rect 298787 91919 298816 91953
rect 298660 91888 298816 91919
rect 298660 91409 298816 91440
rect 298660 91375 298661 91409
rect 298695 91375 298753 91409
rect 298787 91375 298816 91409
rect 298660 91344 298816 91375
rect 298660 90865 298816 90896
rect 298660 90831 298661 90865
rect 298695 90831 298753 90865
rect 298787 90831 298816 90865
rect 298660 90800 298816 90831
rect 298660 90321 298816 90352
rect 298660 90287 298661 90321
rect 298695 90287 298753 90321
rect 298787 90287 298816 90321
rect 298660 90256 298816 90287
rect 298660 89777 298816 89808
rect 298660 89743 298661 89777
rect 298695 89743 298753 89777
rect 298787 89743 298816 89777
rect 298660 89712 298816 89743
rect 298660 89233 298816 89264
rect 298660 89199 298661 89233
rect 298695 89199 298753 89233
rect 298787 89199 298816 89233
rect 298660 89168 298816 89199
rect 298660 88689 298816 88720
rect 298660 88655 298661 88689
rect 298695 88655 298753 88689
rect 298787 88655 298816 88689
rect 298660 88624 298816 88655
rect 298660 88145 298816 88176
rect 298660 88111 298661 88145
rect 298695 88111 298753 88145
rect 298787 88111 298816 88145
rect 298660 88080 298816 88111
rect 298660 87601 298816 87632
rect 298660 87567 298661 87601
rect 298695 87567 298753 87601
rect 298787 87567 298816 87601
rect 298660 87536 298816 87567
rect 298660 87057 298816 87088
rect 298660 87023 298661 87057
rect 298695 87023 298753 87057
rect 298787 87023 298816 87057
rect 298660 86992 298816 87023
rect 298660 86513 298816 86544
rect 298660 86479 298661 86513
rect 298695 86479 298753 86513
rect 298787 86479 298816 86513
rect 298660 86448 298816 86479
rect 298660 85969 298816 86000
rect 298660 85935 298661 85969
rect 298695 85935 298753 85969
rect 298787 85935 298816 85969
rect 298660 85904 298816 85935
rect 298660 85425 298816 85456
rect 298660 85391 298661 85425
rect 298695 85391 298753 85425
rect 298787 85391 298816 85425
rect 298660 85360 298816 85391
rect 298660 84881 298816 84912
rect 298660 84847 298661 84881
rect 298695 84847 298753 84881
rect 298787 84847 298816 84881
rect 298660 84816 298816 84847
rect 298660 84337 298816 84368
rect 298660 84303 298661 84337
rect 298695 84303 298753 84337
rect 298787 84303 298816 84337
rect 298660 84272 298816 84303
rect 298660 83793 298816 83824
rect 298660 83759 298661 83793
rect 298695 83759 298753 83793
rect 298787 83759 298816 83793
rect 298660 83728 298816 83759
rect 298660 83249 298816 83280
rect 298660 83215 298661 83249
rect 298695 83215 298753 83249
rect 298787 83215 298816 83249
rect 298660 83184 298816 83215
rect 298660 82705 298816 82736
rect 298660 82671 298661 82705
rect 298695 82671 298753 82705
rect 298787 82671 298816 82705
rect 298660 82640 298816 82671
rect 298660 82161 298816 82192
rect 298660 82127 298661 82161
rect 298695 82127 298753 82161
rect 298787 82127 298816 82161
rect 298660 82096 298816 82127
rect 298660 81617 298816 81648
rect 298660 81583 298661 81617
rect 298695 81583 298753 81617
rect 298787 81583 298816 81617
rect 298660 81552 298816 81583
rect 298660 81073 298816 81104
rect 298660 81039 298661 81073
rect 298695 81039 298753 81073
rect 298787 81039 298816 81073
rect 298660 81008 298816 81039
rect 298660 80529 298816 80560
rect 298660 80495 298661 80529
rect 298695 80495 298753 80529
rect 298787 80495 298816 80529
rect 298660 80464 298816 80495
rect 298660 79985 298816 80016
rect 298660 79951 298661 79985
rect 298695 79951 298753 79985
rect 298787 79951 298816 79985
rect 298660 79920 298816 79951
rect 298660 79441 298816 79472
rect 298660 79407 298661 79441
rect 298695 79407 298753 79441
rect 298787 79407 298816 79441
rect 298660 79376 298816 79407
rect 298660 78897 298816 78928
rect 298660 78863 298661 78897
rect 298695 78863 298753 78897
rect 298787 78863 298816 78897
rect 298660 78832 298816 78863
rect 298660 78353 298816 78384
rect 298660 78319 298661 78353
rect 298695 78319 298753 78353
rect 298787 78319 298816 78353
rect 298660 78288 298816 78319
rect 298660 77809 298816 77840
rect 298660 77775 298661 77809
rect 298695 77775 298753 77809
rect 298787 77775 298816 77809
rect 298660 77744 298816 77775
rect 298660 77265 298816 77296
rect 298660 77231 298661 77265
rect 298695 77231 298753 77265
rect 298787 77231 298816 77265
rect 298660 77200 298816 77231
rect 298660 76721 298816 76752
rect 298660 76687 298661 76721
rect 298695 76687 298753 76721
rect 298787 76687 298816 76721
rect 298660 76656 298816 76687
rect 298660 76177 298816 76208
rect 298660 76143 298661 76177
rect 298695 76143 298753 76177
rect 298787 76143 298816 76177
rect 298660 76112 298816 76143
rect 298660 75633 298816 75664
rect 298660 75599 298661 75633
rect 298695 75599 298753 75633
rect 298787 75599 298816 75633
rect 298660 75568 298816 75599
rect 298660 75089 298816 75120
rect 298660 75055 298661 75089
rect 298695 75055 298753 75089
rect 298787 75055 298816 75089
rect 298660 75024 298816 75055
rect 298660 74545 298816 74576
rect 298660 74511 298661 74545
rect 298695 74511 298753 74545
rect 298787 74511 298816 74545
rect 298660 74480 298816 74511
rect 298660 74001 298816 74032
rect 298660 73967 298661 74001
rect 298695 73967 298753 74001
rect 298787 73967 298816 74001
rect 298660 73936 298816 73967
rect 298660 73457 298816 73488
rect 298660 73423 298661 73457
rect 298695 73423 298753 73457
rect 298787 73423 298816 73457
rect 298660 73392 298816 73423
rect 298660 72913 298816 72944
rect 298660 72879 298661 72913
rect 298695 72879 298753 72913
rect 298787 72879 298816 72913
rect 298660 72848 298816 72879
rect 298660 72369 298816 72400
rect 298660 72335 298661 72369
rect 298695 72335 298753 72369
rect 298787 72335 298816 72369
rect 298660 72304 298816 72335
rect 298660 71825 298816 71856
rect 298660 71791 298661 71825
rect 298695 71791 298753 71825
rect 298787 71791 298816 71825
rect 298660 71760 298816 71791
rect 298660 71281 298816 71312
rect 298660 71247 298661 71281
rect 298695 71247 298753 71281
rect 298787 71247 298816 71281
rect 298660 71216 298816 71247
rect 298660 70737 298816 70768
rect 298660 70703 298661 70737
rect 298695 70703 298753 70737
rect 298787 70703 298816 70737
rect 298660 70672 298816 70703
rect 298660 70193 298816 70224
rect 298660 70159 298661 70193
rect 298695 70159 298753 70193
rect 298787 70159 298816 70193
rect 298660 70128 298816 70159
rect 298660 69649 298816 69680
rect 298660 69615 298661 69649
rect 298695 69615 298753 69649
rect 298787 69615 298816 69649
rect 298660 69584 298816 69615
rect 298660 69105 298816 69136
rect 298660 69071 298661 69105
rect 298695 69071 298753 69105
rect 298787 69071 298816 69105
rect 298660 69040 298816 69071
rect 298660 68561 298816 68592
rect 298660 68527 298661 68561
rect 298695 68527 298753 68561
rect 298787 68527 298816 68561
rect 298660 68496 298816 68527
rect 298660 68017 298816 68048
rect 298660 67983 298661 68017
rect 298695 67983 298753 68017
rect 298787 67983 298816 68017
rect 298660 67952 298816 67983
rect 298660 67473 298816 67504
rect 298660 67439 298661 67473
rect 298695 67439 298753 67473
rect 298787 67439 298816 67473
rect 298660 67408 298816 67439
rect 298660 66929 298816 66960
rect 298660 66895 298661 66929
rect 298695 66895 298753 66929
rect 298787 66895 298816 66929
rect 298660 66864 298816 66895
rect 298660 66385 298816 66416
rect 298660 66351 298661 66385
rect 298695 66351 298753 66385
rect 298787 66351 298816 66385
rect 298660 66320 298816 66351
rect 298660 65841 298816 65872
rect 298660 65807 298661 65841
rect 298695 65807 298753 65841
rect 298787 65807 298816 65841
rect 298660 65776 298816 65807
rect 298660 65297 298816 65328
rect 298660 65263 298661 65297
rect 298695 65263 298753 65297
rect 298787 65263 298816 65297
rect 298660 65232 298816 65263
rect 298660 64753 298816 64784
rect 298660 64719 298661 64753
rect 298695 64719 298753 64753
rect 298787 64719 298816 64753
rect 298660 64688 298816 64719
rect 298660 64209 298816 64240
rect 298660 64175 298661 64209
rect 298695 64175 298753 64209
rect 298787 64175 298816 64209
rect 298660 64144 298816 64175
rect 298660 63665 298816 63696
rect 298660 63631 298661 63665
rect 298695 63631 298753 63665
rect 298787 63631 298816 63665
rect 298660 63600 298816 63631
rect 298660 63121 298816 63152
rect 298660 63087 298661 63121
rect 298695 63087 298753 63121
rect 298787 63087 298816 63121
rect 298660 63056 298816 63087
rect 298660 62577 298816 62608
rect 298660 62543 298661 62577
rect 298695 62543 298753 62577
rect 298787 62543 298816 62577
rect 298660 62512 298816 62543
rect 298660 62033 298816 62064
rect 298660 61999 298661 62033
rect 298695 61999 298753 62033
rect 298787 61999 298816 62033
rect 298660 61968 298816 61999
rect 298660 61489 298816 61520
rect 298660 61455 298661 61489
rect 298695 61455 298753 61489
rect 298787 61455 298816 61489
rect 298660 61424 298816 61455
rect 298660 60945 298816 60976
rect 298660 60911 298661 60945
rect 298695 60911 298753 60945
rect 298787 60911 298816 60945
rect 298660 60880 298816 60911
rect 298660 60401 298816 60432
rect 298660 60367 298661 60401
rect 298695 60367 298753 60401
rect 298787 60367 298816 60401
rect 298660 60336 298816 60367
rect 298660 59857 298816 59888
rect 298660 59823 298661 59857
rect 298695 59823 298753 59857
rect 298787 59823 298816 59857
rect 298660 59792 298816 59823
rect 298660 59313 298816 59344
rect 298660 59279 298661 59313
rect 298695 59279 298753 59313
rect 298787 59279 298816 59313
rect 298660 59248 298816 59279
rect 298660 58769 298816 58800
rect 298660 58735 298661 58769
rect 298695 58735 298753 58769
rect 298787 58735 298816 58769
rect 298660 58704 298816 58735
rect 298660 58225 298816 58256
rect 298660 58191 298661 58225
rect 298695 58191 298753 58225
rect 298787 58191 298816 58225
rect 298660 58160 298816 58191
rect 298660 57681 298816 57712
rect 298660 57647 298661 57681
rect 298695 57647 298753 57681
rect 298787 57647 298816 57681
rect 298660 57616 298816 57647
rect 298660 57137 298816 57168
rect 298660 57103 298661 57137
rect 298695 57103 298753 57137
rect 298787 57103 298816 57137
rect 298660 57072 298816 57103
rect 298660 56593 298816 56624
rect 298660 56559 298661 56593
rect 298695 56559 298753 56593
rect 298787 56559 298816 56593
rect 298660 56528 298816 56559
rect 298660 56049 298816 56080
rect 298660 56015 298661 56049
rect 298695 56015 298753 56049
rect 298787 56015 298816 56049
rect 298660 55984 298816 56015
rect 298660 55505 298816 55536
rect 298660 55471 298661 55505
rect 298695 55471 298753 55505
rect 298787 55471 298816 55505
rect 298660 55440 298816 55471
rect 298660 54961 298816 54992
rect 298660 54927 298661 54961
rect 298695 54927 298753 54961
rect 298787 54927 298816 54961
rect 298660 54896 298816 54927
rect 298660 54417 298816 54448
rect 298660 54383 298661 54417
rect 298695 54383 298753 54417
rect 298787 54383 298816 54417
rect 298660 54352 298816 54383
rect 298660 53873 298816 53904
rect 298660 53839 298661 53873
rect 298695 53839 298753 53873
rect 298787 53839 298816 53873
rect 298660 53808 298816 53839
rect 298660 53329 298816 53360
rect 298660 53295 298661 53329
rect 298695 53295 298753 53329
rect 298787 53295 298816 53329
rect 298660 53264 298816 53295
rect 298660 52785 298816 52816
rect 298660 52751 298661 52785
rect 298695 52751 298753 52785
rect 298787 52751 298816 52785
rect 298660 52720 298816 52751
rect 298660 52241 298816 52272
rect 298660 52207 298661 52241
rect 298695 52207 298753 52241
rect 298787 52207 298816 52241
rect 298660 52176 298816 52207
rect 298660 51697 298816 51728
rect 298660 51663 298661 51697
rect 298695 51663 298753 51697
rect 298787 51663 298816 51697
rect 298660 51632 298816 51663
rect 298660 51153 298816 51184
rect 298660 51119 298661 51153
rect 298695 51119 298753 51153
rect 298787 51119 298816 51153
rect 298660 51088 298816 51119
rect 298660 50609 298816 50640
rect 298660 50575 298661 50609
rect 298695 50575 298753 50609
rect 298787 50575 298816 50609
rect 298660 50544 298816 50575
rect 298660 50065 298816 50096
rect 298660 50031 298661 50065
rect 298695 50031 298753 50065
rect 298787 50031 298816 50065
rect 298660 50000 298816 50031
rect 298660 49521 298816 49552
rect 298660 49487 298661 49521
rect 298695 49487 298753 49521
rect 298787 49487 298816 49521
rect 298660 49456 298816 49487
rect 298660 48977 298816 49008
rect 298660 48943 298661 48977
rect 298695 48943 298753 48977
rect 298787 48943 298816 48977
rect 298660 48912 298816 48943
rect 298660 48433 298816 48464
rect 298660 48399 298661 48433
rect 298695 48399 298753 48433
rect 298787 48399 298816 48433
rect 298660 48368 298816 48399
rect 298660 47889 298816 47920
rect 298660 47855 298661 47889
rect 298695 47855 298753 47889
rect 298787 47855 298816 47889
rect 298660 47824 298816 47855
rect 298660 47345 298816 47376
rect 298660 47311 298661 47345
rect 298695 47311 298753 47345
rect 298787 47311 298816 47345
rect 298660 47280 298816 47311
rect 298660 46801 298816 46832
rect 298660 46767 298661 46801
rect 298695 46767 298753 46801
rect 298787 46767 298816 46801
rect 298660 46736 298816 46767
rect 298660 46257 298816 46288
rect 298660 46223 298661 46257
rect 298695 46223 298753 46257
rect 298787 46223 298816 46257
rect 298660 46192 298816 46223
rect 298660 45713 298816 45744
rect 298660 45679 298661 45713
rect 298695 45679 298753 45713
rect 298787 45679 298816 45713
rect 298660 45648 298816 45679
rect 298660 45169 298816 45200
rect 298660 45135 298661 45169
rect 298695 45135 298753 45169
rect 298787 45135 298816 45169
rect 298660 45104 298816 45135
rect 298660 44625 298816 44656
rect 298660 44591 298661 44625
rect 298695 44591 298753 44625
rect 298787 44591 298816 44625
rect 298660 44560 298816 44591
rect 298660 44081 298816 44112
rect 298660 44047 298661 44081
rect 298695 44047 298753 44081
rect 298787 44047 298816 44081
rect 298660 44016 298816 44047
rect 298660 43537 298816 43568
rect 298660 43503 298661 43537
rect 298695 43503 298753 43537
rect 298787 43503 298816 43537
rect 298660 43472 298816 43503
rect 298660 42993 298816 43024
rect 298660 42959 298661 42993
rect 298695 42959 298753 42993
rect 298787 42959 298816 42993
rect 298660 42928 298816 42959
rect 298660 42449 298816 42480
rect 298660 42415 298661 42449
rect 298695 42415 298753 42449
rect 298787 42415 298816 42449
rect 298660 42384 298816 42415
rect 298660 41905 298816 41936
rect 298660 41871 298661 41905
rect 298695 41871 298753 41905
rect 298787 41871 298816 41905
rect 298660 41840 298816 41871
rect 298660 41361 298816 41392
rect 298660 41327 298661 41361
rect 298695 41327 298753 41361
rect 298787 41327 298816 41361
rect 298660 41296 298816 41327
rect 298660 40817 298816 40848
rect 298660 40783 298661 40817
rect 298695 40783 298753 40817
rect 298787 40783 298816 40817
rect 298660 40752 298816 40783
rect 298660 40273 298816 40304
rect 298660 40239 298661 40273
rect 298695 40239 298753 40273
rect 298787 40239 298816 40273
rect 298660 40208 298816 40239
rect 298660 39729 298816 39760
rect 298660 39695 298661 39729
rect 298695 39695 298753 39729
rect 298787 39695 298816 39729
rect 298660 39664 298816 39695
rect 298660 39185 298816 39216
rect 298660 39151 298661 39185
rect 298695 39151 298753 39185
rect 298787 39151 298816 39185
rect 298660 39120 298816 39151
rect 298660 38641 298816 38672
rect 298660 38607 298661 38641
rect 298695 38607 298753 38641
rect 298787 38607 298816 38641
rect 298660 38576 298816 38607
rect 298660 38097 298816 38128
rect 298660 38063 298661 38097
rect 298695 38063 298753 38097
rect 298787 38063 298816 38097
rect 298660 38032 298816 38063
rect 298660 37553 298816 37584
rect 298660 37519 298661 37553
rect 298695 37519 298753 37553
rect 298787 37519 298816 37553
rect 298660 37488 298816 37519
rect 298660 37009 298816 37040
rect 298660 36975 298661 37009
rect 298695 36975 298753 37009
rect 298787 36975 298816 37009
rect 298660 36944 298816 36975
rect 298660 36465 298816 36496
rect 298660 36431 298661 36465
rect 298695 36431 298753 36465
rect 298787 36431 298816 36465
rect 298660 36400 298816 36431
rect 298660 35921 298816 35952
rect 298660 35887 298661 35921
rect 298695 35887 298753 35921
rect 298787 35887 298816 35921
rect 298660 35856 298816 35887
rect 298660 35377 298816 35408
rect 298660 35343 298661 35377
rect 298695 35343 298753 35377
rect 298787 35343 298816 35377
rect 298660 35312 298816 35343
rect 298660 34833 298816 34864
rect 298660 34799 298661 34833
rect 298695 34799 298753 34833
rect 298787 34799 298816 34833
rect 298660 34768 298816 34799
rect 298660 34289 298816 34320
rect 298660 34255 298661 34289
rect 298695 34255 298753 34289
rect 298787 34255 298816 34289
rect 298660 34224 298816 34255
rect 298660 33745 298816 33776
rect 298660 33711 298661 33745
rect 298695 33711 298753 33745
rect 298787 33711 298816 33745
rect 298660 33680 298816 33711
rect 298660 33201 298816 33232
rect 298660 33167 298661 33201
rect 298695 33167 298753 33201
rect 298787 33167 298816 33201
rect 298660 33136 298816 33167
rect 298660 32657 298816 32688
rect 298660 32623 298661 32657
rect 298695 32623 298753 32657
rect 298787 32623 298816 32657
rect 298660 32592 298816 32623
rect 298660 32113 298816 32144
rect 298660 32079 298661 32113
rect 298695 32079 298753 32113
rect 298787 32079 298816 32113
rect 298660 32048 298816 32079
rect 298660 31569 298816 31600
rect 298660 31535 298661 31569
rect 298695 31535 298753 31569
rect 298787 31535 298816 31569
rect 298660 31504 298816 31535
rect 298660 31025 298816 31056
rect 298660 30991 298661 31025
rect 298695 30991 298753 31025
rect 298787 30991 298816 31025
rect 298660 30960 298816 30991
rect 298660 30481 298816 30512
rect 298660 30447 298661 30481
rect 298695 30447 298753 30481
rect 298787 30447 298816 30481
rect 298660 30416 298816 30447
rect 298660 29937 298816 29968
rect 298660 29903 298661 29937
rect 298695 29903 298753 29937
rect 298787 29903 298816 29937
rect 298660 29872 298816 29903
rect 298660 29393 298816 29424
rect 298660 29359 298661 29393
rect 298695 29359 298753 29393
rect 298787 29359 298816 29393
rect 298660 29328 298816 29359
rect 298660 28849 298816 28880
rect 298660 28815 298661 28849
rect 298695 28815 298753 28849
rect 298787 28815 298816 28849
rect 298660 28784 298816 28815
rect 298660 28305 298816 28336
rect 298660 28271 298661 28305
rect 298695 28271 298753 28305
rect 298787 28271 298816 28305
rect 298660 28240 298816 28271
rect 298660 27761 298816 27792
rect 298660 27727 298661 27761
rect 298695 27727 298753 27761
rect 298787 27727 298816 27761
rect 298660 27696 298816 27727
rect 298660 27217 298816 27248
rect 298660 27183 298661 27217
rect 298695 27183 298753 27217
rect 298787 27183 298816 27217
rect 298660 27152 298816 27183
rect 298660 26673 298816 26704
rect 298660 26639 298661 26673
rect 298695 26639 298753 26673
rect 298787 26639 298816 26673
rect 298660 26608 298816 26639
rect 298660 26129 298816 26160
rect 298660 26095 298661 26129
rect 298695 26095 298753 26129
rect 298787 26095 298816 26129
rect 298660 26064 298816 26095
rect 298660 25585 298816 25616
rect 298660 25551 298661 25585
rect 298695 25551 298753 25585
rect 298787 25551 298816 25585
rect 298660 25520 298816 25551
rect 298660 25041 298816 25072
rect 298660 25007 298661 25041
rect 298695 25007 298753 25041
rect 298787 25007 298816 25041
rect 298660 24976 298816 25007
rect 298660 24497 298816 24528
rect 298660 24463 298661 24497
rect 298695 24463 298753 24497
rect 298787 24463 298816 24497
rect 298660 24432 298816 24463
rect 298660 23953 298816 23984
rect 298660 23919 298661 23953
rect 298695 23919 298753 23953
rect 298787 23919 298816 23953
rect 298660 23888 298816 23919
rect 298660 23409 298816 23440
rect 298660 23375 298661 23409
rect 298695 23375 298753 23409
rect 298787 23375 298816 23409
rect 298660 23344 298816 23375
rect 298660 22865 298816 22896
rect 298660 22831 298661 22865
rect 298695 22831 298753 22865
rect 298787 22831 298816 22865
rect 298660 22800 298816 22831
rect 298660 22321 298816 22352
rect 298660 22287 298661 22321
rect 298695 22287 298753 22321
rect 298787 22287 298816 22321
rect 298660 22256 298816 22287
rect 298660 21777 298816 21808
rect 298660 21743 298661 21777
rect 298695 21743 298753 21777
rect 298787 21743 298816 21777
rect 298660 21712 298816 21743
rect 298660 21233 298816 21264
rect 298660 21199 298661 21233
rect 298695 21199 298753 21233
rect 298787 21199 298816 21233
rect 298660 21168 298816 21199
rect 298660 20689 298816 20720
rect 298660 20655 298661 20689
rect 298695 20655 298753 20689
rect 298787 20655 298816 20689
rect 298660 20624 298816 20655
rect 298660 20145 298816 20176
rect 298660 20111 298661 20145
rect 298695 20111 298753 20145
rect 298787 20111 298816 20145
rect 298660 20080 298816 20111
rect 298660 19601 298816 19632
rect 298660 19567 298661 19601
rect 298695 19567 298753 19601
rect 298787 19567 298816 19601
rect 298660 19536 298816 19567
rect 298660 19057 298816 19088
rect 298660 19023 298661 19057
rect 298695 19023 298753 19057
rect 298787 19023 298816 19057
rect 298660 18992 298816 19023
rect 298660 18513 298816 18544
rect 298660 18479 298661 18513
rect 298695 18479 298753 18513
rect 298787 18479 298816 18513
rect 298660 18448 298816 18479
rect 298660 17969 298816 18000
rect 298660 17935 298661 17969
rect 298695 17935 298753 17969
rect 298787 17935 298816 17969
rect 298660 17904 298816 17935
rect 298660 17425 298816 17456
rect 298660 17391 298661 17425
rect 298695 17391 298753 17425
rect 298787 17391 298816 17425
rect 298660 17360 298816 17391
rect 298660 16881 298816 16912
rect 298660 16847 298661 16881
rect 298695 16847 298753 16881
rect 298787 16847 298816 16881
rect 298660 16816 298816 16847
rect 298660 16337 298816 16368
rect 298660 16303 298661 16337
rect 298695 16303 298753 16337
rect 298787 16303 298816 16337
rect 298660 16272 298816 16303
rect 298660 15793 298816 15824
rect 298660 15759 298661 15793
rect 298695 15759 298753 15793
rect 298787 15759 298816 15793
rect 298660 15728 298816 15759
rect 298660 15249 298816 15280
rect 298660 15215 298661 15249
rect 298695 15215 298753 15249
rect 298787 15215 298816 15249
rect 298660 15184 298816 15215
rect 298660 14705 298816 14736
rect 298660 14671 298661 14705
rect 298695 14671 298753 14705
rect 298787 14671 298816 14705
rect 298660 14640 298816 14671
rect 298660 14161 298816 14192
rect 298660 14127 298661 14161
rect 298695 14127 298753 14161
rect 298787 14127 298816 14161
rect 298660 14096 298816 14127
rect 298660 13617 298816 13648
rect 298660 13583 298661 13617
rect 298695 13583 298753 13617
rect 298787 13583 298816 13617
rect 298660 13552 298816 13583
rect 298660 13073 298816 13104
rect 298660 13039 298661 13073
rect 298695 13039 298753 13073
rect 298787 13039 298816 13073
rect 298660 13008 298816 13039
rect 298660 12529 298816 12560
rect 298660 12495 298661 12529
rect 298695 12495 298753 12529
rect 298787 12495 298816 12529
rect 298660 12464 298816 12495
rect 298660 11985 298816 12016
rect 298660 11951 298661 11985
rect 298695 11951 298753 11985
rect 298787 11951 298816 11985
rect 298660 11920 298816 11951
rect 298660 11441 298816 11472
rect 298660 11407 298661 11441
rect 298695 11407 298753 11441
rect 298787 11407 298816 11441
rect 298660 11376 298816 11407
rect 298660 10897 298816 10928
rect 298660 10863 298661 10897
rect 298695 10863 298753 10897
rect 298787 10863 298816 10897
rect 298660 10832 298816 10863
rect 298660 10353 298816 10384
rect 298660 10319 298661 10353
rect 298695 10319 298753 10353
rect 298787 10319 298816 10353
rect 298660 10288 298816 10319
rect 298660 9809 298816 9840
rect 298660 9775 298661 9809
rect 298695 9775 298753 9809
rect 298787 9775 298816 9809
rect 298660 9744 298816 9775
rect 298660 9265 298816 9296
rect 298660 9231 298661 9265
rect 298695 9231 298753 9265
rect 298787 9231 298816 9265
rect 298660 9200 298816 9231
rect 298660 8721 298816 8752
rect 298660 8687 298661 8721
rect 298695 8687 298753 8721
rect 298787 8687 298816 8721
rect 298660 8656 298816 8687
rect 298660 8177 298816 8208
rect 298660 8143 298661 8177
rect 298695 8143 298753 8177
rect 298787 8143 298816 8177
rect 298660 8112 298816 8143
rect 298660 7633 298816 7664
rect 298660 7599 298661 7633
rect 298695 7599 298753 7633
rect 298787 7599 298816 7633
rect 298660 7568 298816 7599
rect 298660 7089 298816 7120
rect 298660 7055 298661 7089
rect 298695 7055 298753 7089
rect 298787 7055 298816 7089
rect 298660 7024 298816 7055
rect 298660 6545 298816 6576
rect 298660 6511 298661 6545
rect 298695 6511 298753 6545
rect 298787 6511 298816 6545
rect 298660 6480 298816 6511
rect 298660 6001 298816 6032
rect 298660 5967 298661 6001
rect 298695 5967 298753 6001
rect 298787 5967 298816 6001
rect 298660 5936 298816 5967
rect 298660 5457 298816 5488
rect 298660 5423 298661 5457
rect 298695 5423 298753 5457
rect 298787 5423 298816 5457
rect 298660 5392 298816 5423
rect 298660 4913 298816 4944
rect 298660 4879 298661 4913
rect 298695 4879 298753 4913
rect 298787 4879 298816 4913
rect 298660 4848 298816 4879
rect 298660 4369 298816 4400
rect 298660 4335 298661 4369
rect 298695 4335 298753 4369
rect 298787 4335 298816 4369
rect 298660 4304 298816 4335
rect 298660 3825 298816 3856
rect 298660 3791 298661 3825
rect 298695 3791 298753 3825
rect 298787 3791 298816 3825
rect 298660 3760 298816 3791
rect 298660 3281 298816 3312
rect 298660 3247 298661 3281
rect 298695 3247 298753 3281
rect 298787 3247 298816 3281
rect 298660 3216 298816 3247
rect 298660 2737 298816 2768
rect 298660 2703 298661 2737
rect 298695 2703 298753 2737
rect 298787 2703 298816 2737
rect 298660 2672 298816 2703
rect 298660 2193 298816 2224
rect 298660 2159 298661 2193
rect 298695 2159 298753 2193
rect 298787 2159 298816 2193
rect 298660 2128 298816 2159
<< via1 >>
rect 296 4088 348 4140
rect 848 3408 900 3460
<< obsm1 >>
rect 1340 2128 298660 297616
<< metal2 >>
rect 1278 299400 1390 301200
rect 3854 299400 3966 301200
rect 6430 299400 6542 301200
rect 9098 299400 9210 301200
rect 11674 299400 11786 301200
rect 14250 299400 14362 301200
rect 16918 299400 17030 301200
rect 19494 299400 19606 301200
rect 22070 299400 22182 301200
rect 24738 299400 24850 301200
rect 27314 299400 27426 301200
rect 29890 299400 30002 301200
rect 32558 299400 32670 301200
rect 35134 299400 35246 301200
rect 37710 299400 37822 301200
rect 40378 299400 40490 301200
rect 42954 299400 43066 301200
rect 45622 299400 45734 301200
rect 48198 299400 48310 301200
rect 50774 299400 50886 301200
rect 53442 299400 53554 301200
rect 56018 299400 56130 301200
rect 58594 299400 58706 301200
rect 61262 299400 61374 301200
rect 63838 299400 63950 301200
rect 66414 299400 66526 301200
rect 69082 299400 69194 301200
rect 71658 299400 71770 301200
rect 74234 299400 74346 301200
rect 76902 299400 77014 301200
rect 79478 299400 79590 301200
rect 82146 299400 82258 301200
rect 84722 299400 84834 301200
rect 87298 299400 87410 301200
rect 89966 299400 90078 301200
rect 92542 299400 92654 301200
rect 95118 299400 95230 301200
rect 97786 299400 97898 301200
rect 100362 299400 100474 301200
rect 102938 299400 103050 301200
rect 105606 299400 105718 301200
rect 108182 299400 108294 301200
rect 110758 299400 110870 301200
rect 113426 299400 113538 301200
rect 116002 299400 116114 301200
rect 118670 299400 118782 301200
rect 121246 299400 121358 301200
rect 123822 299400 123934 301200
rect 126490 299400 126602 301200
rect 129066 299400 129178 301200
rect 131642 299400 131754 301200
rect 134310 299400 134422 301200
rect 136886 299400 136998 301200
rect 139462 299400 139574 301200
rect 142130 299400 142242 301200
rect 144706 299400 144818 301200
rect 147282 299400 147394 301200
rect 149950 299400 150062 301200
rect 152526 299400 152638 301200
rect 155194 299400 155306 301200
rect 157770 299400 157882 301200
rect 160346 299400 160458 301200
rect 163014 299400 163126 301200
rect 165590 299400 165702 301200
rect 168166 299400 168278 301200
rect 170834 299400 170946 301200
rect 173410 299400 173522 301200
rect 175986 299400 176098 301200
rect 178654 299400 178766 301200
rect 181230 299400 181342 301200
rect 183806 299400 183918 301200
rect 186474 299400 186586 301200
rect 189050 299400 189162 301200
rect 191718 299400 191830 301200
rect 194294 299400 194406 301200
rect 196870 299400 196982 301200
rect 199538 299400 199650 301200
rect 202114 299400 202226 301200
rect 204690 299400 204802 301200
rect 207358 299400 207470 301200
rect 209934 299400 210046 301200
rect 212510 299400 212622 301200
rect 215178 299400 215290 301200
rect 217754 299400 217866 301200
rect 220330 299400 220442 301200
rect 222998 299400 223110 301200
rect 225574 299400 225686 301200
rect 228242 299400 228354 301200
rect 230818 299400 230930 301200
rect 233394 299400 233506 301200
rect 236062 299400 236174 301200
rect 238638 299400 238750 301200
rect 241214 299400 241326 301200
rect 243882 299400 243994 301200
rect 246458 299400 246570 301200
rect 249034 299400 249146 301200
rect 251702 299400 251814 301200
rect 254278 299400 254390 301200
rect 256854 299400 256966 301200
rect 259522 299400 259634 301200
rect 262098 299400 262210 301200
rect 264766 299400 264878 301200
rect 267342 299400 267454 301200
rect 269918 299400 270030 301200
rect 272586 299400 272698 301200
rect 275162 299400 275274 301200
rect 277738 299400 277850 301200
rect 280406 299400 280518 301200
rect 282982 299400 283094 301200
rect 285558 299400 285670 301200
rect 288226 299400 288338 301200
rect 290802 299400 290914 301200
rect 293378 299400 293490 301200
rect 296046 299400 296158 301200
rect 298622 299400 298734 301200
rect 3896 298660 3924 299400
rect 6472 298660 6500 299400
rect 11716 298660 11744 299400
rect 14292 298660 14320 299400
rect 19536 298660 19564 299400
rect 22112 298660 22140 299400
rect 27356 298660 27384 299400
rect 29932 298660 29960 299400
rect 35176 298660 35204 299400
rect 37752 298660 37780 299400
rect 42996 298660 43024 299400
rect 45664 298660 45692 299400
rect 50816 298660 50844 299400
rect 53484 298660 53512 299400
rect 58636 298660 58664 299400
rect 61304 298660 61332 299400
rect 66456 298660 66484 299400
rect 69124 298660 69152 299400
rect 74276 298660 74304 299400
rect 76944 298660 76972 299400
rect 82188 298660 82216 299400
rect 84764 298660 84792 299400
rect 90008 298660 90036 299400
rect 92584 298660 92612 299400
rect 97828 298660 97856 299400
rect 100404 298660 100432 299400
rect 105648 298660 105676 299400
rect 108224 298660 108252 299400
rect 113468 298660 113496 299400
rect 116044 298660 116072 299400
rect 121288 298660 121316 299400
rect 123864 298660 123892 299400
rect 129108 298660 129136 299400
rect 131684 298660 131712 299400
rect 136928 298660 136956 299400
rect 139504 298660 139532 299400
rect 144748 298660 144776 299400
rect 147324 298660 147352 299400
rect 152568 298660 152596 299400
rect 155236 298660 155264 299400
rect 160388 298660 160416 299400
rect 163056 298660 163084 299400
rect 168208 298660 168236 299400
rect 170876 298660 170904 299400
rect 176028 298660 176056 299400
rect 178696 298660 178724 299400
rect 183848 298660 183876 299400
rect 186516 298660 186544 299400
rect 191760 298660 191788 299400
rect 194336 298660 194364 299400
rect 199580 298660 199608 299400
rect 202156 298660 202184 299400
rect 207400 298660 207428 299400
rect 209976 298660 210004 299400
rect 215220 298660 215248 299400
rect 217796 298660 217824 299400
rect 223040 298660 223068 299400
rect 225616 298660 225644 299400
rect 230860 298660 230888 299400
rect 233436 298660 233464 299400
rect 238680 298660 238708 299400
rect 241256 298660 241284 299400
rect 246500 298660 246528 299400
rect 249076 298660 249104 299400
rect 254320 298660 254348 299400
rect 256896 298660 256924 299400
rect 262140 298660 262168 299400
rect 264808 298660 264836 299400
rect 269960 298660 269988 299400
rect 272628 298660 272656 299400
rect 277780 298660 277808 299400
rect 280448 298660 280476 299400
rect 285600 298660 285628 299400
rect 288268 298660 288296 299400
rect 293420 298660 293448 299400
rect 296088 298660 296116 299400
rect 296 4140 348 4146
rect 296 4082 348 4088
rect 308 600 336 4082
rect 848 3460 900 3466
rect 848 3402 900 3408
rect 860 600 888 3402
rect 1504 600 1532 1340
rect 2056 600 2084 1340
rect 2700 600 2728 1340
rect 3344 600 3372 1340
rect 4540 600 4568 1340
rect 5184 600 5212 1340
rect 5736 600 5764 1340
rect 6932 600 6960 1340
rect 7576 600 7604 1340
rect 8220 600 8248 1340
rect 9416 600 9444 1340
rect 10060 600 10088 1340
rect 10612 600 10640 1340
rect 11808 600 11836 1340
rect 12452 600 12480 1340
rect 13096 600 13124 1340
rect 14292 600 14320 1340
rect 14936 600 14964 1340
rect 16132 600 16160 1340
rect 16684 600 16712 1340
rect 17972 600 18000 1340
rect 18524 600 18552 1340
rect 19812 600 19840 1340
rect 20364 600 20392 1340
rect 21560 600 21588 1340
rect 22204 600 22232 1340
rect 23400 600 23428 1340
rect 24044 600 24072 1340
rect 25240 600 25268 1340
rect 25884 600 25912 1340
rect 27080 600 27108 1340
rect 27724 600 27752 1340
rect 28920 600 28948 1340
rect 29564 600 29592 1340
rect 30760 600 30788 1340
rect 31404 600 31432 1340
rect 32600 600 32628 1340
rect 33152 600 33180 1340
rect 34440 600 34468 1340
rect 34992 600 35020 1340
rect 36280 600 36308 1340
rect 36832 600 36860 1340
rect 38028 600 38056 1340
rect 38672 600 38700 1340
rect 39868 600 39896 1340
rect 40512 600 40540 1340
rect 41800 626 41828 1340
rect 41708 600 41828 626
rect 42352 600 42380 1340
rect 43548 600 43576 1340
rect 44192 600 44220 1340
rect 45388 600 45416 1340
rect 46032 600 46060 1340
rect 47228 600 47256 1340
rect 47780 600 47808 1340
rect 49068 600 49096 1340
rect 49620 600 49648 1340
rect 50908 600 50936 1340
rect 51368 626 51396 1340
rect 51368 600 51488 626
rect 52748 600 52776 1340
rect 53300 600 53328 1340
rect 54312 626 54340 1340
rect 55232 626 55260 1340
rect 54312 600 54524 626
rect 55140 600 55260 626
rect 56152 626 56180 1340
rect 56152 600 56364 626
rect 56980 600 57008 1340
rect 58176 600 58204 1340
rect 58820 600 58848 1340
rect 60108 626 60136 1340
rect 60016 600 60136 626
rect 60660 600 60688 1340
rect 61856 600 61884 1340
rect 62500 600 62528 1340
rect 63696 600 63724 1340
rect 64248 600 64276 1340
rect 65536 600 65564 1340
rect 67376 600 67404 1340
rect 69124 600 69152 1340
rect 70964 600 70992 1340
rect 72804 600 72832 1340
rect 74644 600 74672 1340
rect 76484 600 76512 1340
rect 78600 626 78628 1340
rect 78324 600 78628 626
rect 80164 600 80192 1340
rect 82004 600 82032 1340
rect 84120 626 84148 1340
rect 83844 600 84148 626
rect 85592 600 85620 1340
rect 87432 600 87460 1340
rect 89272 600 89300 1340
rect 91112 600 91140 1340
rect 92952 600 92980 1340
rect 94792 600 94820 1340
rect 96632 600 96660 1340
rect 98472 600 98500 1340
rect 100680 626 100708 1340
rect 100312 600 100708 626
rect 102060 600 102088 1340
rect 103900 600 103928 1340
rect 105740 600 105768 1340
rect 107580 600 107608 1340
rect 109420 600 109448 1340
rect 111260 600 111288 1340
rect 113100 600 113128 1340
rect 114940 600 114968 1340
rect 116688 600 116716 1340
rect 118528 600 118556 1340
rect 120368 600 120396 1340
rect 122208 600 122236 1340
rect 124048 600 124076 1340
rect 125888 600 125916 1340
rect 127728 600 127756 1340
rect 129568 600 129596 1340
rect 131408 600 131436 1340
rect 133156 600 133184 1340
rect 134996 600 135024 1340
rect 136836 600 136864 1340
rect 138952 626 138980 1340
rect 138676 600 138980 626
rect 140516 600 140544 1340
rect 142356 600 142384 1340
rect 144196 600 144224 1340
rect 146036 600 146064 1340
rect 147784 600 147812 1340
rect 149624 600 149652 1340
rect 151464 600 151492 1340
rect 153304 600 153332 1340
rect 155144 600 155172 1340
rect 156984 600 157012 1340
rect 158824 600 158852 1340
rect 160664 600 160692 1340
rect 162504 600 162532 1340
rect 164252 600 164280 1340
rect 166092 600 166120 1340
rect 167932 600 167960 1340
rect 169772 600 169800 1340
rect 171612 600 171640 1340
rect 173452 600 173480 1340
rect 175292 600 175320 1340
rect 177132 600 177160 1340
rect 178972 600 179000 1340
rect 180720 600 180748 1340
rect 182008 600 182036 1340
rect 182560 600 182588 1340
rect 183848 600 183876 1340
rect 184400 600 184428 1340
rect 185596 600 185624 1340
rect 186240 600 186268 1340
rect 187436 600 187464 1340
rect 188080 600 188108 1340
rect 189276 600 189304 1340
rect 189920 600 189948 1340
rect 191116 600 191144 1340
rect 191760 600 191788 1340
rect 192956 600 192984 1340
rect 193600 600 193628 1340
rect 194796 600 194824 1340
rect 195348 600 195376 1340
rect 196636 600 196664 1340
rect 197188 600 197216 1340
rect 198476 600 198504 1340
rect 199028 600 199056 1340
rect 200316 600 200344 1340
rect 200868 600 200896 1340
rect 202064 600 202092 1340
rect 202708 600 202736 1340
rect 203904 600 203932 1340
rect 204548 600 204576 1340
rect 205744 600 205772 1340
rect 206388 600 206416 1340
rect 207584 600 207612 1340
rect 208228 600 208256 1340
rect 209424 600 209452 1340
rect 210068 600 210096 1340
rect 211264 600 211292 1340
rect 211816 600 211844 1340
rect 213104 600 213132 1340
rect 213656 600 213684 1340
rect 214944 600 214972 1340
rect 215496 600 215524 1340
rect 216692 600 216720 1340
rect 217336 600 217364 1340
rect 218532 600 218560 1340
rect 219176 600 219204 1340
rect 220372 600 220400 1340
rect 221016 600 221044 1340
rect 222212 600 222240 1340
rect 222856 600 222884 1340
rect 224052 600 224080 1340
rect 224696 600 224724 1340
rect 225892 600 225920 1340
rect 226536 600 226564 1340
rect 227732 600 227760 1340
rect 228284 600 228312 1340
rect 229572 600 229600 1340
rect 230124 600 230152 1340
rect 231412 600 231440 1340
rect 231964 600 231992 1340
rect 233160 600 233188 1340
rect 233804 600 233832 1340
rect 235000 600 235028 1340
rect 235644 600 235672 1340
rect 236840 600 236868 1340
rect 237484 600 237512 1340
rect 238680 600 238708 1340
rect 239324 600 239352 1340
rect 240520 600 240548 1340
rect 241164 600 241192 1340
rect 242360 600 242388 1340
rect 242912 600 242940 1340
rect 244200 600 244228 1340
rect 244752 600 244780 1340
rect 246040 600 246068 1340
rect 246592 600 246620 1340
rect 247788 600 247816 1340
rect 248432 600 248460 1340
rect 249628 600 249656 1340
rect 250272 600 250300 1340
rect 251468 600 251496 1340
rect 252112 600 252140 1340
rect 253308 600 253336 1340
rect 253952 600 253980 1340
rect 255148 600 255176 1340
rect 255792 600 255820 1340
rect 256988 600 257016 1340
rect 257632 600 257660 1340
rect 258828 600 258856 1340
rect 259380 600 259408 1340
rect 260668 600 260696 1340
rect 261220 600 261248 1340
rect 262508 600 262536 1340
rect 263060 600 263088 1340
rect 264256 600 264284 1340
rect 264900 600 264928 1340
rect 266096 600 266124 1340
rect 266740 600 266768 1340
rect 267936 600 267964 1340
rect 268580 600 268608 1340
rect 269132 762 269160 1340
rect 269132 734 269712 762
rect 269684 626 269712 734
rect 269684 600 269804 626
rect 270420 600 270448 1340
rect 271524 626 271552 1340
rect 271524 600 271644 626
rect 272260 600 272288 1340
rect 274008 600 274036 1340
rect 275848 600 275876 1340
rect 277688 600 277716 1340
rect 279528 600 279556 1340
rect 281368 600 281396 1340
rect 283208 600 283236 1340
rect 285048 600 285076 1340
rect 286888 600 286916 1340
rect 288728 600 288756 1340
rect 290476 600 290504 1340
rect 292316 600 292344 1340
rect 294156 600 294184 1340
rect 295996 600 296024 1340
rect 297836 600 297864 1340
rect 266 -1200 378 600
rect 818 -1200 930 600
rect 1462 -1200 1574 600
rect 2014 -1200 2126 600
rect 2658 -1200 2770 600
rect 3302 -1200 3414 600
rect 3854 -1200 3966 600
rect 4498 -1200 4610 600
rect 5142 -1200 5254 600
rect 5694 -1200 5806 600
rect 6338 -1200 6450 600
rect 6890 -1200 7002 600
rect 7534 -1200 7646 600
rect 8178 -1200 8290 600
rect 8730 -1200 8842 600
rect 9374 -1200 9486 600
rect 10018 -1200 10130 600
rect 10570 -1200 10682 600
rect 11214 -1200 11326 600
rect 11766 -1200 11878 600
rect 12410 -1200 12522 600
rect 13054 -1200 13166 600
rect 13606 -1200 13718 600
rect 14250 -1200 14362 600
rect 14894 -1200 15006 600
rect 15446 -1200 15558 600
rect 16090 -1200 16202 600
rect 16642 -1200 16754 600
rect 17286 -1200 17398 600
rect 17930 -1200 18042 600
rect 18482 -1200 18594 600
rect 19126 -1200 19238 600
rect 19770 -1200 19882 600
rect 20322 -1200 20434 600
rect 20966 -1200 21078 600
rect 21518 -1200 21630 600
rect 22162 -1200 22274 600
rect 22806 -1200 22918 600
rect 23358 -1200 23470 600
rect 24002 -1200 24114 600
rect 24646 -1200 24758 600
rect 25198 -1200 25310 600
rect 25842 -1200 25954 600
rect 26486 -1200 26598 600
rect 27038 -1200 27150 600
rect 27682 -1200 27794 600
rect 28234 -1200 28346 600
rect 28878 -1200 28990 600
rect 29522 -1200 29634 600
rect 30074 -1200 30186 600
rect 30718 -1200 30830 600
rect 31362 -1200 31474 600
rect 31914 -1200 32026 600
rect 32558 -1200 32670 600
rect 33110 -1200 33222 600
rect 33754 -1200 33866 600
rect 34398 -1200 34510 600
rect 34950 -1200 35062 600
rect 35594 -1200 35706 600
rect 36238 -1200 36350 600
rect 36790 -1200 36902 600
rect 37434 -1200 37546 600
rect 37986 -1200 38098 600
rect 38630 -1200 38742 600
rect 39274 -1200 39386 600
rect 39826 -1200 39938 600
rect 40470 -1200 40582 600
rect 41114 -1200 41226 600
rect 41666 598 41828 600
rect 41666 -1200 41778 598
rect 42310 -1200 42422 600
rect 42862 -1200 42974 600
rect 43506 -1200 43618 600
rect 44150 -1200 44262 600
rect 44702 -1200 44814 600
rect 45346 -1200 45458 600
rect 45990 -1200 46102 600
rect 46542 -1200 46654 600
rect 47186 -1200 47298 600
rect 47738 -1200 47850 600
rect 48382 -1200 48494 600
rect 49026 -1200 49138 600
rect 49578 -1200 49690 600
rect 50222 -1200 50334 600
rect 50866 -1200 50978 600
rect 51368 598 51530 600
rect 51418 -1200 51530 598
rect 52062 -1200 52174 600
rect 52706 -1200 52818 600
rect 53258 -1200 53370 600
rect 53902 -1200 54014 600
rect 54312 598 54566 600
rect 54454 -1200 54566 598
rect 55098 598 55260 600
rect 55098 -1200 55210 598
rect 55742 -1200 55854 600
rect 56152 598 56406 600
rect 56294 -1200 56406 598
rect 56938 -1200 57050 600
rect 57582 -1200 57694 600
rect 58134 -1200 58246 600
rect 58778 -1200 58890 600
rect 59330 -1200 59442 600
rect 59974 598 60136 600
rect 59974 -1200 60086 598
rect 60618 -1200 60730 600
rect 61170 -1200 61282 600
rect 61814 -1200 61926 600
rect 62458 -1200 62570 600
rect 63010 -1200 63122 600
rect 63654 -1200 63766 600
rect 64206 -1200 64318 600
rect 64850 -1200 64962 600
rect 65494 -1200 65606 600
rect 66046 -1200 66158 600
rect 66690 -1200 66802 600
rect 67334 -1200 67446 600
rect 67886 -1200 67998 600
rect 68530 -1200 68642 600
rect 69082 -1200 69194 600
rect 69726 -1200 69838 600
rect 70370 -1200 70482 600
rect 70922 -1200 71034 600
rect 71566 -1200 71678 600
rect 72210 -1200 72322 600
rect 72762 -1200 72874 600
rect 73406 -1200 73518 600
rect 73958 -1200 74070 600
rect 74602 -1200 74714 600
rect 75246 -1200 75358 600
rect 75798 -1200 75910 600
rect 76442 -1200 76554 600
rect 77086 -1200 77198 600
rect 77638 -1200 77750 600
rect 78282 598 78628 600
rect 78282 -1200 78394 598
rect 78926 -1200 79038 600
rect 79478 -1200 79590 600
rect 80122 -1200 80234 600
rect 80674 -1200 80786 600
rect 81318 -1200 81430 600
rect 81962 -1200 82074 600
rect 82514 -1200 82626 600
rect 83158 -1200 83270 600
rect 83802 598 84148 600
rect 83802 -1200 83914 598
rect 84354 -1200 84466 600
rect 84998 -1200 85110 600
rect 85550 -1200 85662 600
rect 86194 -1200 86306 600
rect 86838 -1200 86950 600
rect 87390 -1200 87502 600
rect 88034 -1200 88146 600
rect 88678 -1200 88790 600
rect 89230 -1200 89342 600
rect 89874 -1200 89986 600
rect 90426 -1200 90538 600
rect 91070 -1200 91182 600
rect 91714 -1200 91826 600
rect 92266 -1200 92378 600
rect 92910 -1200 93022 600
rect 93554 -1200 93666 600
rect 94106 -1200 94218 600
rect 94750 -1200 94862 600
rect 95302 -1200 95414 600
rect 95946 -1200 96058 600
rect 96590 -1200 96702 600
rect 97142 -1200 97254 600
rect 97786 -1200 97898 600
rect 98430 -1200 98542 600
rect 98982 -1200 99094 600
rect 99626 -1200 99738 600
rect 100270 598 100708 600
rect 100270 -1200 100382 598
rect 100822 -1200 100934 600
rect 101466 -1200 101578 600
rect 102018 -1200 102130 600
rect 102662 -1200 102774 600
rect 103306 -1200 103418 600
rect 103858 -1200 103970 600
rect 104502 -1200 104614 600
rect 105146 -1200 105258 600
rect 105698 -1200 105810 600
rect 106342 -1200 106454 600
rect 106894 -1200 107006 600
rect 107538 -1200 107650 600
rect 108182 -1200 108294 600
rect 108734 -1200 108846 600
rect 109378 -1200 109490 600
rect 110022 -1200 110134 600
rect 110574 -1200 110686 600
rect 111218 -1200 111330 600
rect 111770 -1200 111882 600
rect 112414 -1200 112526 600
rect 113058 -1200 113170 600
rect 113610 -1200 113722 600
rect 114254 -1200 114366 600
rect 114898 -1200 115010 600
rect 115450 -1200 115562 600
rect 116094 -1200 116206 600
rect 116646 -1200 116758 600
rect 117290 -1200 117402 600
rect 117934 -1200 118046 600
rect 118486 -1200 118598 600
rect 119130 -1200 119242 600
rect 119774 -1200 119886 600
rect 120326 -1200 120438 600
rect 120970 -1200 121082 600
rect 121522 -1200 121634 600
rect 122166 -1200 122278 600
rect 122810 -1200 122922 600
rect 123362 -1200 123474 600
rect 124006 -1200 124118 600
rect 124650 -1200 124762 600
rect 125202 -1200 125314 600
rect 125846 -1200 125958 600
rect 126490 -1200 126602 600
rect 127042 -1200 127154 600
rect 127686 -1200 127798 600
rect 128238 -1200 128350 600
rect 128882 -1200 128994 600
rect 129526 -1200 129638 600
rect 130078 -1200 130190 600
rect 130722 -1200 130834 600
rect 131366 -1200 131478 600
rect 131918 -1200 132030 600
rect 132562 -1200 132674 600
rect 133114 -1200 133226 600
rect 133758 -1200 133870 600
rect 134402 -1200 134514 600
rect 134954 -1200 135066 600
rect 135598 -1200 135710 600
rect 136242 -1200 136354 600
rect 136794 -1200 136906 600
rect 137438 -1200 137550 600
rect 137990 -1200 138102 600
rect 138634 598 138980 600
rect 138634 -1200 138746 598
rect 139278 -1200 139390 600
rect 139830 -1200 139942 600
rect 140474 -1200 140586 600
rect 141118 -1200 141230 600
rect 141670 -1200 141782 600
rect 142314 -1200 142426 600
rect 142866 -1200 142978 600
rect 143510 -1200 143622 600
rect 144154 -1200 144266 600
rect 144706 -1200 144818 600
rect 145350 -1200 145462 600
rect 145994 -1200 146106 600
rect 146546 -1200 146658 600
rect 147190 -1200 147302 600
rect 147742 -1200 147854 600
rect 148386 -1200 148498 600
rect 149030 -1200 149142 600
rect 149582 -1200 149694 600
rect 150226 -1200 150338 600
rect 150870 -1200 150982 600
rect 151422 -1200 151534 600
rect 152066 -1200 152178 600
rect 152710 -1200 152822 600
rect 153262 -1200 153374 600
rect 153906 -1200 154018 600
rect 154458 -1200 154570 600
rect 155102 -1200 155214 600
rect 155746 -1200 155858 600
rect 156298 -1200 156410 600
rect 156942 -1200 157054 600
rect 157586 -1200 157698 600
rect 158138 -1200 158250 600
rect 158782 -1200 158894 600
rect 159334 -1200 159446 600
rect 159978 -1200 160090 600
rect 160622 -1200 160734 600
rect 161174 -1200 161286 600
rect 161818 -1200 161930 600
rect 162462 -1200 162574 600
rect 163014 -1200 163126 600
rect 163658 -1200 163770 600
rect 164210 -1200 164322 600
rect 164854 -1200 164966 600
rect 165498 -1200 165610 600
rect 166050 -1200 166162 600
rect 166694 -1200 166806 600
rect 167338 -1200 167450 600
rect 167890 -1200 168002 600
rect 168534 -1200 168646 600
rect 169086 -1200 169198 600
rect 169730 -1200 169842 600
rect 170374 -1200 170486 600
rect 170926 -1200 171038 600
rect 171570 -1200 171682 600
rect 172214 -1200 172326 600
rect 172766 -1200 172878 600
rect 173410 -1200 173522 600
rect 173962 -1200 174074 600
rect 174606 -1200 174718 600
rect 175250 -1200 175362 600
rect 175802 -1200 175914 600
rect 176446 -1200 176558 600
rect 177090 -1200 177202 600
rect 177642 -1200 177754 600
rect 178286 -1200 178398 600
rect 178930 -1200 179042 600
rect 179482 -1200 179594 600
rect 180126 -1200 180238 600
rect 180678 -1200 180790 600
rect 181322 -1200 181434 600
rect 181966 -1200 182078 600
rect 182518 -1200 182630 600
rect 183162 -1200 183274 600
rect 183806 -1200 183918 600
rect 184358 -1200 184470 600
rect 185002 -1200 185114 600
rect 185554 -1200 185666 600
rect 186198 -1200 186310 600
rect 186842 -1200 186954 600
rect 187394 -1200 187506 600
rect 188038 -1200 188150 600
rect 188682 -1200 188794 600
rect 189234 -1200 189346 600
rect 189878 -1200 189990 600
rect 190430 -1200 190542 600
rect 191074 -1200 191186 600
rect 191718 -1200 191830 600
rect 192270 -1200 192382 600
rect 192914 -1200 193026 600
rect 193558 -1200 193670 600
rect 194110 -1200 194222 600
rect 194754 -1200 194866 600
rect 195306 -1200 195418 600
rect 195950 -1200 196062 600
rect 196594 -1200 196706 600
rect 197146 -1200 197258 600
rect 197790 -1200 197902 600
rect 198434 -1200 198546 600
rect 198986 -1200 199098 600
rect 199630 -1200 199742 600
rect 200274 -1200 200386 600
rect 200826 -1200 200938 600
rect 201470 -1200 201582 600
rect 202022 -1200 202134 600
rect 202666 -1200 202778 600
rect 203310 -1200 203422 600
rect 203862 -1200 203974 600
rect 204506 -1200 204618 600
rect 205150 -1200 205262 600
rect 205702 -1200 205814 600
rect 206346 -1200 206458 600
rect 206898 -1200 207010 600
rect 207542 -1200 207654 600
rect 208186 -1200 208298 600
rect 208738 -1200 208850 600
rect 209382 -1200 209494 600
rect 210026 -1200 210138 600
rect 210578 -1200 210690 600
rect 211222 -1200 211334 600
rect 211774 -1200 211886 600
rect 212418 -1200 212530 600
rect 213062 -1200 213174 600
rect 213614 -1200 213726 600
rect 214258 -1200 214370 600
rect 214902 -1200 215014 600
rect 215454 -1200 215566 600
rect 216098 -1200 216210 600
rect 216650 -1200 216762 600
rect 217294 -1200 217406 600
rect 217938 -1200 218050 600
rect 218490 -1200 218602 600
rect 219134 -1200 219246 600
rect 219778 -1200 219890 600
rect 220330 -1200 220442 600
rect 220974 -1200 221086 600
rect 221526 -1200 221638 600
rect 222170 -1200 222282 600
rect 222814 -1200 222926 600
rect 223366 -1200 223478 600
rect 224010 -1200 224122 600
rect 224654 -1200 224766 600
rect 225206 -1200 225318 600
rect 225850 -1200 225962 600
rect 226494 -1200 226606 600
rect 227046 -1200 227158 600
rect 227690 -1200 227802 600
rect 228242 -1200 228354 600
rect 228886 -1200 228998 600
rect 229530 -1200 229642 600
rect 230082 -1200 230194 600
rect 230726 -1200 230838 600
rect 231370 -1200 231482 600
rect 231922 -1200 232034 600
rect 232566 -1200 232678 600
rect 233118 -1200 233230 600
rect 233762 -1200 233874 600
rect 234406 -1200 234518 600
rect 234958 -1200 235070 600
rect 235602 -1200 235714 600
rect 236246 -1200 236358 600
rect 236798 -1200 236910 600
rect 237442 -1200 237554 600
rect 237994 -1200 238106 600
rect 238638 -1200 238750 600
rect 239282 -1200 239394 600
rect 239834 -1200 239946 600
rect 240478 -1200 240590 600
rect 241122 -1200 241234 600
rect 241674 -1200 241786 600
rect 242318 -1200 242430 600
rect 242870 -1200 242982 600
rect 243514 -1200 243626 600
rect 244158 -1200 244270 600
rect 244710 -1200 244822 600
rect 245354 -1200 245466 600
rect 245998 -1200 246110 600
rect 246550 -1200 246662 600
rect 247194 -1200 247306 600
rect 247746 -1200 247858 600
rect 248390 -1200 248502 600
rect 249034 -1200 249146 600
rect 249586 -1200 249698 600
rect 250230 -1200 250342 600
rect 250874 -1200 250986 600
rect 251426 -1200 251538 600
rect 252070 -1200 252182 600
rect 252714 -1200 252826 600
rect 253266 -1200 253378 600
rect 253910 -1200 254022 600
rect 254462 -1200 254574 600
rect 255106 -1200 255218 600
rect 255750 -1200 255862 600
rect 256302 -1200 256414 600
rect 256946 -1200 257058 600
rect 257590 -1200 257702 600
rect 258142 -1200 258254 600
rect 258786 -1200 258898 600
rect 259338 -1200 259450 600
rect 259982 -1200 260094 600
rect 260626 -1200 260738 600
rect 261178 -1200 261290 600
rect 261822 -1200 261934 600
rect 262466 -1200 262578 600
rect 263018 -1200 263130 600
rect 263662 -1200 263774 600
rect 264214 -1200 264326 600
rect 264858 -1200 264970 600
rect 265502 -1200 265614 600
rect 266054 -1200 266166 600
rect 266698 -1200 266810 600
rect 267342 -1200 267454 600
rect 267894 -1200 268006 600
rect 268538 -1200 268650 600
rect 269090 -1200 269202 600
rect 269684 598 269846 600
rect 269734 -1200 269846 598
rect 270378 -1200 270490 600
rect 270930 -1200 271042 600
rect 271524 598 271686 600
rect 271574 -1200 271686 598
rect 272218 -1200 272330 600
rect 272770 -1200 272882 600
rect 273414 -1200 273526 600
rect 273966 -1200 274078 600
rect 274610 -1200 274722 600
rect 275254 -1200 275366 600
rect 275806 -1200 275918 600
rect 276450 -1200 276562 600
rect 277094 -1200 277206 600
rect 277646 -1200 277758 600
rect 278290 -1200 278402 600
rect 278934 -1200 279046 600
rect 279486 -1200 279598 600
rect 280130 -1200 280242 600
rect 280682 -1200 280794 600
rect 281326 -1200 281438 600
rect 281970 -1200 282082 600
rect 282522 -1200 282634 600
rect 283166 -1200 283278 600
rect 283810 -1200 283922 600
rect 284362 -1200 284474 600
rect 285006 -1200 285118 600
rect 285558 -1200 285670 600
rect 286202 -1200 286314 600
rect 286846 -1200 286958 600
rect 287398 -1200 287510 600
rect 288042 -1200 288154 600
rect 288686 -1200 288798 600
rect 289238 -1200 289350 600
rect 289882 -1200 289994 600
rect 290434 -1200 290546 600
rect 291078 -1200 291190 600
rect 291722 -1200 291834 600
rect 292274 -1200 292386 600
rect 292918 -1200 293030 600
rect 293562 -1200 293674 600
rect 294114 -1200 294226 600
rect 294758 -1200 294870 600
rect 295310 -1200 295422 600
rect 295954 -1200 296066 600
rect 296598 -1200 296710 600
rect 297150 -1200 297262 600
rect 297794 -1200 297906 600
rect 298438 -1200 298550 600
rect 298990 -1200 299102 600
rect 299634 -1200 299746 600
<< obsm2 >>
rect 1492 1340 297876 298660
<< metal3 >>
rect -1200 224892 600 225132
rect -1200 74884 600 75124
rect 299400 249780 301200 250020
rect 299400 149820 301200 150060
rect 299400 49860 301200 50100
<< obsm3 >>
rect 4848 2143 297008 297601
<< metal4 >>
rect -136 298786 464 298808
rect -136 298550 46 298786
rect 282 298550 464 298786
rect 4848 298660 5168 298808
rect 20208 298786 20528 298808
rect 20208 298660 20250 298786
rect 20486 298660 20528 298786
rect 35568 298660 35888 298808
rect 50928 298786 51248 298808
rect 50928 298660 50970 298786
rect 51206 298660 51248 298786
rect 66288 298660 66608 298808
rect 81648 298786 81968 298808
rect 81648 298660 81690 298786
rect 81926 298660 81968 298786
rect 97008 298660 97328 298808
rect 112368 298786 112688 298808
rect 112368 298660 112410 298786
rect 112646 298660 112688 298786
rect 127728 298660 128048 298808
rect 143088 298786 143408 298808
rect 143088 298660 143130 298786
rect 143366 298660 143408 298786
rect 158448 298660 158768 298808
rect 173808 298786 174128 298808
rect 173808 298660 173850 298786
rect 174086 298660 174128 298786
rect 189168 298660 189488 298808
rect 204528 298786 204848 298808
rect 204528 298660 204570 298786
rect 204806 298660 204848 298786
rect 219888 298660 220208 298808
rect 235248 298786 235568 298808
rect 235248 298660 235290 298786
rect 235526 298660 235568 298786
rect 250608 298660 250928 298808
rect 265968 298786 266288 298808
rect 265968 298660 266010 298786
rect 266246 298660 266288 298786
rect 281328 298660 281648 298808
rect 296688 298786 297008 298808
rect 296688 298660 296730 298786
rect 296966 298660 297008 298786
rect 299456 298786 300056 298808
rect -136 298466 464 298550
rect -136 298230 46 298466
rect 282 298230 464 298466
rect -136 289647 464 298230
rect -136 289411 46 289647
rect 282 289411 464 289647
rect -136 274329 464 289411
rect -136 274093 46 274329
rect 282 274093 464 274329
rect -136 259011 464 274093
rect -136 258775 46 259011
rect 282 258775 464 259011
rect -136 243693 464 258775
rect -136 243457 46 243693
rect 282 243457 464 243693
rect -136 228375 464 243457
rect -136 228139 46 228375
rect 282 228139 464 228375
rect -136 213057 464 228139
rect -136 212821 46 213057
rect 282 212821 464 213057
rect -136 197739 464 212821
rect -136 197503 46 197739
rect 282 197503 464 197739
rect -136 182421 464 197503
rect -136 182185 46 182421
rect 282 182185 464 182421
rect -136 167103 464 182185
rect -136 166867 46 167103
rect 282 166867 464 167103
rect -136 151785 464 166867
rect -136 151549 46 151785
rect 282 151549 464 151785
rect -136 136467 464 151549
rect -136 136231 46 136467
rect 282 136231 464 136467
rect -136 121149 464 136231
rect -136 120913 46 121149
rect 282 120913 464 121149
rect -136 105831 464 120913
rect -136 105595 46 105831
rect 282 105595 464 105831
rect -136 90513 464 105595
rect -136 90277 46 90513
rect 282 90277 464 90513
rect -136 75195 464 90277
rect -136 74959 46 75195
rect 282 74959 464 75195
rect -136 59877 464 74959
rect -136 59641 46 59877
rect 282 59641 464 59877
rect -136 44559 464 59641
rect -136 44323 46 44559
rect 282 44323 464 44559
rect -136 29241 464 44323
rect -136 29005 46 29241
rect 282 29005 464 29241
rect -136 13923 464 29005
rect -136 13687 46 13923
rect 282 13687 464 13923
rect -136 1514 464 13687
rect 804 297846 1340 297868
rect 804 297610 986 297846
rect 1222 297610 1340 297846
rect 804 297526 1340 297610
rect 804 297290 986 297526
rect 1222 297290 1340 297526
rect 804 281988 1340 297290
rect 804 281752 986 281988
rect 1222 281752 1340 281988
rect 804 266670 1340 281752
rect 804 266434 986 266670
rect 1222 266434 1340 266670
rect 804 251352 1340 266434
rect 804 251116 986 251352
rect 1222 251116 1340 251352
rect 804 236034 1340 251116
rect 804 235798 986 236034
rect 1222 235798 1340 236034
rect 804 220716 1340 235798
rect 804 220480 986 220716
rect 1222 220480 1340 220716
rect 804 205398 1340 220480
rect 804 205162 986 205398
rect 1222 205162 1340 205398
rect 804 190080 1340 205162
rect 804 189844 986 190080
rect 1222 189844 1340 190080
rect 804 174762 1340 189844
rect 804 174526 986 174762
rect 1222 174526 1340 174762
rect 804 159444 1340 174526
rect 804 159208 986 159444
rect 1222 159208 1340 159444
rect 804 144126 1340 159208
rect 804 143890 986 144126
rect 1222 143890 1340 144126
rect 804 128808 1340 143890
rect 804 128572 986 128808
rect 1222 128572 1340 128808
rect 804 113490 1340 128572
rect 804 113254 986 113490
rect 1222 113254 1340 113490
rect 804 98172 1340 113254
rect 804 97936 986 98172
rect 1222 97936 1340 98172
rect 804 82854 1340 97936
rect 804 82618 986 82854
rect 1222 82618 1340 82854
rect 804 67536 1340 82618
rect 804 67300 986 67536
rect 1222 67300 1340 67536
rect 804 52218 1340 67300
rect 804 51982 986 52218
rect 1222 51982 1340 52218
rect 804 36900 1340 51982
rect 804 36664 986 36900
rect 1222 36664 1340 36900
rect 804 21582 1340 36664
rect 804 21346 986 21582
rect 1222 21346 1340 21582
rect 804 6264 1340 21346
rect 804 6028 986 6264
rect 1222 6028 1340 6264
rect 804 2454 1340 6028
rect 804 2218 986 2454
rect 1222 2218 1340 2454
rect 804 2134 1340 2218
rect 804 1898 986 2134
rect 1222 1898 1340 2134
rect 804 1876 1340 1898
rect -136 1278 46 1514
rect 282 1278 464 1514
rect 299456 298550 299638 298786
rect 299874 298550 300056 298786
rect 299456 298466 300056 298550
rect 299456 298230 299638 298466
rect 299874 298230 300056 298466
rect 298660 297846 299116 297868
rect 298660 297610 298698 297846
rect 298934 297610 299116 297846
rect 298660 297526 299116 297610
rect 298660 297290 298698 297526
rect 298934 297290 299116 297526
rect 298660 281988 299116 297290
rect 298660 281752 298698 281988
rect 298934 281752 299116 281988
rect 298660 266670 299116 281752
rect 298660 266434 298698 266670
rect 298934 266434 299116 266670
rect 298660 251352 299116 266434
rect 298660 251116 298698 251352
rect 298934 251116 299116 251352
rect 298660 236034 299116 251116
rect 298660 235798 298698 236034
rect 298934 235798 299116 236034
rect 298660 220716 299116 235798
rect 298660 220480 298698 220716
rect 298934 220480 299116 220716
rect 298660 205398 299116 220480
rect 298660 205162 298698 205398
rect 298934 205162 299116 205398
rect 298660 190080 299116 205162
rect 298660 189844 298698 190080
rect 298934 189844 299116 190080
rect 298660 174762 299116 189844
rect 298660 174526 298698 174762
rect 298934 174526 299116 174762
rect 298660 159444 299116 174526
rect 298660 159208 298698 159444
rect 298934 159208 299116 159444
rect 298660 144126 299116 159208
rect 298660 143890 298698 144126
rect 298934 143890 299116 144126
rect 298660 128808 299116 143890
rect 298660 128572 298698 128808
rect 298934 128572 299116 128808
rect 298660 113490 299116 128572
rect 298660 113254 298698 113490
rect 298934 113254 299116 113490
rect 298660 98172 299116 113254
rect 298660 97936 298698 98172
rect 298934 97936 299116 98172
rect 298660 82854 299116 97936
rect 298660 82618 298698 82854
rect 298934 82618 299116 82854
rect 298660 67536 299116 82618
rect 298660 67300 298698 67536
rect 298934 67300 299116 67536
rect 298660 52218 299116 67300
rect 298660 51982 298698 52218
rect 298934 51982 299116 52218
rect 298660 36900 299116 51982
rect 298660 36664 298698 36900
rect 298934 36664 299116 36900
rect 298660 21582 299116 36664
rect 298660 21346 298698 21582
rect 298934 21346 299116 21582
rect 298660 6264 299116 21346
rect 298660 6028 298698 6264
rect 298934 6028 299116 6264
rect 298660 2454 299116 6028
rect 298660 2218 298698 2454
rect 298934 2218 299116 2454
rect 298660 2134 299116 2218
rect 298660 1898 298698 2134
rect 298934 1898 299116 2134
rect 298660 1876 299116 1898
rect 299456 289647 300056 298230
rect 299456 289411 299638 289647
rect 299874 289411 300056 289647
rect 299456 274329 300056 289411
rect 299456 274093 299638 274329
rect 299874 274093 300056 274329
rect 299456 259011 300056 274093
rect 299456 258775 299638 259011
rect 299874 258775 300056 259011
rect 299456 243693 300056 258775
rect 299456 243457 299638 243693
rect 299874 243457 300056 243693
rect 299456 228375 300056 243457
rect 299456 228139 299638 228375
rect 299874 228139 300056 228375
rect 299456 213057 300056 228139
rect 299456 212821 299638 213057
rect 299874 212821 300056 213057
rect 299456 197739 300056 212821
rect 299456 197503 299638 197739
rect 299874 197503 300056 197739
rect 299456 182421 300056 197503
rect 299456 182185 299638 182421
rect 299874 182185 300056 182421
rect 299456 167103 300056 182185
rect 299456 166867 299638 167103
rect 299874 166867 300056 167103
rect 299456 151785 300056 166867
rect 299456 151549 299638 151785
rect 299874 151549 300056 151785
rect 299456 136467 300056 151549
rect 299456 136231 299638 136467
rect 299874 136231 300056 136467
rect 299456 121149 300056 136231
rect 299456 120913 299638 121149
rect 299874 120913 300056 121149
rect 299456 105831 300056 120913
rect 299456 105595 299638 105831
rect 299874 105595 300056 105831
rect 299456 90513 300056 105595
rect 299456 90277 299638 90513
rect 299874 90277 300056 90513
rect 299456 75195 300056 90277
rect 299456 74959 299638 75195
rect 299874 74959 300056 75195
rect 299456 59877 300056 74959
rect 299456 59641 299638 59877
rect 299874 59641 300056 59877
rect 299456 44559 300056 59641
rect 299456 44323 299638 44559
rect 299874 44323 300056 44559
rect 299456 29241 300056 44323
rect 299456 29005 299638 29241
rect 299874 29005 300056 29241
rect 299456 13923 300056 29005
rect 299456 13687 299638 13923
rect 299874 13687 300056 13923
rect 299456 1514 300056 13687
rect -136 1194 464 1278
rect -136 958 46 1194
rect 282 958 464 1194
rect -136 936 464 958
rect 4848 936 5168 1340
rect 20208 1278 20250 1340
rect 20486 1278 20528 1340
rect 20208 1194 20528 1278
rect 20208 958 20250 1194
rect 20486 958 20528 1194
rect 20208 936 20528 958
rect 35568 936 35888 1340
rect 50928 1278 50970 1340
rect 51206 1278 51248 1340
rect 50928 1194 51248 1278
rect 50928 958 50970 1194
rect 51206 958 51248 1194
rect 50928 936 51248 958
rect 66288 936 66608 1340
rect 81648 1278 81690 1340
rect 81926 1278 81968 1340
rect 81648 1194 81968 1278
rect 81648 958 81690 1194
rect 81926 958 81968 1194
rect 81648 936 81968 958
rect 97008 936 97328 1340
rect 112368 1278 112410 1340
rect 112646 1278 112688 1340
rect 112368 1194 112688 1278
rect 112368 958 112410 1194
rect 112646 958 112688 1194
rect 112368 936 112688 958
rect 127728 936 128048 1340
rect 143088 1278 143130 1340
rect 143366 1278 143408 1340
rect 143088 1194 143408 1278
rect 143088 958 143130 1194
rect 143366 958 143408 1194
rect 143088 936 143408 958
rect 158448 936 158768 1340
rect 173808 1278 173850 1340
rect 174086 1278 174128 1340
rect 173808 1194 174128 1278
rect 173808 958 173850 1194
rect 174086 958 174128 1194
rect 173808 936 174128 958
rect 189168 936 189488 1340
rect 204528 1278 204570 1340
rect 204806 1278 204848 1340
rect 204528 1194 204848 1278
rect 204528 958 204570 1194
rect 204806 958 204848 1194
rect 204528 936 204848 958
rect 219888 936 220208 1340
rect 235248 1278 235290 1340
rect 235526 1278 235568 1340
rect 235248 1194 235568 1278
rect 235248 958 235290 1194
rect 235526 958 235568 1194
rect 235248 936 235568 958
rect 250608 936 250928 1340
rect 265968 1278 266010 1340
rect 266246 1278 266288 1340
rect 265968 1194 266288 1278
rect 265968 958 266010 1194
rect 266246 958 266288 1194
rect 265968 936 266288 958
rect 281328 936 281648 1340
rect 296688 1278 296730 1340
rect 296966 1278 297008 1340
rect 296688 1194 297008 1278
rect 296688 958 296730 1194
rect 296966 958 297008 1194
rect 296688 936 297008 958
rect 299456 1278 299638 1514
rect 299874 1278 300056 1514
rect 299456 1194 300056 1278
rect 299456 958 299638 1194
rect 299874 958 300056 1194
rect 299456 936 300056 958
<< obsm4 >>
rect 1340 1340 298660 298660
<< via4 >>
rect 46 298550 282 298786
rect 20250 298660 20486 298786
rect 50970 298660 51206 298786
rect 81690 298660 81926 298786
rect 112410 298660 112646 298786
rect 143130 298660 143366 298786
rect 173850 298660 174086 298786
rect 204570 298660 204806 298786
rect 235290 298660 235526 298786
rect 266010 298660 266246 298786
rect 296730 298660 296966 298786
rect 46 298230 282 298466
rect 46 289411 282 289647
rect 46 274093 282 274329
rect 46 258775 282 259011
rect 46 243457 282 243693
rect 46 228139 282 228375
rect 46 212821 282 213057
rect 46 197503 282 197739
rect 46 182185 282 182421
rect 46 166867 282 167103
rect 46 151549 282 151785
rect 46 136231 282 136467
rect 46 120913 282 121149
rect 46 105595 282 105831
rect 46 90277 282 90513
rect 46 74959 282 75195
rect 46 59641 282 59877
rect 46 44323 282 44559
rect 46 29005 282 29241
rect 46 13687 282 13923
rect 986 297610 1222 297846
rect 986 297290 1222 297526
rect 986 281752 1222 281988
rect 986 266434 1222 266670
rect 986 251116 1222 251352
rect 986 235798 1222 236034
rect 986 220480 1222 220716
rect 986 205162 1222 205398
rect 986 189844 1222 190080
rect 986 174526 1222 174762
rect 986 159208 1222 159444
rect 986 143890 1222 144126
rect 986 128572 1222 128808
rect 986 113254 1222 113490
rect 986 97936 1222 98172
rect 986 82618 1222 82854
rect 986 67300 1222 67536
rect 986 51982 1222 52218
rect 986 36664 1222 36900
rect 986 21346 1222 21582
rect 986 6028 1222 6264
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 46 1278 282 1514
rect 299638 298550 299874 298786
rect 299638 298230 299874 298466
rect 298698 297610 298934 297846
rect 298698 297290 298934 297526
rect 298698 281752 298934 281988
rect 298698 266434 298934 266670
rect 298698 251116 298934 251352
rect 298698 235798 298934 236034
rect 298698 220480 298934 220716
rect 298698 205162 298934 205398
rect 298698 189844 298934 190080
rect 298698 174526 298934 174762
rect 298698 159208 298934 159444
rect 298698 143890 298934 144126
rect 298698 128572 298934 128808
rect 298698 113254 298934 113490
rect 298698 97936 298934 98172
rect 298698 82618 298934 82854
rect 298698 67300 298934 67536
rect 298698 51982 298934 52218
rect 298698 36664 298934 36900
rect 298698 21346 298934 21582
rect 298698 6028 298934 6264
rect 298698 2218 298934 2454
rect 298698 1898 298934 2134
rect 299638 289411 299874 289647
rect 299638 274093 299874 274329
rect 299638 258775 299874 259011
rect 299638 243457 299874 243693
rect 299638 228139 299874 228375
rect 299638 212821 299874 213057
rect 299638 197503 299874 197739
rect 299638 182185 299874 182421
rect 299638 166867 299874 167103
rect 299638 151549 299874 151785
rect 299638 136231 299874 136467
rect 299638 120913 299874 121149
rect 299638 105595 299874 105831
rect 299638 90277 299874 90513
rect 299638 74959 299874 75195
rect 299638 59641 299874 59877
rect 299638 44323 299874 44559
rect 299638 29005 299874 29241
rect 299638 13687 299874 13923
rect 46 958 282 1194
rect 20250 1278 20486 1340
rect 20250 958 20486 1194
rect 50970 1278 51206 1340
rect 50970 958 51206 1194
rect 81690 1278 81926 1340
rect 81690 958 81926 1194
rect 112410 1278 112646 1340
rect 112410 958 112646 1194
rect 143130 1278 143366 1340
rect 143130 958 143366 1194
rect 173850 1278 174086 1340
rect 173850 958 174086 1194
rect 204570 1278 204806 1340
rect 204570 958 204806 1194
rect 235290 1278 235526 1340
rect 235290 958 235526 1194
rect 266010 1278 266246 1340
rect 266010 958 266246 1194
rect 296730 1278 296966 1340
rect 296730 958 296966 1194
rect 299638 1278 299874 1514
rect 299638 958 299874 1194
<< metal5 >>
rect -136 298808 464 298810
rect 20208 298808 20528 298810
rect 50928 298808 51248 298810
rect 81648 298808 81968 298810
rect 112368 298808 112688 298810
rect 143088 298808 143408 298810
rect 173808 298808 174128 298810
rect 204528 298808 204848 298810
rect 235248 298808 235568 298810
rect 265968 298808 266288 298810
rect 296688 298808 297008 298810
rect 299456 298808 300056 298810
rect -136 298786 300056 298808
rect -136 298550 46 298786
rect 282 298660 20250 298786
rect 20486 298660 50970 298786
rect 51206 298660 81690 298786
rect 81926 298660 112410 298786
rect 112646 298660 143130 298786
rect 143366 298660 173850 298786
rect 174086 298660 204570 298786
rect 204806 298660 235290 298786
rect 235526 298660 266010 298786
rect 266246 298660 296730 298786
rect 296966 298660 299638 298786
rect 282 298550 1340 298660
rect -136 298466 1340 298550
rect -136 298230 46 298466
rect 282 298230 1340 298466
rect -136 298208 1340 298230
rect -136 298206 464 298208
rect 804 297846 1340 297870
rect 804 297610 986 297846
rect 1222 297610 1340 297846
rect 804 297526 1340 297610
rect 804 297290 986 297526
rect 1222 297290 1340 297526
rect 804 297266 1340 297290
rect -136 289647 1340 289689
rect -136 289411 46 289647
rect 282 289411 1340 289647
rect -136 289369 1340 289411
rect -136 281988 1340 282030
rect -136 281752 986 281988
rect 1222 281752 1340 281988
rect -136 281710 1340 281752
rect -136 274329 1340 274371
rect -136 274093 46 274329
rect 282 274093 1340 274329
rect -136 274051 1340 274093
rect -136 266670 1340 266712
rect -136 266434 986 266670
rect 1222 266434 1340 266670
rect -136 266392 1340 266434
rect -136 259011 1340 259053
rect -136 258775 46 259011
rect 282 258775 1340 259011
rect -136 258733 1340 258775
rect -136 251352 1340 251394
rect -136 251116 986 251352
rect 1222 251116 1340 251352
rect -136 251074 1340 251116
rect -136 243693 1340 243735
rect -136 243457 46 243693
rect 282 243457 1340 243693
rect -136 243415 1340 243457
rect -136 236034 1340 236076
rect -136 235798 986 236034
rect 1222 235798 1340 236034
rect -136 235756 1340 235798
rect -136 228375 1340 228417
rect -136 228139 46 228375
rect 282 228139 1340 228375
rect -136 228097 1340 228139
rect -136 220716 1340 220758
rect -136 220480 986 220716
rect 1222 220480 1340 220716
rect -136 220438 1340 220480
rect -136 213057 1340 213099
rect -136 212821 46 213057
rect 282 212821 1340 213057
rect -136 212779 1340 212821
rect -136 205398 1340 205440
rect -136 205162 986 205398
rect 1222 205162 1340 205398
rect -136 205120 1340 205162
rect -136 197739 1340 197781
rect -136 197503 46 197739
rect 282 197503 1340 197739
rect -136 197461 1340 197503
rect -136 190080 1340 190122
rect -136 189844 986 190080
rect 1222 189844 1340 190080
rect -136 189802 1340 189844
rect -136 182421 1340 182463
rect -136 182185 46 182421
rect 282 182185 1340 182421
rect -136 182143 1340 182185
rect -136 174762 1340 174804
rect -136 174526 986 174762
rect 1222 174526 1340 174762
rect -136 174484 1340 174526
rect -136 167103 1340 167145
rect -136 166867 46 167103
rect 282 166867 1340 167103
rect -136 166825 1340 166867
rect -136 159444 1340 159486
rect -136 159208 986 159444
rect 1222 159208 1340 159444
rect -136 159166 1340 159208
rect -136 151785 1340 151827
rect -136 151549 46 151785
rect 282 151549 1340 151785
rect -136 151507 1340 151549
rect -136 144126 1340 144168
rect -136 143890 986 144126
rect 1222 143890 1340 144126
rect -136 143848 1340 143890
rect -136 136467 1340 136509
rect -136 136231 46 136467
rect 282 136231 1340 136467
rect -136 136189 1340 136231
rect -136 128808 1340 128850
rect -136 128572 986 128808
rect 1222 128572 1340 128808
rect -136 128530 1340 128572
rect -136 121149 1340 121191
rect -136 120913 46 121149
rect 282 120913 1340 121149
rect -136 120871 1340 120913
rect -136 113490 1340 113532
rect -136 113254 986 113490
rect 1222 113254 1340 113490
rect -136 113212 1340 113254
rect -136 105831 1340 105873
rect -136 105595 46 105831
rect 282 105595 1340 105831
rect -136 105553 1340 105595
rect -136 98172 1340 98214
rect -136 97936 986 98172
rect 1222 97936 1340 98172
rect -136 97894 1340 97936
rect -136 90513 1340 90555
rect -136 90277 46 90513
rect 282 90277 1340 90513
rect -136 90235 1340 90277
rect -136 82854 1340 82896
rect -136 82618 986 82854
rect 1222 82618 1340 82854
rect -136 82576 1340 82618
rect -136 75195 1340 75237
rect -136 74959 46 75195
rect 282 74959 1340 75195
rect -136 74917 1340 74959
rect -136 67536 1340 67578
rect -136 67300 986 67536
rect 1222 67300 1340 67536
rect -136 67258 1340 67300
rect -136 59877 1340 59919
rect -136 59641 46 59877
rect 282 59641 1340 59877
rect -136 59599 1340 59641
rect -136 52218 1340 52260
rect -136 51982 986 52218
rect 1222 51982 1340 52218
rect -136 51940 1340 51982
rect -136 44559 1340 44601
rect -136 44323 46 44559
rect 282 44323 1340 44559
rect -136 44281 1340 44323
rect -136 36900 1340 36942
rect -136 36664 986 36900
rect 1222 36664 1340 36900
rect -136 36622 1340 36664
rect -136 29241 1340 29283
rect -136 29005 46 29241
rect 282 29005 1340 29241
rect -136 28963 1340 29005
rect -136 21582 1340 21624
rect -136 21346 986 21582
rect 1222 21346 1340 21582
rect -136 21304 1340 21346
rect -136 13923 1340 13965
rect -136 13687 46 13923
rect 282 13687 1340 13923
rect -136 13645 1340 13687
rect -136 6264 1340 6306
rect -136 6028 986 6264
rect 1222 6028 1340 6264
rect -136 5986 1340 6028
rect 804 2454 1340 2478
rect 804 2218 986 2454
rect 1222 2218 1340 2454
rect 804 2134 1340 2218
rect 804 1898 986 2134
rect 1222 1898 1340 2134
rect 804 1874 1340 1898
rect -136 1536 464 1538
rect -136 1514 1340 1536
rect -136 1278 46 1514
rect 282 1340 1340 1514
rect 298660 298550 299638 298660
rect 299874 298550 300056 298786
rect 298660 298466 300056 298550
rect 298660 298230 299638 298466
rect 299874 298230 300056 298466
rect 298660 298208 300056 298230
rect 299456 298206 300056 298208
rect 298660 297846 299116 297870
rect 298660 297610 298698 297846
rect 298934 297610 299116 297846
rect 298660 297526 299116 297610
rect 298660 297290 298698 297526
rect 298934 297290 299116 297526
rect 298660 297266 299116 297290
rect 298660 289647 300056 289689
rect 298660 289411 299638 289647
rect 299874 289411 300056 289647
rect 298660 289369 300056 289411
rect 298660 281988 300056 282030
rect 298660 281752 298698 281988
rect 298934 281752 300056 281988
rect 298660 281710 300056 281752
rect 298660 274329 300056 274371
rect 298660 274093 299638 274329
rect 299874 274093 300056 274329
rect 298660 274051 300056 274093
rect 298660 266670 300056 266712
rect 298660 266434 298698 266670
rect 298934 266434 300056 266670
rect 298660 266392 300056 266434
rect 298660 259011 300056 259053
rect 298660 258775 299638 259011
rect 299874 258775 300056 259011
rect 298660 258733 300056 258775
rect 298660 251352 300056 251394
rect 298660 251116 298698 251352
rect 298934 251116 300056 251352
rect 298660 251074 300056 251116
rect 298660 243693 300056 243735
rect 298660 243457 299638 243693
rect 299874 243457 300056 243693
rect 298660 243415 300056 243457
rect 298660 236034 300056 236076
rect 298660 235798 298698 236034
rect 298934 235798 300056 236034
rect 298660 235756 300056 235798
rect 298660 228375 300056 228417
rect 298660 228139 299638 228375
rect 299874 228139 300056 228375
rect 298660 228097 300056 228139
rect 298660 220716 300056 220758
rect 298660 220480 298698 220716
rect 298934 220480 300056 220716
rect 298660 220438 300056 220480
rect 298660 213057 300056 213099
rect 298660 212821 299638 213057
rect 299874 212821 300056 213057
rect 298660 212779 300056 212821
rect 298660 205398 300056 205440
rect 298660 205162 298698 205398
rect 298934 205162 300056 205398
rect 298660 205120 300056 205162
rect 298660 197739 300056 197781
rect 298660 197503 299638 197739
rect 299874 197503 300056 197739
rect 298660 197461 300056 197503
rect 298660 190080 300056 190122
rect 298660 189844 298698 190080
rect 298934 189844 300056 190080
rect 298660 189802 300056 189844
rect 298660 182421 300056 182463
rect 298660 182185 299638 182421
rect 299874 182185 300056 182421
rect 298660 182143 300056 182185
rect 298660 174762 300056 174804
rect 298660 174526 298698 174762
rect 298934 174526 300056 174762
rect 298660 174484 300056 174526
rect 298660 167103 300056 167145
rect 298660 166867 299638 167103
rect 299874 166867 300056 167103
rect 298660 166825 300056 166867
rect 298660 159444 300056 159486
rect 298660 159208 298698 159444
rect 298934 159208 300056 159444
rect 298660 159166 300056 159208
rect 298660 151785 300056 151827
rect 298660 151549 299638 151785
rect 299874 151549 300056 151785
rect 298660 151507 300056 151549
rect 298660 144126 300056 144168
rect 298660 143890 298698 144126
rect 298934 143890 300056 144126
rect 298660 143848 300056 143890
rect 298660 136467 300056 136509
rect 298660 136231 299638 136467
rect 299874 136231 300056 136467
rect 298660 136189 300056 136231
rect 298660 128808 300056 128850
rect 298660 128572 298698 128808
rect 298934 128572 300056 128808
rect 298660 128530 300056 128572
rect 298660 121149 300056 121191
rect 298660 120913 299638 121149
rect 299874 120913 300056 121149
rect 298660 120871 300056 120913
rect 298660 113490 300056 113532
rect 298660 113254 298698 113490
rect 298934 113254 300056 113490
rect 298660 113212 300056 113254
rect 298660 105831 300056 105873
rect 298660 105595 299638 105831
rect 299874 105595 300056 105831
rect 298660 105553 300056 105595
rect 298660 98172 300056 98214
rect 298660 97936 298698 98172
rect 298934 97936 300056 98172
rect 298660 97894 300056 97936
rect 298660 90513 300056 90555
rect 298660 90277 299638 90513
rect 299874 90277 300056 90513
rect 298660 90235 300056 90277
rect 298660 82854 300056 82896
rect 298660 82618 298698 82854
rect 298934 82618 300056 82854
rect 298660 82576 300056 82618
rect 298660 75195 300056 75237
rect 298660 74959 299638 75195
rect 299874 74959 300056 75195
rect 298660 74917 300056 74959
rect 298660 67536 300056 67578
rect 298660 67300 298698 67536
rect 298934 67300 300056 67536
rect 298660 67258 300056 67300
rect 298660 59877 300056 59919
rect 298660 59641 299638 59877
rect 299874 59641 300056 59877
rect 298660 59599 300056 59641
rect 298660 52218 300056 52260
rect 298660 51982 298698 52218
rect 298934 51982 300056 52218
rect 298660 51940 300056 51982
rect 298660 44559 300056 44601
rect 298660 44323 299638 44559
rect 299874 44323 300056 44559
rect 298660 44281 300056 44323
rect 298660 36900 300056 36942
rect 298660 36664 298698 36900
rect 298934 36664 300056 36900
rect 298660 36622 300056 36664
rect 298660 29241 300056 29283
rect 298660 29005 299638 29241
rect 299874 29005 300056 29241
rect 298660 28963 300056 29005
rect 298660 21582 300056 21624
rect 298660 21346 298698 21582
rect 298934 21346 300056 21582
rect 298660 21304 300056 21346
rect 298660 13923 300056 13965
rect 298660 13687 299638 13923
rect 299874 13687 300056 13923
rect 298660 13645 300056 13687
rect 298660 6264 300056 6306
rect 298660 6028 298698 6264
rect 298934 6028 300056 6264
rect 298660 5986 300056 6028
rect 298660 2454 299116 2478
rect 298660 2218 298698 2454
rect 298934 2218 299116 2454
rect 298660 2134 299116 2218
rect 298660 1898 298698 2134
rect 298934 1898 299116 2134
rect 298660 1874 299116 1898
rect 299456 1536 300056 1538
rect 298660 1514 300056 1536
rect 298660 1340 299638 1514
rect 282 1278 20250 1340
rect 20486 1278 50970 1340
rect 51206 1278 81690 1340
rect 81926 1278 112410 1340
rect 112646 1278 143130 1340
rect 143366 1278 173850 1340
rect 174086 1278 204570 1340
rect 204806 1278 235290 1340
rect 235526 1278 266010 1340
rect 266246 1278 296730 1340
rect 296966 1278 299638 1340
rect 299874 1278 300056 1514
rect -136 1194 300056 1278
rect -136 958 46 1194
rect 282 958 20250 1194
rect 20486 958 50970 1194
rect 51206 958 81690 1194
rect 81926 958 112410 1194
rect 112646 958 143130 1194
rect 143366 958 173850 1194
rect 174086 958 204570 1194
rect 204806 958 235290 1194
rect 235526 958 266010 1194
rect 266246 958 296730 1194
rect 296966 958 299638 1194
rect 299874 958 300056 1194
rect -136 936 300056 958
rect -136 934 464 936
rect 20208 934 20528 936
rect 50928 934 51248 936
rect 81648 934 81968 936
rect 112368 934 112688 936
rect 143088 934 143408 936
rect 173808 934 174128 936
rect 204528 934 204848 936
rect 235248 934 235568 936
rect 265968 934 266288 936
rect 296688 934 297008 936
rect 299456 934 300056 936
<< obsm5 >>
rect 1340 1340 298660 298660
<< labels >>
rlabel metal2 s 1278 299400 1390 301200 6 io_in[0]
port 1 nsew default input
rlabel metal2 s 79478 299400 79590 301200 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 87298 299400 87410 301200 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 95118 299400 95230 301200 6 io_in[12]
port 4 nsew default input
rlabel metal2 s 102938 299400 103050 301200 6 io_in[13]
port 5 nsew default input
rlabel metal2 s 110758 299400 110870 301200 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 118670 299400 118782 301200 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 126490 299400 126602 301200 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 134310 299400 134422 301200 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 142130 299400 142242 301200 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 149950 299400 150062 301200 6 io_in[19]
port 11 nsew default input
rlabel metal2 s 9098 299400 9210 301200 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 157770 299400 157882 301200 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 165590 299400 165702 301200 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 173410 299400 173522 301200 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 181230 299400 181342 301200 6 io_in[23]
port 16 nsew default input
rlabel metal2 s 189050 299400 189162 301200 6 io_in[24]
port 17 nsew default input
rlabel metal2 s 196870 299400 196982 301200 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 204690 299400 204802 301200 6 io_in[26]
port 19 nsew default input
rlabel metal2 s 212510 299400 212622 301200 6 io_in[27]
port 20 nsew default input
rlabel metal2 s 220330 299400 220442 301200 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 228242 299400 228354 301200 6 io_in[29]
port 22 nsew default input
rlabel metal2 s 16918 299400 17030 301200 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 236062 299400 236174 301200 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 243882 299400 243994 301200 6 io_in[31]
port 25 nsew default input
rlabel metal2 s 251702 299400 251814 301200 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 259522 299400 259634 301200 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 267342 299400 267454 301200 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 275162 299400 275274 301200 6 io_in[35]
port 29 nsew default input
rlabel metal2 s 282982 299400 283094 301200 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 290802 299400 290914 301200 6 io_in[37]
port 31 nsew default input
rlabel metal2 s 24738 299400 24850 301200 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 32558 299400 32670 301200 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 40378 299400 40490 301200 6 io_in[5]
port 34 nsew default input
rlabel metal2 s 48198 299400 48310 301200 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 56018 299400 56130 301200 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 63838 299400 63950 301200 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 71658 299400 71770 301200 6 io_in[9]
port 38 nsew default input
rlabel metal2 s 3896 298660 3924 299400 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 3854 299400 3966 301200 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 82188 298660 82216 299400 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 82146 299400 82258 301200 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 90008 298660 90036 299400 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 89966 299400 90078 301200 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 97828 298660 97856 299400 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 97786 299400 97898 301200 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 105648 298660 105676 299400 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 105606 299400 105718 301200 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 113468 298660 113496 299400 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 113426 299400 113538 301200 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 121288 298660 121316 299400 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 121246 299400 121358 301200 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 129108 298660 129136 299400 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 129066 299400 129178 301200 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 136928 298660 136956 299400 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 136886 299400 136998 301200 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 144748 298660 144776 299400 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 144706 299400 144818 301200 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 152568 298660 152596 299400 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 152526 299400 152638 301200 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 11716 298660 11744 299400 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 11674 299400 11786 301200 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 160388 298660 160416 299400 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 160346 299400 160458 301200 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 168208 298660 168236 299400 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 168166 299400 168278 301200 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 176028 298660 176056 299400 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 175986 299400 176098 301200 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 183848 298660 183876 299400 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 183806 299400 183918 301200 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 191760 298660 191788 299400 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 191718 299400 191830 301200 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 199580 298660 199608 299400 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 199538 299400 199650 301200 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 207400 298660 207428 299400 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 207358 299400 207470 301200 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 215220 298660 215248 299400 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 215178 299400 215290 301200 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 223040 298660 223068 299400 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 222998 299400 223110 301200 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 230860 298660 230888 299400 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 230818 299400 230930 301200 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 19536 298660 19564 299400 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 19494 299400 19606 301200 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 238680 298660 238708 299400 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 238638 299400 238750 301200 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 246500 298660 246528 299400 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 246458 299400 246570 301200 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 254320 298660 254348 299400 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 254278 299400 254390 301200 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 262140 298660 262168 299400 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 262098 299400 262210 301200 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 269960 298660 269988 299400 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 269918 299400 270030 301200 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 277780 298660 277808 299400 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 277738 299400 277850 301200 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 285600 298660 285628 299400 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 285558 299400 285670 301200 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 293420 298660 293448 299400 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 293378 299400 293490 301200 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 27356 298660 27384 299400 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 27314 299400 27426 301200 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 35176 298660 35204 299400 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 35134 299400 35246 301200 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 42996 298660 43024 299400 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 42954 299400 43066 301200 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 50816 298660 50844 299400 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 50774 299400 50886 301200 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 58636 298660 58664 299400 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 58594 299400 58706 301200 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 66456 298660 66484 299400 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 66414 299400 66526 301200 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 74276 298660 74304 299400 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 74234 299400 74346 301200 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 6472 298660 6500 299400 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 6430 299400 6542 301200 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 84764 298660 84792 299400 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 84722 299400 84834 301200 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 92584 298660 92612 299400 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 92542 299400 92654 301200 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 100404 298660 100432 299400 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 100362 299400 100474 301200 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 108224 298660 108252 299400 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 108182 299400 108294 301200 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 116044 298660 116072 299400 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 116002 299400 116114 301200 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 123864 298660 123892 299400 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 123822 299400 123934 301200 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 131684 298660 131712 299400 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 131642 299400 131754 301200 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 139504 298660 139532 299400 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 139462 299400 139574 301200 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 147324 298660 147352 299400 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 147282 299400 147394 301200 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 155236 298660 155264 299400 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 155194 299400 155306 301200 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 14292 298660 14320 299400 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 14250 299400 14362 301200 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 163056 298660 163084 299400 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 163014 299400 163126 301200 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 170876 298660 170904 299400 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 170834 299400 170946 301200 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 178696 298660 178724 299400 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 178654 299400 178766 301200 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 186516 298660 186544 299400 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 186474 299400 186586 301200 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 194336 298660 194364 299400 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 194294 299400 194406 301200 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 202156 298660 202184 299400 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 202114 299400 202226 301200 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 209976 298660 210004 299400 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 209934 299400 210046 301200 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 217796 298660 217824 299400 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 217754 299400 217866 301200 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 225616 298660 225644 299400 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 225574 299400 225686 301200 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 233436 298660 233464 299400 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 233394 299400 233506 301200 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 22112 298660 22140 299400 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 22070 299400 22182 301200 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 241256 298660 241284 299400 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 241214 299400 241326 301200 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 249076 298660 249104 299400 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 249034 299400 249146 301200 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 256896 298660 256924 299400 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 256854 299400 256966 301200 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 264808 298660 264836 299400 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 264766 299400 264878 301200 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 272628 298660 272656 299400 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 272586 299400 272698 301200 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 280448 298660 280476 299400 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 280406 299400 280518 301200 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 288268 298660 288296 299400 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 288226 299400 288338 301200 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 296088 298660 296116 299400 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 296046 299400 296158 301200 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 29932 298660 29960 299400 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 29890 299400 30002 301200 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 37752 298660 37780 299400 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 37710 299400 37822 301200 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 45664 298660 45692 299400 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 45622 299400 45734 301200 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 53484 298660 53512 299400 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 53442 299400 53554 301200 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 61304 298660 61332 299400 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 61262 299400 61374 301200 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 69124 298660 69152 299400 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 69082 299400 69194 301200 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 76944 298660 76972 299400 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 76902 299400 77014 301200 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 64850 -1200 64962 600 8 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 247746 -1200 247858 600 8 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 247788 600 247816 1340 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 249586 -1200 249698 600 8 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 249628 600 249656 1340 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 251426 -1200 251538 600 8 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 251468 600 251496 1340 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 253266 -1200 253378 600 8 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 253308 600 253336 1340 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 255106 -1200 255218 600 8 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 255148 600 255176 1340 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 256946 -1200 257058 600 8 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 256988 600 257016 1340 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 258786 -1200 258898 600 8 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 258828 600 258856 1340 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 260626 -1200 260738 600 8 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 260668 600 260696 1340 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 262466 -1200 262578 600 8 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 262508 600 262536 1340 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 264214 -1200 264326 600 8 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 264256 600 264284 1340 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 83158 -1200 83270 600 8 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 266054 -1200 266166 600 8 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 266096 600 266124 1340 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 267894 -1200 268006 600 8 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 267936 600 267964 1340 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 269734 -1200 269846 598 8 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 269684 598 269846 600 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 269684 600 269804 626 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 269684 626 269712 734 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 269132 734 269712 762 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 269132 762 269160 1340 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 271574 -1200 271686 598 8 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 271524 598 271686 600 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 271524 600 271644 626 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 271524 626 271552 1340 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 273414 -1200 273526 600 8 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 275254 -1200 275366 600 8 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 277094 -1200 277206 600 8 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 278934 -1200 279046 600 8 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 280682 -1200 280794 600 8 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 282522 -1200 282634 600 8 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 84998 -1200 85110 600 8 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 284362 -1200 284474 600 8 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 286202 -1200 286314 600 8 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 288042 -1200 288154 600 8 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 289882 -1200 289994 600 8 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 291722 -1200 291834 600 8 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 293562 -1200 293674 600 8 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 295310 -1200 295422 600 8 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 297150 -1200 297262 600 8 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 86838 -1200 86950 600 8 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 88678 -1200 88790 600 8 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 90426 -1200 90538 600 8 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 92266 -1200 92378 600 8 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 94106 -1200 94218 600 8 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 95946 -1200 96058 600 8 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 97786 -1200 97898 600 8 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 99626 -1200 99738 600 8 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 66690 -1200 66802 600 8 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 101466 -1200 101578 600 8 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 103306 -1200 103418 600 8 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 105146 -1200 105258 600 8 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 106894 -1200 107006 600 8 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 108734 -1200 108846 600 8 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 110574 -1200 110686 600 8 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 112414 -1200 112526 600 8 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 114254 -1200 114366 600 8 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 116094 -1200 116206 600 8 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 117934 -1200 118046 600 8 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 68530 -1200 68642 600 8 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 119774 -1200 119886 600 8 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 121522 -1200 121634 600 8 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 123362 -1200 123474 600 8 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 125202 -1200 125314 600 8 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 127042 -1200 127154 600 8 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 128882 -1200 128994 600 8 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 130722 -1200 130834 600 8 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 132562 -1200 132674 600 8 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 134402 -1200 134514 600 8 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 136242 -1200 136354 600 8 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 70370 -1200 70482 600 8 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 137990 -1200 138102 600 8 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 139830 -1200 139942 600 8 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 141670 -1200 141782 600 8 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 143510 -1200 143622 600 8 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 145350 -1200 145462 600 8 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 147190 -1200 147302 600 8 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 149030 -1200 149142 600 8 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 150870 -1200 150982 600 8 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 152710 -1200 152822 600 8 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 154458 -1200 154570 600 8 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 72210 -1200 72322 600 8 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 156298 -1200 156410 600 8 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 158138 -1200 158250 600 8 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 159978 -1200 160090 600 8 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 161818 -1200 161930 600 8 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 163658 -1200 163770 600 8 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 165498 -1200 165610 600 8 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 167338 -1200 167450 600 8 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 169086 -1200 169198 600 8 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 170926 -1200 171038 600 8 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 172766 -1200 172878 600 8 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 73958 -1200 74070 600 8 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 174606 -1200 174718 600 8 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 176446 -1200 176558 600 8 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 178286 -1200 178398 600 8 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 180126 -1200 180238 600 8 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 181966 -1200 182078 600 8 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 182008 600 182036 1340 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 183806 -1200 183918 600 8 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 183848 600 183876 1340 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 185554 -1200 185666 600 8 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 185596 600 185624 1340 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 187394 -1200 187506 600 8 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 187436 600 187464 1340 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 189234 -1200 189346 600 8 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 189276 600 189304 1340 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 191074 -1200 191186 600 8 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 191116 600 191144 1340 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 75798 -1200 75910 600 8 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 192914 -1200 193026 600 8 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 192956 600 192984 1340 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 194754 -1200 194866 600 8 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 194796 600 194824 1340 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 196594 -1200 196706 600 8 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 196636 600 196664 1340 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 198434 -1200 198546 600 8 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 198476 600 198504 1340 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 200274 -1200 200386 600 8 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 200316 600 200344 1340 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 202022 -1200 202134 600 8 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 202064 600 202092 1340 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 203862 -1200 203974 600 8 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 203904 600 203932 1340 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 205702 -1200 205814 600 8 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 205744 600 205772 1340 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 207542 -1200 207654 600 8 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 207584 600 207612 1340 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 209382 -1200 209494 600 8 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 209424 600 209452 1340 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 77638 -1200 77750 600 8 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 211222 -1200 211334 600 8 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 211264 600 211292 1340 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 213062 -1200 213174 600 8 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 213104 600 213132 1340 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 214902 -1200 215014 600 8 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 214944 600 214972 1340 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 216650 -1200 216762 600 8 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 216692 600 216720 1340 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 218490 -1200 218602 600 8 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 218532 600 218560 1340 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 220330 -1200 220442 600 8 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 220372 600 220400 1340 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 222170 -1200 222282 600 8 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 222212 600 222240 1340 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 224010 -1200 224122 600 8 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 224052 600 224080 1340 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 225850 -1200 225962 600 8 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 225892 600 225920 1340 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 227690 -1200 227802 600 8 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 227732 600 227760 1340 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 79478 -1200 79590 600 8 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 229530 -1200 229642 600 8 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 229572 600 229600 1340 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 231370 -1200 231482 600 8 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 231412 600 231440 1340 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 233118 -1200 233230 600 8 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 233160 600 233188 1340 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 234958 -1200 235070 600 8 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 235000 600 235028 1340 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 236798 -1200 236910 600 8 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 236840 600 236868 1340 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 238638 -1200 238750 600 8 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 238680 600 238708 1340 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 240478 -1200 240590 600 8 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 240520 600 240548 1340 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 242318 -1200 242430 600 8 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 242360 600 242388 1340 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 244158 -1200 244270 600 8 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 244200 600 244228 1340 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 245998 -1200 246110 600 8 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 246040 600 246068 1340 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 81318 -1200 81430 600 8 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 65494 -1200 65606 600 8 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 65536 600 65564 1340 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 248390 -1200 248502 600 8 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 248432 600 248460 1340 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 250230 -1200 250342 600 8 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 250272 600 250300 1340 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 252070 -1200 252182 600 8 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 252112 600 252140 1340 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 253910 -1200 254022 600 8 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 253952 600 253980 1340 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 255750 -1200 255862 600 8 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 255792 600 255820 1340 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 257590 -1200 257702 600 8 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 257632 600 257660 1340 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 259338 -1200 259450 600 8 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 259380 600 259408 1340 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 261178 -1200 261290 600 8 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 261220 600 261248 1340 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 263018 -1200 263130 600 8 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 263060 600 263088 1340 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 264858 -1200 264970 600 8 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 264900 600 264928 1340 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 83802 -1200 83914 598 8 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 83802 598 84148 600 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 83844 600 84148 626 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 84120 626 84148 1340 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 266698 -1200 266810 600 8 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 266740 600 266768 1340 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 268538 -1200 268650 600 8 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 268580 600 268608 1340 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 270378 -1200 270490 600 8 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 270420 600 270448 1340 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 272218 -1200 272330 600 8 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 272260 600 272288 1340 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 273966 -1200 274078 600 8 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 274008 600 274036 1340 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 275806 -1200 275918 600 8 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 275848 600 275876 1340 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 277646 -1200 277758 600 8 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 277688 600 277716 1340 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 279486 -1200 279598 600 8 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 279528 600 279556 1340 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 281326 -1200 281438 600 8 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 281368 600 281396 1340 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 283166 -1200 283278 600 8 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 283208 600 283236 1340 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 85550 -1200 85662 600 8 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 85592 600 85620 1340 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 285006 -1200 285118 600 8 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 285048 600 285076 1340 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 286846 -1200 286958 600 8 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 286888 600 286916 1340 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 288686 -1200 288798 600 8 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 288728 600 288756 1340 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 290434 -1200 290546 600 8 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 290476 600 290504 1340 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 292274 -1200 292386 600 8 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 292316 600 292344 1340 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 294114 -1200 294226 600 8 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 294156 600 294184 1340 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 295954 -1200 296066 600 8 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 295996 600 296024 1340 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 297794 -1200 297906 600 8 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 297836 600 297864 1340 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 87390 -1200 87502 600 8 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 87432 600 87460 1340 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 89230 -1200 89342 600 8 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 89272 600 89300 1340 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 91070 -1200 91182 600 8 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 91112 600 91140 1340 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 92910 -1200 93022 600 8 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 92952 600 92980 1340 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 94750 -1200 94862 600 8 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 94792 600 94820 1340 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 96590 -1200 96702 600 8 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 96632 600 96660 1340 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 98430 -1200 98542 600 8 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 98472 600 98500 1340 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 100270 -1200 100382 598 8 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 100270 598 100708 600 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 100312 600 100708 626 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 100680 626 100708 1340 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 67334 -1200 67446 600 8 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 67376 600 67404 1340 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 102018 -1200 102130 600 8 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 102060 600 102088 1340 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 103858 -1200 103970 600 8 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 103900 600 103928 1340 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 105698 -1200 105810 600 8 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 105740 600 105768 1340 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 107538 -1200 107650 600 8 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 107580 600 107608 1340 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 109378 -1200 109490 600 8 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 109420 600 109448 1340 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 111218 -1200 111330 600 8 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 111260 600 111288 1340 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 113058 -1200 113170 600 8 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 113100 600 113128 1340 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 114898 -1200 115010 600 8 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 114940 600 114968 1340 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 116646 -1200 116758 600 8 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 116688 600 116716 1340 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 118486 -1200 118598 600 8 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 118528 600 118556 1340 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 69082 -1200 69194 600 8 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 69124 600 69152 1340 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 120326 -1200 120438 600 8 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 120368 600 120396 1340 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 122166 -1200 122278 600 8 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 122208 600 122236 1340 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 124006 -1200 124118 600 8 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 124048 600 124076 1340 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 125846 -1200 125958 600 8 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 125888 600 125916 1340 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 127686 -1200 127798 600 8 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 127728 600 127756 1340 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 129526 -1200 129638 600 8 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 129568 600 129596 1340 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 131366 -1200 131478 600 8 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 131408 600 131436 1340 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 133114 -1200 133226 600 8 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 133156 600 133184 1340 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 134954 -1200 135066 600 8 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 134996 600 135024 1340 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 136794 -1200 136906 600 8 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 136836 600 136864 1340 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 70922 -1200 71034 600 8 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 70964 600 70992 1340 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 138634 -1200 138746 598 8 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 138634 598 138980 600 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 138676 600 138980 626 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 138952 626 138980 1340 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 140474 -1200 140586 600 8 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 140516 600 140544 1340 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 142314 -1200 142426 600 8 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 142356 600 142384 1340 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 144154 -1200 144266 600 8 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 144196 600 144224 1340 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 145994 -1200 146106 600 8 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 146036 600 146064 1340 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 147742 -1200 147854 600 8 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 147784 600 147812 1340 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 149582 -1200 149694 600 8 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 149624 600 149652 1340 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 151422 -1200 151534 600 8 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 151464 600 151492 1340 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 153262 -1200 153374 600 8 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 153304 600 153332 1340 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 155102 -1200 155214 600 8 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 155144 600 155172 1340 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 72762 -1200 72874 600 8 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 72804 600 72832 1340 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 156942 -1200 157054 600 8 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 156984 600 157012 1340 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 158782 -1200 158894 600 8 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 158824 600 158852 1340 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 160622 -1200 160734 600 8 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 160664 600 160692 1340 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 162462 -1200 162574 600 8 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 162504 600 162532 1340 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 164210 -1200 164322 600 8 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 164252 600 164280 1340 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 166050 -1200 166162 600 8 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 166092 600 166120 1340 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 167890 -1200 168002 600 8 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 167932 600 167960 1340 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 169730 -1200 169842 600 8 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 169772 600 169800 1340 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 171570 -1200 171682 600 8 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 171612 600 171640 1340 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 173410 -1200 173522 600 8 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 173452 600 173480 1340 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 74602 -1200 74714 600 8 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 74644 600 74672 1340 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 175250 -1200 175362 600 8 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 175292 600 175320 1340 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 177090 -1200 177202 600 8 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 177132 600 177160 1340 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 178930 -1200 179042 600 8 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 178972 600 179000 1340 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 180678 -1200 180790 600 8 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 180720 600 180748 1340 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 182518 -1200 182630 600 8 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 182560 600 182588 1340 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 184358 -1200 184470 600 8 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 184400 600 184428 1340 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 186198 -1200 186310 600 8 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 186240 600 186268 1340 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 188038 -1200 188150 600 8 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 188080 600 188108 1340 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 189878 -1200 189990 600 8 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 189920 600 189948 1340 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 191718 -1200 191830 600 8 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 191760 600 191788 1340 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 76442 -1200 76554 600 8 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 76484 600 76512 1340 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 193558 -1200 193670 600 8 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 193600 600 193628 1340 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 195306 -1200 195418 600 8 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 195348 600 195376 1340 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 197146 -1200 197258 600 8 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 197188 600 197216 1340 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 198986 -1200 199098 600 8 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 199028 600 199056 1340 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 200826 -1200 200938 600 8 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 200868 600 200896 1340 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 202666 -1200 202778 600 8 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 202708 600 202736 1340 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 204506 -1200 204618 600 8 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 204548 600 204576 1340 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 206346 -1200 206458 600 8 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 206388 600 206416 1340 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 208186 -1200 208298 600 8 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 208228 600 208256 1340 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 210026 -1200 210138 600 8 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 210068 600 210096 1340 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 78282 -1200 78394 598 8 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 78282 598 78628 600 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 78324 600 78628 626 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 78600 626 78628 1340 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 211774 -1200 211886 600 8 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 211816 600 211844 1340 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 213614 -1200 213726 600 8 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 213656 600 213684 1340 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 215454 -1200 215566 600 8 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 215496 600 215524 1340 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 217294 -1200 217406 600 8 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 217336 600 217364 1340 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 219134 -1200 219246 600 8 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 219176 600 219204 1340 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 220974 -1200 221086 600 8 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 221016 600 221044 1340 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 222814 -1200 222926 600 8 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 222856 600 222884 1340 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 224654 -1200 224766 600 8 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 224696 600 224724 1340 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 226494 -1200 226606 600 8 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 226536 600 226564 1340 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 228242 -1200 228354 600 8 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 228284 600 228312 1340 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 80122 -1200 80234 600 8 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 80164 600 80192 1340 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 230082 -1200 230194 600 8 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 230124 600 230152 1340 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 231922 -1200 232034 600 8 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 231964 600 231992 1340 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 233762 -1200 233874 600 8 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 233804 600 233832 1340 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 235602 -1200 235714 600 8 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 235644 600 235672 1340 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 237442 -1200 237554 600 8 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 237484 600 237512 1340 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 239282 -1200 239394 600 8 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 239324 600 239352 1340 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 241122 -1200 241234 600 8 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 241164 600 241192 1340 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 242870 -1200 242982 600 8 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 242912 600 242940 1340 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 244710 -1200 244822 600 8 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 244752 600 244780 1340 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 246550 -1200 246662 600 8 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 246592 600 246620 1340 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 81962 -1200 82074 600 8 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 82004 600 82032 1340 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 66046 -1200 66158 600 8 la_oen[0]
port 371 nsew default input
rlabel metal2 s 249034 -1200 249146 600 8 la_oen[100]
port 372 nsew default input
rlabel metal2 s 250874 -1200 250986 600 8 la_oen[101]
port 373 nsew default input
rlabel metal2 s 252714 -1200 252826 600 8 la_oen[102]
port 374 nsew default input
rlabel metal2 s 254462 -1200 254574 600 8 la_oen[103]
port 375 nsew default input
rlabel metal2 s 256302 -1200 256414 600 8 la_oen[104]
port 376 nsew default input
rlabel metal2 s 258142 -1200 258254 600 8 la_oen[105]
port 377 nsew default input
rlabel metal2 s 259982 -1200 260094 600 8 la_oen[106]
port 378 nsew default input
rlabel metal2 s 261822 -1200 261934 600 8 la_oen[107]
port 379 nsew default input
rlabel metal2 s 263662 -1200 263774 600 8 la_oen[108]
port 380 nsew default input
rlabel metal2 s 265502 -1200 265614 600 8 la_oen[109]
port 381 nsew default input
rlabel metal2 s 84354 -1200 84466 600 8 la_oen[10]
port 382 nsew default input
rlabel metal2 s 267342 -1200 267454 600 8 la_oen[110]
port 383 nsew default input
rlabel metal2 s 269090 -1200 269202 600 8 la_oen[111]
port 384 nsew default input
rlabel metal2 s 270930 -1200 271042 600 8 la_oen[112]
port 385 nsew default input
rlabel metal2 s 272770 -1200 272882 600 8 la_oen[113]
port 386 nsew default input
rlabel metal2 s 274610 -1200 274722 600 8 la_oen[114]
port 387 nsew default input
rlabel metal2 s 276450 -1200 276562 600 8 la_oen[115]
port 388 nsew default input
rlabel metal2 s 278290 -1200 278402 600 8 la_oen[116]
port 389 nsew default input
rlabel metal2 s 280130 -1200 280242 600 8 la_oen[117]
port 390 nsew default input
rlabel metal2 s 281970 -1200 282082 600 8 la_oen[118]
port 391 nsew default input
rlabel metal2 s 283810 -1200 283922 600 8 la_oen[119]
port 392 nsew default input
rlabel metal2 s 86194 -1200 86306 600 8 la_oen[11]
port 393 nsew default input
rlabel metal2 s 285558 -1200 285670 600 8 la_oen[120]
port 394 nsew default input
rlabel metal2 s 287398 -1200 287510 600 8 la_oen[121]
port 395 nsew default input
rlabel metal2 s 289238 -1200 289350 600 8 la_oen[122]
port 396 nsew default input
rlabel metal2 s 291078 -1200 291190 600 8 la_oen[123]
port 397 nsew default input
rlabel metal2 s 292918 -1200 293030 600 8 la_oen[124]
port 398 nsew default input
rlabel metal2 s 294758 -1200 294870 600 8 la_oen[125]
port 399 nsew default input
rlabel metal2 s 296598 -1200 296710 600 8 la_oen[126]
port 400 nsew default input
rlabel metal2 s 298438 -1200 298550 600 8 la_oen[127]
port 401 nsew default input
rlabel metal2 s 88034 -1200 88146 600 8 la_oen[12]
port 402 nsew default input
rlabel metal2 s 89874 -1200 89986 600 8 la_oen[13]
port 403 nsew default input
rlabel metal2 s 91714 -1200 91826 600 8 la_oen[14]
port 404 nsew default input
rlabel metal2 s 93554 -1200 93666 600 8 la_oen[15]
port 405 nsew default input
rlabel metal2 s 95302 -1200 95414 600 8 la_oen[16]
port 406 nsew default input
rlabel metal2 s 97142 -1200 97254 600 8 la_oen[17]
port 407 nsew default input
rlabel metal2 s 98982 -1200 99094 600 8 la_oen[18]
port 408 nsew default input
rlabel metal2 s 100822 -1200 100934 600 8 la_oen[19]
port 409 nsew default input
rlabel metal2 s 67886 -1200 67998 600 8 la_oen[1]
port 410 nsew default input
rlabel metal2 s 102662 -1200 102774 600 8 la_oen[20]
port 411 nsew default input
rlabel metal2 s 104502 -1200 104614 600 8 la_oen[21]
port 412 nsew default input
rlabel metal2 s 106342 -1200 106454 600 8 la_oen[22]
port 413 nsew default input
rlabel metal2 s 108182 -1200 108294 600 8 la_oen[23]
port 414 nsew default input
rlabel metal2 s 110022 -1200 110134 600 8 la_oen[24]
port 415 nsew default input
rlabel metal2 s 111770 -1200 111882 600 8 la_oen[25]
port 416 nsew default input
rlabel metal2 s 113610 -1200 113722 600 8 la_oen[26]
port 417 nsew default input
rlabel metal2 s 115450 -1200 115562 600 8 la_oen[27]
port 418 nsew default input
rlabel metal2 s 117290 -1200 117402 600 8 la_oen[28]
port 419 nsew default input
rlabel metal2 s 119130 -1200 119242 600 8 la_oen[29]
port 420 nsew default input
rlabel metal2 s 69726 -1200 69838 600 8 la_oen[2]
port 421 nsew default input
rlabel metal2 s 120970 -1200 121082 600 8 la_oen[30]
port 422 nsew default input
rlabel metal2 s 122810 -1200 122922 600 8 la_oen[31]
port 423 nsew default input
rlabel metal2 s 124650 -1200 124762 600 8 la_oen[32]
port 424 nsew default input
rlabel metal2 s 126490 -1200 126602 600 8 la_oen[33]
port 425 nsew default input
rlabel metal2 s 128238 -1200 128350 600 8 la_oen[34]
port 426 nsew default input
rlabel metal2 s 130078 -1200 130190 600 8 la_oen[35]
port 427 nsew default input
rlabel metal2 s 131918 -1200 132030 600 8 la_oen[36]
port 428 nsew default input
rlabel metal2 s 133758 -1200 133870 600 8 la_oen[37]
port 429 nsew default input
rlabel metal2 s 135598 -1200 135710 600 8 la_oen[38]
port 430 nsew default input
rlabel metal2 s 137438 -1200 137550 600 8 la_oen[39]
port 431 nsew default input
rlabel metal2 s 71566 -1200 71678 600 8 la_oen[3]
port 432 nsew default input
rlabel metal2 s 139278 -1200 139390 600 8 la_oen[40]
port 433 nsew default input
rlabel metal2 s 141118 -1200 141230 600 8 la_oen[41]
port 434 nsew default input
rlabel metal2 s 142866 -1200 142978 600 8 la_oen[42]
port 435 nsew default input
rlabel metal2 s 144706 -1200 144818 600 8 la_oen[43]
port 436 nsew default input
rlabel metal2 s 146546 -1200 146658 600 8 la_oen[44]
port 437 nsew default input
rlabel metal2 s 148386 -1200 148498 600 8 la_oen[45]
port 438 nsew default input
rlabel metal2 s 150226 -1200 150338 600 8 la_oen[46]
port 439 nsew default input
rlabel metal2 s 152066 -1200 152178 600 8 la_oen[47]
port 440 nsew default input
rlabel metal2 s 153906 -1200 154018 600 8 la_oen[48]
port 441 nsew default input
rlabel metal2 s 155746 -1200 155858 600 8 la_oen[49]
port 442 nsew default input
rlabel metal2 s 73406 -1200 73518 600 8 la_oen[4]
port 443 nsew default input
rlabel metal2 s 157586 -1200 157698 600 8 la_oen[50]
port 444 nsew default input
rlabel metal2 s 159334 -1200 159446 600 8 la_oen[51]
port 445 nsew default input
rlabel metal2 s 161174 -1200 161286 600 8 la_oen[52]
port 446 nsew default input
rlabel metal2 s 163014 -1200 163126 600 8 la_oen[53]
port 447 nsew default input
rlabel metal2 s 164854 -1200 164966 600 8 la_oen[54]
port 448 nsew default input
rlabel metal2 s 166694 -1200 166806 600 8 la_oen[55]
port 449 nsew default input
rlabel metal2 s 168534 -1200 168646 600 8 la_oen[56]
port 450 nsew default input
rlabel metal2 s 170374 -1200 170486 600 8 la_oen[57]
port 451 nsew default input
rlabel metal2 s 172214 -1200 172326 600 8 la_oen[58]
port 452 nsew default input
rlabel metal2 s 173962 -1200 174074 600 8 la_oen[59]
port 453 nsew default input
rlabel metal2 s 75246 -1200 75358 600 8 la_oen[5]
port 454 nsew default input
rlabel metal2 s 175802 -1200 175914 600 8 la_oen[60]
port 455 nsew default input
rlabel metal2 s 177642 -1200 177754 600 8 la_oen[61]
port 456 nsew default input
rlabel metal2 s 179482 -1200 179594 600 8 la_oen[62]
port 457 nsew default input
rlabel metal2 s 181322 -1200 181434 600 8 la_oen[63]
port 458 nsew default input
rlabel metal2 s 183162 -1200 183274 600 8 la_oen[64]
port 459 nsew default input
rlabel metal2 s 185002 -1200 185114 600 8 la_oen[65]
port 460 nsew default input
rlabel metal2 s 186842 -1200 186954 600 8 la_oen[66]
port 461 nsew default input
rlabel metal2 s 188682 -1200 188794 600 8 la_oen[67]
port 462 nsew default input
rlabel metal2 s 190430 -1200 190542 600 8 la_oen[68]
port 463 nsew default input
rlabel metal2 s 192270 -1200 192382 600 8 la_oen[69]
port 464 nsew default input
rlabel metal2 s 77086 -1200 77198 600 8 la_oen[6]
port 465 nsew default input
rlabel metal2 s 194110 -1200 194222 600 8 la_oen[70]
port 466 nsew default input
rlabel metal2 s 195950 -1200 196062 600 8 la_oen[71]
port 467 nsew default input
rlabel metal2 s 197790 -1200 197902 600 8 la_oen[72]
port 468 nsew default input
rlabel metal2 s 199630 -1200 199742 600 8 la_oen[73]
port 469 nsew default input
rlabel metal2 s 201470 -1200 201582 600 8 la_oen[74]
port 470 nsew default input
rlabel metal2 s 203310 -1200 203422 600 8 la_oen[75]
port 471 nsew default input
rlabel metal2 s 205150 -1200 205262 600 8 la_oen[76]
port 472 nsew default input
rlabel metal2 s 206898 -1200 207010 600 8 la_oen[77]
port 473 nsew default input
rlabel metal2 s 208738 -1200 208850 600 8 la_oen[78]
port 474 nsew default input
rlabel metal2 s 210578 -1200 210690 600 8 la_oen[79]
port 475 nsew default input
rlabel metal2 s 78926 -1200 79038 600 8 la_oen[7]
port 476 nsew default input
rlabel metal2 s 212418 -1200 212530 600 8 la_oen[80]
port 477 nsew default input
rlabel metal2 s 214258 -1200 214370 600 8 la_oen[81]
port 478 nsew default input
rlabel metal2 s 216098 -1200 216210 600 8 la_oen[82]
port 479 nsew default input
rlabel metal2 s 217938 -1200 218050 600 8 la_oen[83]
port 480 nsew default input
rlabel metal2 s 219778 -1200 219890 600 8 la_oen[84]
port 481 nsew default input
rlabel metal2 s 221526 -1200 221638 600 8 la_oen[85]
port 482 nsew default input
rlabel metal2 s 223366 -1200 223478 600 8 la_oen[86]
port 483 nsew default input
rlabel metal2 s 225206 -1200 225318 600 8 la_oen[87]
port 484 nsew default input
rlabel metal2 s 227046 -1200 227158 600 8 la_oen[88]
port 485 nsew default input
rlabel metal2 s 228886 -1200 228998 600 8 la_oen[89]
port 486 nsew default input
rlabel metal2 s 80674 -1200 80786 600 8 la_oen[8]
port 487 nsew default input
rlabel metal2 s 230726 -1200 230838 600 8 la_oen[90]
port 488 nsew default input
rlabel metal2 s 232566 -1200 232678 600 8 la_oen[91]
port 489 nsew default input
rlabel metal2 s 234406 -1200 234518 600 8 la_oen[92]
port 490 nsew default input
rlabel metal2 s 236246 -1200 236358 600 8 la_oen[93]
port 491 nsew default input
rlabel metal2 s 237994 -1200 238106 600 8 la_oen[94]
port 492 nsew default input
rlabel metal2 s 239834 -1200 239946 600 8 la_oen[95]
port 493 nsew default input
rlabel metal2 s 241674 -1200 241786 600 8 la_oen[96]
port 494 nsew default input
rlabel metal2 s 243514 -1200 243626 600 8 la_oen[97]
port 495 nsew default input
rlabel metal2 s 245354 -1200 245466 600 8 la_oen[98]
port 496 nsew default input
rlabel metal2 s 247194 -1200 247306 600 8 la_oen[99]
port 497 nsew default input
rlabel metal2 s 82514 -1200 82626 600 8 la_oen[9]
port 498 nsew default input
rlabel metal2 s 298622 299400 298734 301200 6 vccd1
port 499 nsew default bidirectional
rlabel metal3 s -1200 74884 600 75124 4 vccd2
port 500 nsew default bidirectional
rlabel metal3 s 299400 49860 301200 50100 6 vdda1
port 501 nsew default bidirectional
rlabel metal3 s -1200 224892 600 225132 4 vdda2
port 502 nsew default bidirectional
rlabel metal2 s 298990 -1200 299102 600 8 vssa1
port 503 nsew default bidirectional
rlabel metal2 s 299634 -1200 299746 600 8 vssa2
port 504 nsew default bidirectional
rlabel metal3 s 299400 149820 301200 150060 6 vssd1
port 505 nsew default bidirectional
rlabel metal3 s 299400 249780 301200 250020 6 vssd2
port 506 nsew default bidirectional
rlabel metal2 s 266 -1200 378 600 8 wb_clk_i
port 507 nsew default input
rlabel metal2 s 308 600 336 4082 6 wb_clk_i
port 507 nsew default input
rlabel metal2 s 296 4082 348 4146 6 wb_clk_i
port 507 nsew default input
rlabel via1 s 296 4088 348 4140 6 wb_clk_i
port 507 nsew default input
rlabel metal1 s 290 4088 354 4100 6 wb_clk_i
port 507 nsew default input
rlabel metal1 s 290 4100 1340 4128 6 wb_clk_i
port 507 nsew default input
rlabel metal1 s 290 4128 354 4140 6 wb_clk_i
port 507 nsew default input
rlabel metal2 s 818 -1200 930 600 8 wb_rst_i
port 508 nsew default input
rlabel metal2 s 860 600 888 3402 6 wb_rst_i
port 508 nsew default input
rlabel metal2 s 848 3402 900 3466 6 wb_rst_i
port 508 nsew default input
rlabel via1 s 848 3408 900 3460 6 wb_rst_i
port 508 nsew default input
rlabel metal1 s 842 3408 906 3420 6 wb_rst_i
port 508 nsew default input
rlabel metal1 s 842 3420 1340 3448 6 wb_rst_i
port 508 nsew default input
rlabel metal1 s 842 3448 906 3460 6 wb_rst_i
port 508 nsew default input
rlabel metal2 s 1462 -1200 1574 600 8 wbs_ack_o
port 509 nsew default output
rlabel metal2 s 1504 600 1532 1340 6 wbs_ack_o
port 509 nsew default output
rlabel metal2 s 3854 -1200 3966 600 8 wbs_adr_i[0]
port 510 nsew default input
rlabel metal2 s 24646 -1200 24758 600 8 wbs_adr_i[10]
port 511 nsew default input
rlabel metal2 s 26486 -1200 26598 600 8 wbs_adr_i[11]
port 512 nsew default input
rlabel metal2 s 28234 -1200 28346 600 8 wbs_adr_i[12]
port 513 nsew default input
rlabel metal2 s 30074 -1200 30186 600 8 wbs_adr_i[13]
port 514 nsew default input
rlabel metal2 s 31914 -1200 32026 600 8 wbs_adr_i[14]
port 515 nsew default input
rlabel metal2 s 33754 -1200 33866 600 8 wbs_adr_i[15]
port 516 nsew default input
rlabel metal2 s 35594 -1200 35706 600 8 wbs_adr_i[16]
port 517 nsew default input
rlabel metal2 s 37434 -1200 37546 600 8 wbs_adr_i[17]
port 518 nsew default input
rlabel metal2 s 39274 -1200 39386 600 8 wbs_adr_i[18]
port 519 nsew default input
rlabel metal2 s 41114 -1200 41226 600 8 wbs_adr_i[19]
port 520 nsew default input
rlabel metal2 s 6338 -1200 6450 600 8 wbs_adr_i[1]
port 521 nsew default input
rlabel metal2 s 42862 -1200 42974 600 8 wbs_adr_i[20]
port 522 nsew default input
rlabel metal2 s 44702 -1200 44814 600 8 wbs_adr_i[21]
port 523 nsew default input
rlabel metal2 s 46542 -1200 46654 600 8 wbs_adr_i[22]
port 524 nsew default input
rlabel metal2 s 48382 -1200 48494 600 8 wbs_adr_i[23]
port 525 nsew default input
rlabel metal2 s 50222 -1200 50334 600 8 wbs_adr_i[24]
port 526 nsew default input
rlabel metal2 s 52062 -1200 52174 600 8 wbs_adr_i[25]
port 527 nsew default input
rlabel metal2 s 53902 -1200 54014 600 8 wbs_adr_i[26]
port 528 nsew default input
rlabel metal2 s 55742 -1200 55854 600 8 wbs_adr_i[27]
port 529 nsew default input
rlabel metal2 s 57582 -1200 57694 600 8 wbs_adr_i[28]
port 530 nsew default input
rlabel metal2 s 59330 -1200 59442 600 8 wbs_adr_i[29]
port 531 nsew default input
rlabel metal2 s 8730 -1200 8842 600 8 wbs_adr_i[2]
port 532 nsew default input
rlabel metal2 s 61170 -1200 61282 600 8 wbs_adr_i[30]
port 533 nsew default input
rlabel metal2 s 63010 -1200 63122 600 8 wbs_adr_i[31]
port 534 nsew default input
rlabel metal2 s 11214 -1200 11326 600 8 wbs_adr_i[3]
port 535 nsew default input
rlabel metal2 s 13606 -1200 13718 600 8 wbs_adr_i[4]
port 536 nsew default input
rlabel metal2 s 15446 -1200 15558 600 8 wbs_adr_i[5]
port 537 nsew default input
rlabel metal2 s 17286 -1200 17398 600 8 wbs_adr_i[6]
port 538 nsew default input
rlabel metal2 s 19126 -1200 19238 600 8 wbs_adr_i[7]
port 539 nsew default input
rlabel metal2 s 20966 -1200 21078 600 8 wbs_adr_i[8]
port 540 nsew default input
rlabel metal2 s 22806 -1200 22918 600 8 wbs_adr_i[9]
port 541 nsew default input
rlabel metal2 s 2014 -1200 2126 600 8 wbs_cyc_i
port 542 nsew default input
rlabel metal2 s 2056 600 2084 1340 6 wbs_cyc_i
port 542 nsew default input
rlabel metal2 s 4498 -1200 4610 600 8 wbs_dat_i[0]
port 543 nsew default input
rlabel metal2 s 4540 600 4568 1340 6 wbs_dat_i[0]
port 543 nsew default input
rlabel metal2 s 25198 -1200 25310 600 8 wbs_dat_i[10]
port 544 nsew default input
rlabel metal2 s 25240 600 25268 1340 6 wbs_dat_i[10]
port 544 nsew default input
rlabel metal2 s 27038 -1200 27150 600 8 wbs_dat_i[11]
port 545 nsew default input
rlabel metal2 s 27080 600 27108 1340 6 wbs_dat_i[11]
port 545 nsew default input
rlabel metal2 s 28878 -1200 28990 600 8 wbs_dat_i[12]
port 546 nsew default input
rlabel metal2 s 28920 600 28948 1340 6 wbs_dat_i[12]
port 546 nsew default input
rlabel metal2 s 30718 -1200 30830 600 8 wbs_dat_i[13]
port 547 nsew default input
rlabel metal2 s 30760 600 30788 1340 6 wbs_dat_i[13]
port 547 nsew default input
rlabel metal2 s 32558 -1200 32670 600 8 wbs_dat_i[14]
port 548 nsew default input
rlabel metal2 s 32600 600 32628 1340 6 wbs_dat_i[14]
port 548 nsew default input
rlabel metal2 s 34398 -1200 34510 600 8 wbs_dat_i[15]
port 549 nsew default input
rlabel metal2 s 34440 600 34468 1340 6 wbs_dat_i[15]
port 549 nsew default input
rlabel metal2 s 36238 -1200 36350 600 8 wbs_dat_i[16]
port 550 nsew default input
rlabel metal2 s 36280 600 36308 1340 6 wbs_dat_i[16]
port 550 nsew default input
rlabel metal2 s 37986 -1200 38098 600 8 wbs_dat_i[17]
port 551 nsew default input
rlabel metal2 s 38028 600 38056 1340 6 wbs_dat_i[17]
port 551 nsew default input
rlabel metal2 s 39826 -1200 39938 600 8 wbs_dat_i[18]
port 552 nsew default input
rlabel metal2 s 39868 600 39896 1340 6 wbs_dat_i[18]
port 552 nsew default input
rlabel metal2 s 41666 -1200 41778 598 8 wbs_dat_i[19]
port 553 nsew default input
rlabel metal2 s 41666 598 41828 600 6 wbs_dat_i[19]
port 553 nsew default input
rlabel metal2 s 41708 600 41828 626 6 wbs_dat_i[19]
port 553 nsew default input
rlabel metal2 s 41800 626 41828 1340 6 wbs_dat_i[19]
port 553 nsew default input
rlabel metal2 s 6890 -1200 7002 600 8 wbs_dat_i[1]
port 554 nsew default input
rlabel metal2 s 6932 600 6960 1340 6 wbs_dat_i[1]
port 554 nsew default input
rlabel metal2 s 43506 -1200 43618 600 8 wbs_dat_i[20]
port 555 nsew default input
rlabel metal2 s 43548 600 43576 1340 6 wbs_dat_i[20]
port 555 nsew default input
rlabel metal2 s 45346 -1200 45458 600 8 wbs_dat_i[21]
port 556 nsew default input
rlabel metal2 s 45388 600 45416 1340 6 wbs_dat_i[21]
port 556 nsew default input
rlabel metal2 s 47186 -1200 47298 600 8 wbs_dat_i[22]
port 557 nsew default input
rlabel metal2 s 47228 600 47256 1340 6 wbs_dat_i[22]
port 557 nsew default input
rlabel metal2 s 49026 -1200 49138 600 8 wbs_dat_i[23]
port 558 nsew default input
rlabel metal2 s 49068 600 49096 1340 6 wbs_dat_i[23]
port 558 nsew default input
rlabel metal2 s 50866 -1200 50978 600 8 wbs_dat_i[24]
port 559 nsew default input
rlabel metal2 s 50908 600 50936 1340 6 wbs_dat_i[24]
port 559 nsew default input
rlabel metal2 s 52706 -1200 52818 600 8 wbs_dat_i[25]
port 560 nsew default input
rlabel metal2 s 52748 600 52776 1340 6 wbs_dat_i[25]
port 560 nsew default input
rlabel metal2 s 54454 -1200 54566 598 8 wbs_dat_i[26]
port 561 nsew default input
rlabel metal2 s 54312 598 54566 600 6 wbs_dat_i[26]
port 561 nsew default input
rlabel metal2 s 54312 600 54524 626 6 wbs_dat_i[26]
port 561 nsew default input
rlabel metal2 s 54312 626 54340 1340 6 wbs_dat_i[26]
port 561 nsew default input
rlabel metal2 s 56294 -1200 56406 598 8 wbs_dat_i[27]
port 562 nsew default input
rlabel metal2 s 56152 598 56406 600 6 wbs_dat_i[27]
port 562 nsew default input
rlabel metal2 s 56152 600 56364 626 6 wbs_dat_i[27]
port 562 nsew default input
rlabel metal2 s 56152 626 56180 1340 6 wbs_dat_i[27]
port 562 nsew default input
rlabel metal2 s 58134 -1200 58246 600 8 wbs_dat_i[28]
port 563 nsew default input
rlabel metal2 s 58176 600 58204 1340 6 wbs_dat_i[28]
port 563 nsew default input
rlabel metal2 s 59974 -1200 60086 598 8 wbs_dat_i[29]
port 564 nsew default input
rlabel metal2 s 59974 598 60136 600 6 wbs_dat_i[29]
port 564 nsew default input
rlabel metal2 s 60016 600 60136 626 6 wbs_dat_i[29]
port 564 nsew default input
rlabel metal2 s 60108 626 60136 1340 6 wbs_dat_i[29]
port 564 nsew default input
rlabel metal2 s 9374 -1200 9486 600 8 wbs_dat_i[2]
port 565 nsew default input
rlabel metal2 s 9416 600 9444 1340 6 wbs_dat_i[2]
port 565 nsew default input
rlabel metal2 s 61814 -1200 61926 600 8 wbs_dat_i[30]
port 566 nsew default input
rlabel metal2 s 61856 600 61884 1340 6 wbs_dat_i[30]
port 566 nsew default input
rlabel metal2 s 63654 -1200 63766 600 8 wbs_dat_i[31]
port 567 nsew default input
rlabel metal2 s 63696 600 63724 1340 6 wbs_dat_i[31]
port 567 nsew default input
rlabel metal2 s 11766 -1200 11878 600 8 wbs_dat_i[3]
port 568 nsew default input
rlabel metal2 s 11808 600 11836 1340 6 wbs_dat_i[3]
port 568 nsew default input
rlabel metal2 s 14250 -1200 14362 600 8 wbs_dat_i[4]
port 569 nsew default input
rlabel metal2 s 14292 600 14320 1340 6 wbs_dat_i[4]
port 569 nsew default input
rlabel metal2 s 16090 -1200 16202 600 8 wbs_dat_i[5]
port 570 nsew default input
rlabel metal2 s 16132 600 16160 1340 6 wbs_dat_i[5]
port 570 nsew default input
rlabel metal2 s 17930 -1200 18042 600 8 wbs_dat_i[6]
port 571 nsew default input
rlabel metal2 s 17972 600 18000 1340 6 wbs_dat_i[6]
port 571 nsew default input
rlabel metal2 s 19770 -1200 19882 600 8 wbs_dat_i[7]
port 572 nsew default input
rlabel metal2 s 19812 600 19840 1340 6 wbs_dat_i[7]
port 572 nsew default input
rlabel metal2 s 21518 -1200 21630 600 8 wbs_dat_i[8]
port 573 nsew default input
rlabel metal2 s 21560 600 21588 1340 6 wbs_dat_i[8]
port 573 nsew default input
rlabel metal2 s 23358 -1200 23470 600 8 wbs_dat_i[9]
port 574 nsew default input
rlabel metal2 s 23400 600 23428 1340 6 wbs_dat_i[9]
port 574 nsew default input
rlabel metal2 s 5142 -1200 5254 600 8 wbs_dat_o[0]
port 575 nsew default output
rlabel metal2 s 5184 600 5212 1340 6 wbs_dat_o[0]
port 575 nsew default output
rlabel metal2 s 25842 -1200 25954 600 8 wbs_dat_o[10]
port 576 nsew default output
rlabel metal2 s 25884 600 25912 1340 6 wbs_dat_o[10]
port 576 nsew default output
rlabel metal2 s 27682 -1200 27794 600 8 wbs_dat_o[11]
port 577 nsew default output
rlabel metal2 s 27724 600 27752 1340 6 wbs_dat_o[11]
port 577 nsew default output
rlabel metal2 s 29522 -1200 29634 600 8 wbs_dat_o[12]
port 578 nsew default output
rlabel metal2 s 29564 600 29592 1340 6 wbs_dat_o[12]
port 578 nsew default output
rlabel metal2 s 31362 -1200 31474 600 8 wbs_dat_o[13]
port 579 nsew default output
rlabel metal2 s 31404 600 31432 1340 6 wbs_dat_o[13]
port 579 nsew default output
rlabel metal2 s 33110 -1200 33222 600 8 wbs_dat_o[14]
port 580 nsew default output
rlabel metal2 s 33152 600 33180 1340 6 wbs_dat_o[14]
port 580 nsew default output
rlabel metal2 s 34950 -1200 35062 600 8 wbs_dat_o[15]
port 581 nsew default output
rlabel metal2 s 34992 600 35020 1340 6 wbs_dat_o[15]
port 581 nsew default output
rlabel metal2 s 36790 -1200 36902 600 8 wbs_dat_o[16]
port 582 nsew default output
rlabel metal2 s 36832 600 36860 1340 6 wbs_dat_o[16]
port 582 nsew default output
rlabel metal2 s 38630 -1200 38742 600 8 wbs_dat_o[17]
port 583 nsew default output
rlabel metal2 s 38672 600 38700 1340 6 wbs_dat_o[17]
port 583 nsew default output
rlabel metal2 s 40470 -1200 40582 600 8 wbs_dat_o[18]
port 584 nsew default output
rlabel metal2 s 40512 600 40540 1340 6 wbs_dat_o[18]
port 584 nsew default output
rlabel metal2 s 42310 -1200 42422 600 8 wbs_dat_o[19]
port 585 nsew default output
rlabel metal2 s 42352 600 42380 1340 6 wbs_dat_o[19]
port 585 nsew default output
rlabel metal2 s 7534 -1200 7646 600 8 wbs_dat_o[1]
port 586 nsew default output
rlabel metal2 s 7576 600 7604 1340 6 wbs_dat_o[1]
port 586 nsew default output
rlabel metal2 s 44150 -1200 44262 600 8 wbs_dat_o[20]
port 587 nsew default output
rlabel metal2 s 44192 600 44220 1340 6 wbs_dat_o[20]
port 587 nsew default output
rlabel metal2 s 45990 -1200 46102 600 8 wbs_dat_o[21]
port 588 nsew default output
rlabel metal2 s 46032 600 46060 1340 6 wbs_dat_o[21]
port 588 nsew default output
rlabel metal2 s 47738 -1200 47850 600 8 wbs_dat_o[22]
port 589 nsew default output
rlabel metal2 s 47780 600 47808 1340 6 wbs_dat_o[22]
port 589 nsew default output
rlabel metal2 s 49578 -1200 49690 600 8 wbs_dat_o[23]
port 590 nsew default output
rlabel metal2 s 49620 600 49648 1340 6 wbs_dat_o[23]
port 590 nsew default output
rlabel metal2 s 51418 -1200 51530 598 8 wbs_dat_o[24]
port 591 nsew default output
rlabel metal2 s 51368 598 51530 600 6 wbs_dat_o[24]
port 591 nsew default output
rlabel metal2 s 51368 600 51488 626 6 wbs_dat_o[24]
port 591 nsew default output
rlabel metal2 s 51368 626 51396 1340 6 wbs_dat_o[24]
port 591 nsew default output
rlabel metal2 s 53258 -1200 53370 600 8 wbs_dat_o[25]
port 592 nsew default output
rlabel metal2 s 53300 600 53328 1340 6 wbs_dat_o[25]
port 592 nsew default output
rlabel metal2 s 55098 -1200 55210 598 8 wbs_dat_o[26]
port 593 nsew default output
rlabel metal2 s 55098 598 55260 600 6 wbs_dat_o[26]
port 593 nsew default output
rlabel metal2 s 55140 600 55260 626 6 wbs_dat_o[26]
port 593 nsew default output
rlabel metal2 s 55232 626 55260 1340 6 wbs_dat_o[26]
port 593 nsew default output
rlabel metal2 s 56938 -1200 57050 600 8 wbs_dat_o[27]
port 594 nsew default output
rlabel metal2 s 56980 600 57008 1340 6 wbs_dat_o[27]
port 594 nsew default output
rlabel metal2 s 58778 -1200 58890 600 8 wbs_dat_o[28]
port 595 nsew default output
rlabel metal2 s 58820 600 58848 1340 6 wbs_dat_o[28]
port 595 nsew default output
rlabel metal2 s 60618 -1200 60730 600 8 wbs_dat_o[29]
port 596 nsew default output
rlabel metal2 s 60660 600 60688 1340 6 wbs_dat_o[29]
port 596 nsew default output
rlabel metal2 s 10018 -1200 10130 600 8 wbs_dat_o[2]
port 597 nsew default output
rlabel metal2 s 10060 600 10088 1340 6 wbs_dat_o[2]
port 597 nsew default output
rlabel metal2 s 62458 -1200 62570 600 8 wbs_dat_o[30]
port 598 nsew default output
rlabel metal2 s 62500 600 62528 1340 6 wbs_dat_o[30]
port 598 nsew default output
rlabel metal2 s 64206 -1200 64318 600 8 wbs_dat_o[31]
port 599 nsew default output
rlabel metal2 s 64248 600 64276 1340 6 wbs_dat_o[31]
port 599 nsew default output
rlabel metal2 s 12410 -1200 12522 600 8 wbs_dat_o[3]
port 600 nsew default output
rlabel metal2 s 12452 600 12480 1340 6 wbs_dat_o[3]
port 600 nsew default output
rlabel metal2 s 14894 -1200 15006 600 8 wbs_dat_o[4]
port 601 nsew default output
rlabel metal2 s 14936 600 14964 1340 6 wbs_dat_o[4]
port 601 nsew default output
rlabel metal2 s 16642 -1200 16754 600 8 wbs_dat_o[5]
port 602 nsew default output
rlabel metal2 s 16684 600 16712 1340 6 wbs_dat_o[5]
port 602 nsew default output
rlabel metal2 s 18482 -1200 18594 600 8 wbs_dat_o[6]
port 603 nsew default output
rlabel metal2 s 18524 600 18552 1340 6 wbs_dat_o[6]
port 603 nsew default output
rlabel metal2 s 20322 -1200 20434 600 8 wbs_dat_o[7]
port 604 nsew default output
rlabel metal2 s 20364 600 20392 1340 6 wbs_dat_o[7]
port 604 nsew default output
rlabel metal2 s 22162 -1200 22274 600 8 wbs_dat_o[8]
port 605 nsew default output
rlabel metal2 s 22204 600 22232 1340 6 wbs_dat_o[8]
port 605 nsew default output
rlabel metal2 s 24002 -1200 24114 600 8 wbs_dat_o[9]
port 606 nsew default output
rlabel metal2 s 24044 600 24072 1340 6 wbs_dat_o[9]
port 606 nsew default output
rlabel metal2 s 5694 -1200 5806 600 8 wbs_sel_i[0]
port 607 nsew default input
rlabel metal2 s 5736 600 5764 1340 6 wbs_sel_i[0]
port 607 nsew default input
rlabel metal2 s 8178 -1200 8290 600 8 wbs_sel_i[1]
port 608 nsew default input
rlabel metal2 s 8220 600 8248 1340 6 wbs_sel_i[1]
port 608 nsew default input
rlabel metal2 s 10570 -1200 10682 600 8 wbs_sel_i[2]
port 609 nsew default input
rlabel metal2 s 10612 600 10640 1340 6 wbs_sel_i[2]
port 609 nsew default input
rlabel metal2 s 13054 -1200 13166 600 8 wbs_sel_i[3]
port 610 nsew default input
rlabel metal2 s 13096 600 13124 1340 6 wbs_sel_i[3]
port 610 nsew default input
rlabel metal2 s 2658 -1200 2770 600 8 wbs_stb_i
port 611 nsew default input
rlabel metal2 s 2700 600 2728 1340 6 wbs_stb_i
port 611 nsew default input
rlabel metal2 s 3302 -1200 3414 600 8 wbs_we_i
port 612 nsew default input
rlabel metal2 s 3344 600 3372 1340 6 wbs_we_i
port 612 nsew default input
rlabel metal5 s 298660 1874 299116 2478 6 VPWR
port 613 nsew power input
rlabel metal5 s 804 1874 1340 2478 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 5986 300056 6306 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 5986 1340 6306 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 21304 300056 21624 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 21304 1340 21624 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 36622 300056 36942 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 36622 1340 36942 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 51940 300056 52260 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 51940 1340 52260 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 67258 300056 67578 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 67258 1340 67578 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 82576 300056 82896 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 82576 1340 82896 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 97894 300056 98214 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 97894 1340 98214 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 113212 300056 113532 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 113212 1340 113532 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 128530 300056 128850 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 128530 1340 128850 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 143848 300056 144168 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 143848 1340 144168 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 159166 300056 159486 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 159166 1340 159486 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 174484 300056 174804 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 174484 1340 174804 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 189802 300056 190122 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 189802 1340 190122 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 205120 300056 205440 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 205120 1340 205440 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 220438 300056 220758 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 220438 1340 220758 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 235756 300056 236076 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 235756 1340 236076 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 251074 300056 251394 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 251074 1340 251394 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 266392 300056 266712 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 266392 1340 266712 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 281710 300056 282030 6 VPWR
port 613 nsew power input
rlabel metal5 s -136 281710 1340 282030 6 VPWR
port 613 nsew power input
rlabel metal5 s 298660 297266 299116 297870 6 VPWR
port 613 nsew power input
rlabel metal5 s 804 297266 1340 297870 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 1898 298934 2134 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 2218 298934 2454 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 6028 298934 6264 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 21346 298934 21582 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 36664 298934 36900 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 51982 298934 52218 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 67300 298934 67536 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 82618 298934 82854 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 97936 298934 98172 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 113254 298934 113490 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 128572 298934 128808 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 143890 298934 144126 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 159208 298934 159444 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 174526 298934 174762 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 189844 298934 190080 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 205162 298934 205398 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 220480 298934 220716 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 235798 298934 236034 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 251116 298934 251352 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 266434 298934 266670 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 281752 298934 281988 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 297290 298934 297526 6 VPWR
port 613 nsew power input
rlabel via4 s 298698 297610 298934 297846 6 VPWR
port 613 nsew power input
rlabel via4 s 986 1898 1222 2134 6 VPWR
port 613 nsew power input
rlabel via4 s 986 2218 1222 2454 6 VPWR
port 613 nsew power input
rlabel via4 s 986 6028 1222 6264 6 VPWR
port 613 nsew power input
rlabel via4 s 986 21346 1222 21582 6 VPWR
port 613 nsew power input
rlabel via4 s 986 36664 1222 36900 6 VPWR
port 613 nsew power input
rlabel via4 s 986 51982 1222 52218 6 VPWR
port 613 nsew power input
rlabel via4 s 986 67300 1222 67536 6 VPWR
port 613 nsew power input
rlabel via4 s 986 82618 1222 82854 6 VPWR
port 613 nsew power input
rlabel via4 s 986 97936 1222 98172 6 VPWR
port 613 nsew power input
rlabel via4 s 986 113254 1222 113490 6 VPWR
port 613 nsew power input
rlabel via4 s 986 128572 1222 128808 6 VPWR
port 613 nsew power input
rlabel via4 s 986 143890 1222 144126 6 VPWR
port 613 nsew power input
rlabel via4 s 986 159208 1222 159444 6 VPWR
port 613 nsew power input
rlabel via4 s 986 174526 1222 174762 6 VPWR
port 613 nsew power input
rlabel via4 s 986 189844 1222 190080 6 VPWR
port 613 nsew power input
rlabel via4 s 986 205162 1222 205398 6 VPWR
port 613 nsew power input
rlabel via4 s 986 220480 1222 220716 6 VPWR
port 613 nsew power input
rlabel via4 s 986 235798 1222 236034 6 VPWR
port 613 nsew power input
rlabel via4 s 986 251116 1222 251352 6 VPWR
port 613 nsew power input
rlabel via4 s 986 266434 1222 266670 6 VPWR
port 613 nsew power input
rlabel via4 s 986 281752 1222 281988 6 VPWR
port 613 nsew power input
rlabel via4 s 986 297290 1222 297526 6 VPWR
port 613 nsew power input
rlabel via4 s 986 297610 1222 297846 6 VPWR
port 613 nsew power input
rlabel metal4 s 281328 936 281648 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 250608 936 250928 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 219888 936 220208 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 189168 936 189488 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 158448 936 158768 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 127728 936 128048 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 97008 936 97328 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 66288 936 66608 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 35568 936 35888 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 4848 936 5168 1340 6 VPWR
port 613 nsew power input
rlabel metal4 s 298660 1876 299116 297868 6 VPWR
port 613 nsew power input
rlabel metal4 s 804 1876 1340 297868 6 VPWR
port 613 nsew power input
rlabel metal4 s 281328 298660 281648 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 250608 298660 250928 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 219888 298660 220208 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 189168 298660 189488 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 158448 298660 158768 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 127728 298660 128048 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 97008 298660 97328 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 66288 298660 66608 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 35568 298660 35888 298808 6 VPWR
port 613 nsew power input
rlabel metal4 s 4848 298660 5168 298808 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 2128 298816 2224 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 2128 1340 2224 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 3216 298816 3312 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 3216 1340 3312 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 4304 298816 4400 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 4304 1340 4400 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 5392 298816 5488 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 5392 1340 5488 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 6480 298816 6576 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 6480 1340 6576 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 7568 298816 7664 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 7568 1340 7664 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 8656 298816 8752 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 8656 1340 8752 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 9744 298816 9840 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 9744 1340 9840 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 10832 298816 10928 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 10832 1340 10928 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 11920 298816 12016 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 11920 1340 12016 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 13008 298816 13104 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 13008 1340 13104 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 14096 298816 14192 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 14096 1340 14192 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 15184 298816 15280 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 15184 1340 15280 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 16272 298816 16368 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 16272 1340 16368 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 17360 298816 17456 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 17360 1340 17456 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 18448 298816 18544 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 18448 1340 18544 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 19536 298816 19632 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 19536 1340 19632 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 20624 298816 20720 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 20624 1340 20720 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 21712 298816 21808 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 21712 1340 21808 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 22800 298816 22896 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 22800 1340 22896 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 23888 298816 23984 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 23888 1340 23984 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 24976 298816 25072 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 24976 1340 25072 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 26064 298816 26160 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 26064 1340 26160 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 27152 298816 27248 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 27152 1340 27248 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 28240 298816 28336 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 28240 1340 28336 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 29328 298816 29424 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 29328 1340 29424 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 30416 298816 30512 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 30416 1340 30512 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 31504 298816 31600 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 31504 1340 31600 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 32592 298816 32688 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 32592 1340 32688 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 33680 298816 33776 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 33680 1340 33776 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 34768 298816 34864 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 34768 1340 34864 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 35856 298816 35952 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 35856 1340 35952 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 36944 298816 37040 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 36944 1340 37040 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 38032 298816 38128 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 38032 1340 38128 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 39120 298816 39216 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 39120 1340 39216 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 40208 298816 40304 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 40208 1340 40304 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 41296 298816 41392 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 41296 1340 41392 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 42384 298816 42480 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 42384 1340 42480 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 43472 298816 43568 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 43472 1340 43568 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 44560 298816 44656 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 44560 1340 44656 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 45648 298816 45744 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 45648 1340 45744 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 46736 298816 46832 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 46736 1340 46832 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 47824 298816 47920 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 47824 1340 47920 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 48912 298816 49008 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 48912 1340 49008 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 50000 298816 50096 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 50000 1340 50096 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 51088 298816 51184 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 51088 1340 51184 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 52176 298816 52272 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 52176 1340 52272 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 53264 298816 53360 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 53264 1340 53360 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 54352 298816 54448 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 54352 1340 54448 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 55440 298816 55536 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 55440 1340 55536 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 56528 298816 56624 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 56528 1340 56624 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 57616 298816 57712 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 57616 1340 57712 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 58704 298816 58800 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 58704 1340 58800 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 59792 298816 59888 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 59792 1340 59888 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 60880 298816 60976 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 60880 1340 60976 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 61968 298816 62064 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 61968 1340 62064 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 63056 298816 63152 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 63056 1340 63152 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 64144 298816 64240 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 64144 1340 64240 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 65232 298816 65328 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 65232 1340 65328 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 66320 298816 66416 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 66320 1340 66416 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 67408 298816 67504 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 67408 1340 67504 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 68496 298816 68592 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 68496 1340 68592 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 69584 298816 69680 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 69584 1340 69680 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 70672 298816 70768 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 70672 1340 70768 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 71760 298816 71856 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 71760 1340 71856 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 72848 298816 72944 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 72848 1340 72944 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 73936 298816 74032 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 73936 1340 74032 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 75024 298816 75120 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 75024 1340 75120 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 76112 298816 76208 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 76112 1340 76208 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 77200 298816 77296 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 77200 1340 77296 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 78288 298816 78384 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 78288 1340 78384 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 79376 298816 79472 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 79376 1340 79472 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 80464 298816 80560 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 80464 1340 80560 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 81552 298816 81648 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 81552 1340 81648 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 82640 298816 82736 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 82640 1340 82736 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 83728 298816 83824 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 83728 1340 83824 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 84816 298816 84912 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 84816 1340 84912 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 85904 298816 86000 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 85904 1340 86000 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 86992 298816 87088 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 86992 1340 87088 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 88080 298816 88176 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 88080 1340 88176 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 89168 298816 89264 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 89168 1340 89264 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 90256 298816 90352 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 90256 1340 90352 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 91344 298816 91440 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 91344 1340 91440 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 92432 298816 92528 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 92432 1340 92528 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 93520 298816 93616 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 93520 1340 93616 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 94608 298816 94704 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 94608 1340 94704 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 95696 298816 95792 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 95696 1340 95792 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 96784 298816 96880 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 96784 1340 96880 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 97872 298816 97968 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 97872 1340 97968 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 98960 298816 99056 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 98960 1340 99056 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 100048 298816 100144 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 100048 1340 100144 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 101136 298816 101232 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 101136 1340 101232 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 102224 298816 102320 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 102224 1340 102320 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 103312 298816 103408 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 103312 1340 103408 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 104400 298816 104496 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 104400 1340 104496 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 105488 298816 105584 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 105488 1340 105584 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 106576 298816 106672 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 106576 1340 106672 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 107664 298816 107760 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 107664 1340 107760 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 108752 298816 108848 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 108752 1340 108848 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 109840 298816 109936 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 109840 1340 109936 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 110928 298816 111024 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 110928 1340 111024 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 112016 298816 112112 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 112016 1340 112112 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 113104 298816 113200 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 113104 1340 113200 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 114192 298816 114288 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 114192 1340 114288 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 115280 298816 115376 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 115280 1340 115376 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 116368 298816 116464 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 116368 1340 116464 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 117456 298816 117552 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 117456 1340 117552 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 118544 298816 118640 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 118544 1340 118640 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 119632 298816 119728 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 119632 1340 119728 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 120720 298816 120816 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 120720 1340 120816 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 121808 298816 121904 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 121808 1340 121904 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 122896 298816 122992 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 122896 1340 122992 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 123984 298816 124080 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 123984 1340 124080 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 125072 298816 125168 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 125072 1340 125168 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 126160 298816 126256 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 126160 1340 126256 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 127248 298816 127344 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 127248 1340 127344 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 128336 298816 128432 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 128336 1340 128432 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 129424 298816 129520 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 129424 1340 129520 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 130512 298816 130608 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 130512 1340 130608 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 131600 298816 131696 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 131600 1340 131696 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 132688 298816 132784 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 132688 1340 132784 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 133776 298816 133872 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 133776 1340 133872 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 134864 298816 134960 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 134864 1340 134960 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 135952 298816 136048 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 135952 1340 136048 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 137040 298816 137136 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 137040 1340 137136 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 138128 298816 138224 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 138128 1340 138224 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 139216 298816 139312 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 139216 1340 139312 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 140304 298816 140400 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 140304 1340 140400 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 141392 298816 141488 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 141392 1340 141488 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 142480 298816 142576 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 142480 1340 142576 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 143568 298816 143664 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 143568 1340 143664 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 144656 298816 144752 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 144656 1340 144752 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 145744 298816 145840 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 145744 1340 145840 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 146832 298816 146928 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 146832 1340 146928 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 147920 298816 148016 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 147920 1340 148016 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 149008 298816 149104 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 149008 1340 149104 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 150096 298816 150192 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 150096 1340 150192 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 151184 298816 151280 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 151184 1340 151280 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 152272 298816 152368 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 152272 1340 152368 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 153360 298816 153456 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 153360 1340 153456 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 154448 298816 154544 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 154448 1340 154544 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 155536 298816 155632 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 155536 1340 155632 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 156624 298816 156720 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 156624 1340 156720 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 157712 298816 157808 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 157712 1340 157808 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 158800 298816 158896 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 158800 1340 158896 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 159888 298816 159984 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 159888 1340 159984 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 160976 298816 161072 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 160976 1340 161072 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 162064 298816 162160 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 162064 1340 162160 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 163152 298816 163248 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 163152 1340 163248 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 164240 298816 164336 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 164240 1340 164336 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 165328 298816 165424 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 165328 1340 165424 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 166416 298816 166512 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 166416 1340 166512 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 167504 298816 167600 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 167504 1340 167600 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 168592 298816 168688 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 168592 1340 168688 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 169680 298816 169776 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 169680 1340 169776 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 170768 298816 170864 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 170768 1340 170864 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 171856 298816 171952 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 171856 1340 171952 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 172944 298816 173040 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 172944 1340 173040 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 174032 298816 174128 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 174032 1340 174128 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 175120 298816 175216 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 175120 1340 175216 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 176208 298816 176304 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 176208 1340 176304 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 177296 298816 177392 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 177296 1340 177392 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 178384 298816 178480 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 178384 1340 178480 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 179472 298816 179568 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 179472 1340 179568 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 180560 298816 180656 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 180560 1340 180656 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 181648 298816 181744 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 181648 1340 181744 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 182736 298816 182832 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 182736 1340 182832 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 183824 298816 183920 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 183824 1340 183920 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 184912 298816 185008 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 184912 1340 185008 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 186000 298816 186096 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 186000 1340 186096 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 187088 298816 187184 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 187088 1340 187184 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 188176 298816 188272 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 188176 1340 188272 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 189264 298816 189360 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 189264 1340 189360 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 190352 298816 190448 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 190352 1340 190448 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 191440 298816 191536 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 191440 1340 191536 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 192528 298816 192624 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 192528 1340 192624 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 193616 298816 193712 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 193616 1340 193712 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 194704 298816 194800 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 194704 1340 194800 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 195792 298816 195888 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 195792 1340 195888 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 196880 298816 196976 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 196880 1340 196976 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 197968 298816 198064 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 197968 1340 198064 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 199056 298816 199152 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 199056 1340 199152 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 200144 298816 200240 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 200144 1340 200240 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 201232 298816 201328 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 201232 1340 201328 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 202320 298816 202416 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 202320 1340 202416 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 203408 298816 203504 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 203408 1340 203504 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 204496 298816 204592 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 204496 1340 204592 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 205584 298816 205680 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 205584 1340 205680 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 206672 298816 206768 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 206672 1340 206768 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 207760 298816 207856 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 207760 1340 207856 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 208848 298816 208944 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 208848 1340 208944 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 209936 298816 210032 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 209936 1340 210032 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 211024 298816 211120 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 211024 1340 211120 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 212112 298816 212208 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 212112 1340 212208 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 213200 298816 213296 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 213200 1340 213296 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 214288 298816 214384 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 214288 1340 214384 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 215376 298816 215472 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 215376 1340 215472 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 216464 298816 216560 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 216464 1340 216560 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 217552 298816 217648 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 217552 1340 217648 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 218640 298816 218736 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 218640 1340 218736 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 219728 298816 219824 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 219728 1340 219824 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 220816 298816 220912 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 220816 1340 220912 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 221904 298816 222000 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 221904 1340 222000 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 222992 298816 223088 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 222992 1340 223088 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 224080 298816 224176 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 224080 1340 224176 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 225168 298816 225264 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 225168 1340 225264 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 226256 298816 226352 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 226256 1340 226352 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 227344 298816 227440 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 227344 1340 227440 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 228432 298816 228528 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 228432 1340 228528 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 229520 298816 229616 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 229520 1340 229616 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 230608 298816 230704 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 230608 1340 230704 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 231696 298816 231792 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 231696 1340 231792 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 232784 298816 232880 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 232784 1340 232880 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 233872 298816 233968 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 233872 1340 233968 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 234960 298816 235056 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 234960 1340 235056 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 236048 298816 236144 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 236048 1340 236144 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 237136 298816 237232 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 237136 1340 237232 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 238224 298816 238320 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 238224 1340 238320 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 239312 298816 239408 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 239312 1340 239408 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 240400 298816 240496 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 240400 1340 240496 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 241488 298816 241584 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 241488 1340 241584 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 242576 298816 242672 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 242576 1340 242672 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 243664 298816 243760 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 243664 1340 243760 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 244752 298816 244848 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 244752 1340 244848 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 245840 298816 245936 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 245840 1340 245936 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 246928 298816 247024 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 246928 1340 247024 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 248016 298816 248112 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 248016 1340 248112 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 249104 298816 249200 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 249104 1340 249200 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 250192 298816 250288 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 250192 1340 250288 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 251280 298816 251376 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 251280 1340 251376 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 252368 298816 252464 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 252368 1340 252464 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 253456 298816 253552 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 253456 1340 253552 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 254544 298816 254640 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 254544 1340 254640 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 255632 298816 255728 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 255632 1340 255728 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 256720 298816 256816 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 256720 1340 256816 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 257808 298816 257904 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 257808 1340 257904 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 258896 298816 258992 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 258896 1340 258992 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 259984 298816 260080 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 259984 1340 260080 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 261072 298816 261168 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 261072 1340 261168 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 262160 298816 262256 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 262160 1340 262256 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 263248 298816 263344 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 263248 1340 263344 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 264336 298816 264432 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 264336 1340 264432 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 265424 298816 265520 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 265424 1340 265520 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 266512 298816 266608 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 266512 1340 266608 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 267600 298816 267696 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 267600 1340 267696 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 268688 298816 268784 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 268688 1340 268784 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 269776 298816 269872 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 269776 1340 269872 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 270864 298816 270960 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 270864 1340 270960 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 271952 298816 272048 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 271952 1340 272048 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 273040 298816 273136 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 273040 1340 273136 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 274128 298816 274224 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 274128 1340 274224 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 275216 298816 275312 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 275216 1340 275312 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 276304 298816 276400 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 276304 1340 276400 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 277392 298816 277488 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 277392 1340 277488 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 278480 298816 278576 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 278480 1340 278576 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 279568 298816 279664 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 279568 1340 279664 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 280656 298816 280752 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 280656 1340 280752 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 281744 298816 281840 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 281744 1340 281840 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 282832 298816 282928 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 282832 1340 282928 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 283920 298816 284016 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 283920 1340 284016 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 285008 298816 285104 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 285008 1340 285104 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 286096 298816 286192 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 286096 1340 286192 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 287184 298816 287280 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 287184 1340 287280 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 288272 298816 288368 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 288272 1340 288368 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 289360 298816 289456 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 289360 1340 289456 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 290448 298816 290544 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 290448 1340 290544 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 291536 298816 291632 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 291536 1340 291632 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 292624 298816 292720 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 292624 1340 292720 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 293712 298816 293808 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 293712 1340 293808 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 294800 298816 294896 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 294800 1340 294896 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 295888 298816 295984 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 295888 1340 295984 6 VPWR
port 613 nsew power input
rlabel metal1 s 298660 296976 298816 297072 6 VPWR
port 613 nsew power input
rlabel metal1 s 1104 296976 1340 297072 6 VPWR
port 613 nsew power input
rlabel viali s 298753 2159 298787 2193 6 VPWR
port 613 nsew power input
rlabel viali s 298661 2159 298695 2193 6 VPWR
port 613 nsew power input
rlabel viali s 1317 2159 1340 2193 6 VPWR
port 613 nsew power input
rlabel viali s 1225 2159 1259 2193 6 VPWR
port 613 nsew power input
rlabel viali s 1133 2159 1167 2193 6 VPWR
port 613 nsew power input
rlabel viali s 298753 3247 298787 3281 6 VPWR
port 613 nsew power input
rlabel viali s 298661 3247 298695 3281 6 VPWR
port 613 nsew power input
rlabel viali s 1317 3247 1340 3281 6 VPWR
port 613 nsew power input
rlabel viali s 1225 3247 1259 3281 6 VPWR
port 613 nsew power input
rlabel viali s 1133 3247 1167 3281 6 VPWR
port 613 nsew power input
rlabel viali s 298753 4335 298787 4369 6 VPWR
port 613 nsew power input
rlabel viali s 298661 4335 298695 4369 6 VPWR
port 613 nsew power input
rlabel viali s 1317 4335 1340 4369 6 VPWR
port 613 nsew power input
rlabel viali s 1225 4335 1259 4369 6 VPWR
port 613 nsew power input
rlabel viali s 1133 4335 1167 4369 6 VPWR
port 613 nsew power input
rlabel viali s 298753 5423 298787 5457 6 VPWR
port 613 nsew power input
rlabel viali s 298661 5423 298695 5457 6 VPWR
port 613 nsew power input
rlabel viali s 1317 5423 1340 5457 6 VPWR
port 613 nsew power input
rlabel viali s 1225 5423 1259 5457 6 VPWR
port 613 nsew power input
rlabel viali s 1133 5423 1167 5457 6 VPWR
port 613 nsew power input
rlabel viali s 298753 6511 298787 6545 6 VPWR
port 613 nsew power input
rlabel viali s 298661 6511 298695 6545 6 VPWR
port 613 nsew power input
rlabel viali s 1317 6511 1340 6545 6 VPWR
port 613 nsew power input
rlabel viali s 1225 6511 1259 6545 6 VPWR
port 613 nsew power input
rlabel viali s 1133 6511 1167 6545 6 VPWR
port 613 nsew power input
rlabel viali s 298753 7599 298787 7633 6 VPWR
port 613 nsew power input
rlabel viali s 298661 7599 298695 7633 6 VPWR
port 613 nsew power input
rlabel viali s 1317 7599 1340 7633 6 VPWR
port 613 nsew power input
rlabel viali s 1225 7599 1259 7633 6 VPWR
port 613 nsew power input
rlabel viali s 1133 7599 1167 7633 6 VPWR
port 613 nsew power input
rlabel viali s 298753 8687 298787 8721 6 VPWR
port 613 nsew power input
rlabel viali s 298661 8687 298695 8721 6 VPWR
port 613 nsew power input
rlabel viali s 1317 8687 1340 8721 6 VPWR
port 613 nsew power input
rlabel viali s 1225 8687 1259 8721 6 VPWR
port 613 nsew power input
rlabel viali s 1133 8687 1167 8721 6 VPWR
port 613 nsew power input
rlabel viali s 298753 9775 298787 9809 6 VPWR
port 613 nsew power input
rlabel viali s 298661 9775 298695 9809 6 VPWR
port 613 nsew power input
rlabel viali s 1317 9775 1340 9809 6 VPWR
port 613 nsew power input
rlabel viali s 1225 9775 1259 9809 6 VPWR
port 613 nsew power input
rlabel viali s 1133 9775 1167 9809 6 VPWR
port 613 nsew power input
rlabel viali s 298753 10863 298787 10897 6 VPWR
port 613 nsew power input
rlabel viali s 298661 10863 298695 10897 6 VPWR
port 613 nsew power input
rlabel viali s 1317 10863 1340 10897 6 VPWR
port 613 nsew power input
rlabel viali s 1225 10863 1259 10897 6 VPWR
port 613 nsew power input
rlabel viali s 1133 10863 1167 10897 6 VPWR
port 613 nsew power input
rlabel viali s 298753 11951 298787 11985 6 VPWR
port 613 nsew power input
rlabel viali s 298661 11951 298695 11985 6 VPWR
port 613 nsew power input
rlabel viali s 1317 11951 1340 11985 6 VPWR
port 613 nsew power input
rlabel viali s 1225 11951 1259 11985 6 VPWR
port 613 nsew power input
rlabel viali s 1133 11951 1167 11985 6 VPWR
port 613 nsew power input
rlabel viali s 298753 13039 298787 13073 6 VPWR
port 613 nsew power input
rlabel viali s 298661 13039 298695 13073 6 VPWR
port 613 nsew power input
rlabel viali s 1317 13039 1340 13073 6 VPWR
port 613 nsew power input
rlabel viali s 1225 13039 1259 13073 6 VPWR
port 613 nsew power input
rlabel viali s 1133 13039 1167 13073 6 VPWR
port 613 nsew power input
rlabel viali s 298753 14127 298787 14161 6 VPWR
port 613 nsew power input
rlabel viali s 298661 14127 298695 14161 6 VPWR
port 613 nsew power input
rlabel viali s 1317 14127 1340 14161 6 VPWR
port 613 nsew power input
rlabel viali s 1225 14127 1259 14161 6 VPWR
port 613 nsew power input
rlabel viali s 1133 14127 1167 14161 6 VPWR
port 613 nsew power input
rlabel viali s 298753 15215 298787 15249 6 VPWR
port 613 nsew power input
rlabel viali s 298661 15215 298695 15249 6 VPWR
port 613 nsew power input
rlabel viali s 1317 15215 1340 15249 6 VPWR
port 613 nsew power input
rlabel viali s 1225 15215 1259 15249 6 VPWR
port 613 nsew power input
rlabel viali s 1133 15215 1167 15249 6 VPWR
port 613 nsew power input
rlabel viali s 298753 16303 298787 16337 6 VPWR
port 613 nsew power input
rlabel viali s 298661 16303 298695 16337 6 VPWR
port 613 nsew power input
rlabel viali s 1317 16303 1340 16337 6 VPWR
port 613 nsew power input
rlabel viali s 1225 16303 1259 16337 6 VPWR
port 613 nsew power input
rlabel viali s 1133 16303 1167 16337 6 VPWR
port 613 nsew power input
rlabel viali s 298753 17391 298787 17425 6 VPWR
port 613 nsew power input
rlabel viali s 298661 17391 298695 17425 6 VPWR
port 613 nsew power input
rlabel viali s 1317 17391 1340 17425 6 VPWR
port 613 nsew power input
rlabel viali s 1225 17391 1259 17425 6 VPWR
port 613 nsew power input
rlabel viali s 1133 17391 1167 17425 6 VPWR
port 613 nsew power input
rlabel viali s 298753 18479 298787 18513 6 VPWR
port 613 nsew power input
rlabel viali s 298661 18479 298695 18513 6 VPWR
port 613 nsew power input
rlabel viali s 1317 18479 1340 18513 6 VPWR
port 613 nsew power input
rlabel viali s 1225 18479 1259 18513 6 VPWR
port 613 nsew power input
rlabel viali s 1133 18479 1167 18513 6 VPWR
port 613 nsew power input
rlabel viali s 298753 19567 298787 19601 6 VPWR
port 613 nsew power input
rlabel viali s 298661 19567 298695 19601 6 VPWR
port 613 nsew power input
rlabel viali s 1317 19567 1340 19601 6 VPWR
port 613 nsew power input
rlabel viali s 1225 19567 1259 19601 6 VPWR
port 613 nsew power input
rlabel viali s 1133 19567 1167 19601 6 VPWR
port 613 nsew power input
rlabel viali s 298753 20655 298787 20689 6 VPWR
port 613 nsew power input
rlabel viali s 298661 20655 298695 20689 6 VPWR
port 613 nsew power input
rlabel viali s 1317 20655 1340 20689 6 VPWR
port 613 nsew power input
rlabel viali s 1225 20655 1259 20689 6 VPWR
port 613 nsew power input
rlabel viali s 1133 20655 1167 20689 6 VPWR
port 613 nsew power input
rlabel viali s 298753 21743 298787 21777 6 VPWR
port 613 nsew power input
rlabel viali s 298661 21743 298695 21777 6 VPWR
port 613 nsew power input
rlabel viali s 1317 21743 1340 21777 6 VPWR
port 613 nsew power input
rlabel viali s 1225 21743 1259 21777 6 VPWR
port 613 nsew power input
rlabel viali s 1133 21743 1167 21777 6 VPWR
port 613 nsew power input
rlabel viali s 298753 22831 298787 22865 6 VPWR
port 613 nsew power input
rlabel viali s 298661 22831 298695 22865 6 VPWR
port 613 nsew power input
rlabel viali s 1317 22831 1340 22865 6 VPWR
port 613 nsew power input
rlabel viali s 1225 22831 1259 22865 6 VPWR
port 613 nsew power input
rlabel viali s 1133 22831 1167 22865 6 VPWR
port 613 nsew power input
rlabel viali s 298753 23919 298787 23953 6 VPWR
port 613 nsew power input
rlabel viali s 298661 23919 298695 23953 6 VPWR
port 613 nsew power input
rlabel viali s 1317 23919 1340 23953 6 VPWR
port 613 nsew power input
rlabel viali s 1225 23919 1259 23953 6 VPWR
port 613 nsew power input
rlabel viali s 1133 23919 1167 23953 6 VPWR
port 613 nsew power input
rlabel viali s 298753 25007 298787 25041 6 VPWR
port 613 nsew power input
rlabel viali s 298661 25007 298695 25041 6 VPWR
port 613 nsew power input
rlabel viali s 1317 25007 1340 25041 6 VPWR
port 613 nsew power input
rlabel viali s 1225 25007 1259 25041 6 VPWR
port 613 nsew power input
rlabel viali s 1133 25007 1167 25041 6 VPWR
port 613 nsew power input
rlabel viali s 298753 26095 298787 26129 6 VPWR
port 613 nsew power input
rlabel viali s 298661 26095 298695 26129 6 VPWR
port 613 nsew power input
rlabel viali s 1317 26095 1340 26129 6 VPWR
port 613 nsew power input
rlabel viali s 1225 26095 1259 26129 6 VPWR
port 613 nsew power input
rlabel viali s 1133 26095 1167 26129 6 VPWR
port 613 nsew power input
rlabel viali s 298753 27183 298787 27217 6 VPWR
port 613 nsew power input
rlabel viali s 298661 27183 298695 27217 6 VPWR
port 613 nsew power input
rlabel viali s 1317 27183 1340 27217 6 VPWR
port 613 nsew power input
rlabel viali s 1225 27183 1259 27217 6 VPWR
port 613 nsew power input
rlabel viali s 1133 27183 1167 27217 6 VPWR
port 613 nsew power input
rlabel viali s 298753 28271 298787 28305 6 VPWR
port 613 nsew power input
rlabel viali s 298661 28271 298695 28305 6 VPWR
port 613 nsew power input
rlabel viali s 1317 28271 1340 28305 6 VPWR
port 613 nsew power input
rlabel viali s 1225 28271 1259 28305 6 VPWR
port 613 nsew power input
rlabel viali s 1133 28271 1167 28305 6 VPWR
port 613 nsew power input
rlabel viali s 298753 29359 298787 29393 6 VPWR
port 613 nsew power input
rlabel viali s 298661 29359 298695 29393 6 VPWR
port 613 nsew power input
rlabel viali s 1317 29359 1340 29393 6 VPWR
port 613 nsew power input
rlabel viali s 1225 29359 1259 29393 6 VPWR
port 613 nsew power input
rlabel viali s 1133 29359 1167 29393 6 VPWR
port 613 nsew power input
rlabel viali s 298753 30447 298787 30481 6 VPWR
port 613 nsew power input
rlabel viali s 298661 30447 298695 30481 6 VPWR
port 613 nsew power input
rlabel viali s 1317 30447 1340 30481 6 VPWR
port 613 nsew power input
rlabel viali s 1225 30447 1259 30481 6 VPWR
port 613 nsew power input
rlabel viali s 1133 30447 1167 30481 6 VPWR
port 613 nsew power input
rlabel viali s 298753 31535 298787 31569 6 VPWR
port 613 nsew power input
rlabel viali s 298661 31535 298695 31569 6 VPWR
port 613 nsew power input
rlabel viali s 1317 31535 1340 31569 6 VPWR
port 613 nsew power input
rlabel viali s 1225 31535 1259 31569 6 VPWR
port 613 nsew power input
rlabel viali s 1133 31535 1167 31569 6 VPWR
port 613 nsew power input
rlabel viali s 298753 32623 298787 32657 6 VPWR
port 613 nsew power input
rlabel viali s 298661 32623 298695 32657 6 VPWR
port 613 nsew power input
rlabel viali s 1317 32623 1340 32657 6 VPWR
port 613 nsew power input
rlabel viali s 1225 32623 1259 32657 6 VPWR
port 613 nsew power input
rlabel viali s 1133 32623 1167 32657 6 VPWR
port 613 nsew power input
rlabel viali s 298753 33711 298787 33745 6 VPWR
port 613 nsew power input
rlabel viali s 298661 33711 298695 33745 6 VPWR
port 613 nsew power input
rlabel viali s 1317 33711 1340 33745 6 VPWR
port 613 nsew power input
rlabel viali s 1225 33711 1259 33745 6 VPWR
port 613 nsew power input
rlabel viali s 1133 33711 1167 33745 6 VPWR
port 613 nsew power input
rlabel viali s 298753 34799 298787 34833 6 VPWR
port 613 nsew power input
rlabel viali s 298661 34799 298695 34833 6 VPWR
port 613 nsew power input
rlabel viali s 1317 34799 1340 34833 6 VPWR
port 613 nsew power input
rlabel viali s 1225 34799 1259 34833 6 VPWR
port 613 nsew power input
rlabel viali s 1133 34799 1167 34833 6 VPWR
port 613 nsew power input
rlabel viali s 298753 35887 298787 35921 6 VPWR
port 613 nsew power input
rlabel viali s 298661 35887 298695 35921 6 VPWR
port 613 nsew power input
rlabel viali s 1317 35887 1340 35921 6 VPWR
port 613 nsew power input
rlabel viali s 1225 35887 1259 35921 6 VPWR
port 613 nsew power input
rlabel viali s 1133 35887 1167 35921 6 VPWR
port 613 nsew power input
rlabel viali s 298753 36975 298787 37009 6 VPWR
port 613 nsew power input
rlabel viali s 298661 36975 298695 37009 6 VPWR
port 613 nsew power input
rlabel viali s 1317 36975 1340 37009 6 VPWR
port 613 nsew power input
rlabel viali s 1225 36975 1259 37009 6 VPWR
port 613 nsew power input
rlabel viali s 1133 36975 1167 37009 6 VPWR
port 613 nsew power input
rlabel viali s 298753 38063 298787 38097 6 VPWR
port 613 nsew power input
rlabel viali s 298661 38063 298695 38097 6 VPWR
port 613 nsew power input
rlabel viali s 1317 38063 1340 38097 6 VPWR
port 613 nsew power input
rlabel viali s 1225 38063 1259 38097 6 VPWR
port 613 nsew power input
rlabel viali s 1133 38063 1167 38097 6 VPWR
port 613 nsew power input
rlabel viali s 298753 39151 298787 39185 6 VPWR
port 613 nsew power input
rlabel viali s 298661 39151 298695 39185 6 VPWR
port 613 nsew power input
rlabel viali s 1317 39151 1340 39185 6 VPWR
port 613 nsew power input
rlabel viali s 1225 39151 1259 39185 6 VPWR
port 613 nsew power input
rlabel viali s 1133 39151 1167 39185 6 VPWR
port 613 nsew power input
rlabel viali s 298753 40239 298787 40273 6 VPWR
port 613 nsew power input
rlabel viali s 298661 40239 298695 40273 6 VPWR
port 613 nsew power input
rlabel viali s 1317 40239 1340 40273 6 VPWR
port 613 nsew power input
rlabel viali s 1225 40239 1259 40273 6 VPWR
port 613 nsew power input
rlabel viali s 1133 40239 1167 40273 6 VPWR
port 613 nsew power input
rlabel viali s 298753 41327 298787 41361 6 VPWR
port 613 nsew power input
rlabel viali s 298661 41327 298695 41361 6 VPWR
port 613 nsew power input
rlabel viali s 1317 41327 1340 41361 6 VPWR
port 613 nsew power input
rlabel viali s 1225 41327 1259 41361 6 VPWR
port 613 nsew power input
rlabel viali s 1133 41327 1167 41361 6 VPWR
port 613 nsew power input
rlabel viali s 298753 42415 298787 42449 6 VPWR
port 613 nsew power input
rlabel viali s 298661 42415 298695 42449 6 VPWR
port 613 nsew power input
rlabel viali s 1317 42415 1340 42449 6 VPWR
port 613 nsew power input
rlabel viali s 1225 42415 1259 42449 6 VPWR
port 613 nsew power input
rlabel viali s 1133 42415 1167 42449 6 VPWR
port 613 nsew power input
rlabel viali s 298753 43503 298787 43537 6 VPWR
port 613 nsew power input
rlabel viali s 298661 43503 298695 43537 6 VPWR
port 613 nsew power input
rlabel viali s 1317 43503 1340 43537 6 VPWR
port 613 nsew power input
rlabel viali s 1225 43503 1259 43537 6 VPWR
port 613 nsew power input
rlabel viali s 1133 43503 1167 43537 6 VPWR
port 613 nsew power input
rlabel viali s 298753 44591 298787 44625 6 VPWR
port 613 nsew power input
rlabel viali s 298661 44591 298695 44625 6 VPWR
port 613 nsew power input
rlabel viali s 1317 44591 1340 44625 6 VPWR
port 613 nsew power input
rlabel viali s 1225 44591 1259 44625 6 VPWR
port 613 nsew power input
rlabel viali s 1133 44591 1167 44625 6 VPWR
port 613 nsew power input
rlabel viali s 298753 45679 298787 45713 6 VPWR
port 613 nsew power input
rlabel viali s 298661 45679 298695 45713 6 VPWR
port 613 nsew power input
rlabel viali s 1317 45679 1340 45713 6 VPWR
port 613 nsew power input
rlabel viali s 1225 45679 1259 45713 6 VPWR
port 613 nsew power input
rlabel viali s 1133 45679 1167 45713 6 VPWR
port 613 nsew power input
rlabel viali s 298753 46767 298787 46801 6 VPWR
port 613 nsew power input
rlabel viali s 298661 46767 298695 46801 6 VPWR
port 613 nsew power input
rlabel viali s 1317 46767 1340 46801 6 VPWR
port 613 nsew power input
rlabel viali s 1225 46767 1259 46801 6 VPWR
port 613 nsew power input
rlabel viali s 1133 46767 1167 46801 6 VPWR
port 613 nsew power input
rlabel viali s 298753 47855 298787 47889 6 VPWR
port 613 nsew power input
rlabel viali s 298661 47855 298695 47889 6 VPWR
port 613 nsew power input
rlabel viali s 1317 47855 1340 47889 6 VPWR
port 613 nsew power input
rlabel viali s 1225 47855 1259 47889 6 VPWR
port 613 nsew power input
rlabel viali s 1133 47855 1167 47889 6 VPWR
port 613 nsew power input
rlabel viali s 298753 48943 298787 48977 6 VPWR
port 613 nsew power input
rlabel viali s 298661 48943 298695 48977 6 VPWR
port 613 nsew power input
rlabel viali s 1317 48943 1340 48977 6 VPWR
port 613 nsew power input
rlabel viali s 1225 48943 1259 48977 6 VPWR
port 613 nsew power input
rlabel viali s 1133 48943 1167 48977 6 VPWR
port 613 nsew power input
rlabel viali s 298753 50031 298787 50065 6 VPWR
port 613 nsew power input
rlabel viali s 298661 50031 298695 50065 6 VPWR
port 613 nsew power input
rlabel viali s 1317 50031 1340 50065 6 VPWR
port 613 nsew power input
rlabel viali s 1225 50031 1259 50065 6 VPWR
port 613 nsew power input
rlabel viali s 1133 50031 1167 50065 6 VPWR
port 613 nsew power input
rlabel viali s 298753 51119 298787 51153 6 VPWR
port 613 nsew power input
rlabel viali s 298661 51119 298695 51153 6 VPWR
port 613 nsew power input
rlabel viali s 1317 51119 1340 51153 6 VPWR
port 613 nsew power input
rlabel viali s 1225 51119 1259 51153 6 VPWR
port 613 nsew power input
rlabel viali s 1133 51119 1167 51153 6 VPWR
port 613 nsew power input
rlabel viali s 298753 52207 298787 52241 6 VPWR
port 613 nsew power input
rlabel viali s 298661 52207 298695 52241 6 VPWR
port 613 nsew power input
rlabel viali s 1317 52207 1340 52241 6 VPWR
port 613 nsew power input
rlabel viali s 1225 52207 1259 52241 6 VPWR
port 613 nsew power input
rlabel viali s 1133 52207 1167 52241 6 VPWR
port 613 nsew power input
rlabel viali s 298753 53295 298787 53329 6 VPWR
port 613 nsew power input
rlabel viali s 298661 53295 298695 53329 6 VPWR
port 613 nsew power input
rlabel viali s 1317 53295 1340 53329 6 VPWR
port 613 nsew power input
rlabel viali s 1225 53295 1259 53329 6 VPWR
port 613 nsew power input
rlabel viali s 1133 53295 1167 53329 6 VPWR
port 613 nsew power input
rlabel viali s 298753 54383 298787 54417 6 VPWR
port 613 nsew power input
rlabel viali s 298661 54383 298695 54417 6 VPWR
port 613 nsew power input
rlabel viali s 1317 54383 1340 54417 6 VPWR
port 613 nsew power input
rlabel viali s 1225 54383 1259 54417 6 VPWR
port 613 nsew power input
rlabel viali s 1133 54383 1167 54417 6 VPWR
port 613 nsew power input
rlabel viali s 298753 55471 298787 55505 6 VPWR
port 613 nsew power input
rlabel viali s 298661 55471 298695 55505 6 VPWR
port 613 nsew power input
rlabel viali s 1317 55471 1340 55505 6 VPWR
port 613 nsew power input
rlabel viali s 1225 55471 1259 55505 6 VPWR
port 613 nsew power input
rlabel viali s 1133 55471 1167 55505 6 VPWR
port 613 nsew power input
rlabel viali s 298753 56559 298787 56593 6 VPWR
port 613 nsew power input
rlabel viali s 298661 56559 298695 56593 6 VPWR
port 613 nsew power input
rlabel viali s 1317 56559 1340 56593 6 VPWR
port 613 nsew power input
rlabel viali s 1225 56559 1259 56593 6 VPWR
port 613 nsew power input
rlabel viali s 1133 56559 1167 56593 6 VPWR
port 613 nsew power input
rlabel viali s 298753 57647 298787 57681 6 VPWR
port 613 nsew power input
rlabel viali s 298661 57647 298695 57681 6 VPWR
port 613 nsew power input
rlabel viali s 1317 57647 1340 57681 6 VPWR
port 613 nsew power input
rlabel viali s 1225 57647 1259 57681 6 VPWR
port 613 nsew power input
rlabel viali s 1133 57647 1167 57681 6 VPWR
port 613 nsew power input
rlabel viali s 298753 58735 298787 58769 6 VPWR
port 613 nsew power input
rlabel viali s 298661 58735 298695 58769 6 VPWR
port 613 nsew power input
rlabel viali s 1317 58735 1340 58769 6 VPWR
port 613 nsew power input
rlabel viali s 1225 58735 1259 58769 6 VPWR
port 613 nsew power input
rlabel viali s 1133 58735 1167 58769 6 VPWR
port 613 nsew power input
rlabel viali s 298753 59823 298787 59857 6 VPWR
port 613 nsew power input
rlabel viali s 298661 59823 298695 59857 6 VPWR
port 613 nsew power input
rlabel viali s 1317 59823 1340 59857 6 VPWR
port 613 nsew power input
rlabel viali s 1225 59823 1259 59857 6 VPWR
port 613 nsew power input
rlabel viali s 1133 59823 1167 59857 6 VPWR
port 613 nsew power input
rlabel viali s 298753 60911 298787 60945 6 VPWR
port 613 nsew power input
rlabel viali s 298661 60911 298695 60945 6 VPWR
port 613 nsew power input
rlabel viali s 1317 60911 1340 60945 6 VPWR
port 613 nsew power input
rlabel viali s 1225 60911 1259 60945 6 VPWR
port 613 nsew power input
rlabel viali s 1133 60911 1167 60945 6 VPWR
port 613 nsew power input
rlabel viali s 298753 61999 298787 62033 6 VPWR
port 613 nsew power input
rlabel viali s 298661 61999 298695 62033 6 VPWR
port 613 nsew power input
rlabel viali s 1317 61999 1340 62033 6 VPWR
port 613 nsew power input
rlabel viali s 1225 61999 1259 62033 6 VPWR
port 613 nsew power input
rlabel viali s 1133 61999 1167 62033 6 VPWR
port 613 nsew power input
rlabel viali s 298753 63087 298787 63121 6 VPWR
port 613 nsew power input
rlabel viali s 298661 63087 298695 63121 6 VPWR
port 613 nsew power input
rlabel viali s 1317 63087 1340 63121 6 VPWR
port 613 nsew power input
rlabel viali s 1225 63087 1259 63121 6 VPWR
port 613 nsew power input
rlabel viali s 1133 63087 1167 63121 6 VPWR
port 613 nsew power input
rlabel viali s 298753 64175 298787 64209 6 VPWR
port 613 nsew power input
rlabel viali s 298661 64175 298695 64209 6 VPWR
port 613 nsew power input
rlabel viali s 1317 64175 1340 64209 6 VPWR
port 613 nsew power input
rlabel viali s 1225 64175 1259 64209 6 VPWR
port 613 nsew power input
rlabel viali s 1133 64175 1167 64209 6 VPWR
port 613 nsew power input
rlabel viali s 298753 65263 298787 65297 6 VPWR
port 613 nsew power input
rlabel viali s 298661 65263 298695 65297 6 VPWR
port 613 nsew power input
rlabel viali s 1317 65263 1340 65297 6 VPWR
port 613 nsew power input
rlabel viali s 1225 65263 1259 65297 6 VPWR
port 613 nsew power input
rlabel viali s 1133 65263 1167 65297 6 VPWR
port 613 nsew power input
rlabel viali s 298753 66351 298787 66385 6 VPWR
port 613 nsew power input
rlabel viali s 298661 66351 298695 66385 6 VPWR
port 613 nsew power input
rlabel viali s 1317 66351 1340 66385 6 VPWR
port 613 nsew power input
rlabel viali s 1225 66351 1259 66385 6 VPWR
port 613 nsew power input
rlabel viali s 1133 66351 1167 66385 6 VPWR
port 613 nsew power input
rlabel viali s 298753 67439 298787 67473 6 VPWR
port 613 nsew power input
rlabel viali s 298661 67439 298695 67473 6 VPWR
port 613 nsew power input
rlabel viali s 1317 67439 1340 67473 6 VPWR
port 613 nsew power input
rlabel viali s 1225 67439 1259 67473 6 VPWR
port 613 nsew power input
rlabel viali s 1133 67439 1167 67473 6 VPWR
port 613 nsew power input
rlabel viali s 298753 68527 298787 68561 6 VPWR
port 613 nsew power input
rlabel viali s 298661 68527 298695 68561 6 VPWR
port 613 nsew power input
rlabel viali s 1317 68527 1340 68561 6 VPWR
port 613 nsew power input
rlabel viali s 1225 68527 1259 68561 6 VPWR
port 613 nsew power input
rlabel viali s 1133 68527 1167 68561 6 VPWR
port 613 nsew power input
rlabel viali s 298753 69615 298787 69649 6 VPWR
port 613 nsew power input
rlabel viali s 298661 69615 298695 69649 6 VPWR
port 613 nsew power input
rlabel viali s 1317 69615 1340 69649 6 VPWR
port 613 nsew power input
rlabel viali s 1225 69615 1259 69649 6 VPWR
port 613 nsew power input
rlabel viali s 1133 69615 1167 69649 6 VPWR
port 613 nsew power input
rlabel viali s 298753 70703 298787 70737 6 VPWR
port 613 nsew power input
rlabel viali s 298661 70703 298695 70737 6 VPWR
port 613 nsew power input
rlabel viali s 1317 70703 1340 70737 6 VPWR
port 613 nsew power input
rlabel viali s 1225 70703 1259 70737 6 VPWR
port 613 nsew power input
rlabel viali s 1133 70703 1167 70737 6 VPWR
port 613 nsew power input
rlabel viali s 298753 71791 298787 71825 6 VPWR
port 613 nsew power input
rlabel viali s 298661 71791 298695 71825 6 VPWR
port 613 nsew power input
rlabel viali s 1317 71791 1340 71825 6 VPWR
port 613 nsew power input
rlabel viali s 1225 71791 1259 71825 6 VPWR
port 613 nsew power input
rlabel viali s 1133 71791 1167 71825 6 VPWR
port 613 nsew power input
rlabel viali s 298753 72879 298787 72913 6 VPWR
port 613 nsew power input
rlabel viali s 298661 72879 298695 72913 6 VPWR
port 613 nsew power input
rlabel viali s 1317 72879 1340 72913 6 VPWR
port 613 nsew power input
rlabel viali s 1225 72879 1259 72913 6 VPWR
port 613 nsew power input
rlabel viali s 1133 72879 1167 72913 6 VPWR
port 613 nsew power input
rlabel viali s 298753 73967 298787 74001 6 VPWR
port 613 nsew power input
rlabel viali s 298661 73967 298695 74001 6 VPWR
port 613 nsew power input
rlabel viali s 1317 73967 1340 74001 6 VPWR
port 613 nsew power input
rlabel viali s 1225 73967 1259 74001 6 VPWR
port 613 nsew power input
rlabel viali s 1133 73967 1167 74001 6 VPWR
port 613 nsew power input
rlabel viali s 298753 75055 298787 75089 6 VPWR
port 613 nsew power input
rlabel viali s 298661 75055 298695 75089 6 VPWR
port 613 nsew power input
rlabel viali s 1317 75055 1340 75089 6 VPWR
port 613 nsew power input
rlabel viali s 1225 75055 1259 75089 6 VPWR
port 613 nsew power input
rlabel viali s 1133 75055 1167 75089 6 VPWR
port 613 nsew power input
rlabel viali s 298753 76143 298787 76177 6 VPWR
port 613 nsew power input
rlabel viali s 298661 76143 298695 76177 6 VPWR
port 613 nsew power input
rlabel viali s 1317 76143 1340 76177 6 VPWR
port 613 nsew power input
rlabel viali s 1225 76143 1259 76177 6 VPWR
port 613 nsew power input
rlabel viali s 1133 76143 1167 76177 6 VPWR
port 613 nsew power input
rlabel viali s 298753 77231 298787 77265 6 VPWR
port 613 nsew power input
rlabel viali s 298661 77231 298695 77265 6 VPWR
port 613 nsew power input
rlabel viali s 1317 77231 1340 77265 6 VPWR
port 613 nsew power input
rlabel viali s 1225 77231 1259 77265 6 VPWR
port 613 nsew power input
rlabel viali s 1133 77231 1167 77265 6 VPWR
port 613 nsew power input
rlabel viali s 298753 78319 298787 78353 6 VPWR
port 613 nsew power input
rlabel viali s 298661 78319 298695 78353 6 VPWR
port 613 nsew power input
rlabel viali s 1317 78319 1340 78353 6 VPWR
port 613 nsew power input
rlabel viali s 1225 78319 1259 78353 6 VPWR
port 613 nsew power input
rlabel viali s 1133 78319 1167 78353 6 VPWR
port 613 nsew power input
rlabel viali s 298753 79407 298787 79441 6 VPWR
port 613 nsew power input
rlabel viali s 298661 79407 298695 79441 6 VPWR
port 613 nsew power input
rlabel viali s 1317 79407 1340 79441 6 VPWR
port 613 nsew power input
rlabel viali s 1225 79407 1259 79441 6 VPWR
port 613 nsew power input
rlabel viali s 1133 79407 1167 79441 6 VPWR
port 613 nsew power input
rlabel viali s 298753 80495 298787 80529 6 VPWR
port 613 nsew power input
rlabel viali s 298661 80495 298695 80529 6 VPWR
port 613 nsew power input
rlabel viali s 1317 80495 1340 80529 6 VPWR
port 613 nsew power input
rlabel viali s 1225 80495 1259 80529 6 VPWR
port 613 nsew power input
rlabel viali s 1133 80495 1167 80529 6 VPWR
port 613 nsew power input
rlabel viali s 298753 81583 298787 81617 6 VPWR
port 613 nsew power input
rlabel viali s 298661 81583 298695 81617 6 VPWR
port 613 nsew power input
rlabel viali s 1317 81583 1340 81617 6 VPWR
port 613 nsew power input
rlabel viali s 1225 81583 1259 81617 6 VPWR
port 613 nsew power input
rlabel viali s 1133 81583 1167 81617 6 VPWR
port 613 nsew power input
rlabel viali s 298753 82671 298787 82705 6 VPWR
port 613 nsew power input
rlabel viali s 298661 82671 298695 82705 6 VPWR
port 613 nsew power input
rlabel viali s 1317 82671 1340 82705 6 VPWR
port 613 nsew power input
rlabel viali s 1225 82671 1259 82705 6 VPWR
port 613 nsew power input
rlabel viali s 1133 82671 1167 82705 6 VPWR
port 613 nsew power input
rlabel viali s 298753 83759 298787 83793 6 VPWR
port 613 nsew power input
rlabel viali s 298661 83759 298695 83793 6 VPWR
port 613 nsew power input
rlabel viali s 1317 83759 1340 83793 6 VPWR
port 613 nsew power input
rlabel viali s 1225 83759 1259 83793 6 VPWR
port 613 nsew power input
rlabel viali s 1133 83759 1167 83793 6 VPWR
port 613 nsew power input
rlabel viali s 298753 84847 298787 84881 6 VPWR
port 613 nsew power input
rlabel viali s 298661 84847 298695 84881 6 VPWR
port 613 nsew power input
rlabel viali s 1317 84847 1340 84881 6 VPWR
port 613 nsew power input
rlabel viali s 1225 84847 1259 84881 6 VPWR
port 613 nsew power input
rlabel viali s 1133 84847 1167 84881 6 VPWR
port 613 nsew power input
rlabel viali s 298753 85935 298787 85969 6 VPWR
port 613 nsew power input
rlabel viali s 298661 85935 298695 85969 6 VPWR
port 613 nsew power input
rlabel viali s 1317 85935 1340 85969 6 VPWR
port 613 nsew power input
rlabel viali s 1225 85935 1259 85969 6 VPWR
port 613 nsew power input
rlabel viali s 1133 85935 1167 85969 6 VPWR
port 613 nsew power input
rlabel viali s 298753 87023 298787 87057 6 VPWR
port 613 nsew power input
rlabel viali s 298661 87023 298695 87057 6 VPWR
port 613 nsew power input
rlabel viali s 1317 87023 1340 87057 6 VPWR
port 613 nsew power input
rlabel viali s 1225 87023 1259 87057 6 VPWR
port 613 nsew power input
rlabel viali s 1133 87023 1167 87057 6 VPWR
port 613 nsew power input
rlabel viali s 298753 88111 298787 88145 6 VPWR
port 613 nsew power input
rlabel viali s 298661 88111 298695 88145 6 VPWR
port 613 nsew power input
rlabel viali s 1317 88111 1340 88145 6 VPWR
port 613 nsew power input
rlabel viali s 1225 88111 1259 88145 6 VPWR
port 613 nsew power input
rlabel viali s 1133 88111 1167 88145 6 VPWR
port 613 nsew power input
rlabel viali s 298753 89199 298787 89233 6 VPWR
port 613 nsew power input
rlabel viali s 298661 89199 298695 89233 6 VPWR
port 613 nsew power input
rlabel viali s 1317 89199 1340 89233 6 VPWR
port 613 nsew power input
rlabel viali s 1225 89199 1259 89233 6 VPWR
port 613 nsew power input
rlabel viali s 1133 89199 1167 89233 6 VPWR
port 613 nsew power input
rlabel viali s 298753 90287 298787 90321 6 VPWR
port 613 nsew power input
rlabel viali s 298661 90287 298695 90321 6 VPWR
port 613 nsew power input
rlabel viali s 1317 90287 1340 90321 6 VPWR
port 613 nsew power input
rlabel viali s 1225 90287 1259 90321 6 VPWR
port 613 nsew power input
rlabel viali s 1133 90287 1167 90321 6 VPWR
port 613 nsew power input
rlabel viali s 298753 91375 298787 91409 6 VPWR
port 613 nsew power input
rlabel viali s 298661 91375 298695 91409 6 VPWR
port 613 nsew power input
rlabel viali s 1317 91375 1340 91409 6 VPWR
port 613 nsew power input
rlabel viali s 1225 91375 1259 91409 6 VPWR
port 613 nsew power input
rlabel viali s 1133 91375 1167 91409 6 VPWR
port 613 nsew power input
rlabel viali s 298753 92463 298787 92497 6 VPWR
port 613 nsew power input
rlabel viali s 298661 92463 298695 92497 6 VPWR
port 613 nsew power input
rlabel viali s 1317 92463 1340 92497 6 VPWR
port 613 nsew power input
rlabel viali s 1225 92463 1259 92497 6 VPWR
port 613 nsew power input
rlabel viali s 1133 92463 1167 92497 6 VPWR
port 613 nsew power input
rlabel viali s 298753 93551 298787 93585 6 VPWR
port 613 nsew power input
rlabel viali s 298661 93551 298695 93585 6 VPWR
port 613 nsew power input
rlabel viali s 1317 93551 1340 93585 6 VPWR
port 613 nsew power input
rlabel viali s 1225 93551 1259 93585 6 VPWR
port 613 nsew power input
rlabel viali s 1133 93551 1167 93585 6 VPWR
port 613 nsew power input
rlabel viali s 298753 94639 298787 94673 6 VPWR
port 613 nsew power input
rlabel viali s 298661 94639 298695 94673 6 VPWR
port 613 nsew power input
rlabel viali s 1317 94639 1340 94673 6 VPWR
port 613 nsew power input
rlabel viali s 1225 94639 1259 94673 6 VPWR
port 613 nsew power input
rlabel viali s 1133 94639 1167 94673 6 VPWR
port 613 nsew power input
rlabel viali s 298753 95727 298787 95761 6 VPWR
port 613 nsew power input
rlabel viali s 298661 95727 298695 95761 6 VPWR
port 613 nsew power input
rlabel viali s 1317 95727 1340 95761 6 VPWR
port 613 nsew power input
rlabel viali s 1225 95727 1259 95761 6 VPWR
port 613 nsew power input
rlabel viali s 1133 95727 1167 95761 6 VPWR
port 613 nsew power input
rlabel viali s 298753 96815 298787 96849 6 VPWR
port 613 nsew power input
rlabel viali s 298661 96815 298695 96849 6 VPWR
port 613 nsew power input
rlabel viali s 1317 96815 1340 96849 6 VPWR
port 613 nsew power input
rlabel viali s 1225 96815 1259 96849 6 VPWR
port 613 nsew power input
rlabel viali s 1133 96815 1167 96849 6 VPWR
port 613 nsew power input
rlabel viali s 298753 97903 298787 97937 6 VPWR
port 613 nsew power input
rlabel viali s 298661 97903 298695 97937 6 VPWR
port 613 nsew power input
rlabel viali s 1317 97903 1340 97937 6 VPWR
port 613 nsew power input
rlabel viali s 1225 97903 1259 97937 6 VPWR
port 613 nsew power input
rlabel viali s 1133 97903 1167 97937 6 VPWR
port 613 nsew power input
rlabel viali s 298753 98991 298787 99025 6 VPWR
port 613 nsew power input
rlabel viali s 298661 98991 298695 99025 6 VPWR
port 613 nsew power input
rlabel viali s 1317 98991 1340 99025 6 VPWR
port 613 nsew power input
rlabel viali s 1225 98991 1259 99025 6 VPWR
port 613 nsew power input
rlabel viali s 1133 98991 1167 99025 6 VPWR
port 613 nsew power input
rlabel viali s 298753 100079 298787 100113 6 VPWR
port 613 nsew power input
rlabel viali s 298661 100079 298695 100113 6 VPWR
port 613 nsew power input
rlabel viali s 1317 100079 1340 100113 6 VPWR
port 613 nsew power input
rlabel viali s 1225 100079 1259 100113 6 VPWR
port 613 nsew power input
rlabel viali s 1133 100079 1167 100113 6 VPWR
port 613 nsew power input
rlabel viali s 298753 101167 298787 101201 6 VPWR
port 613 nsew power input
rlabel viali s 298661 101167 298695 101201 6 VPWR
port 613 nsew power input
rlabel viali s 1317 101167 1340 101201 6 VPWR
port 613 nsew power input
rlabel viali s 1225 101167 1259 101201 6 VPWR
port 613 nsew power input
rlabel viali s 1133 101167 1167 101201 6 VPWR
port 613 nsew power input
rlabel viali s 298753 102255 298787 102289 6 VPWR
port 613 nsew power input
rlabel viali s 298661 102255 298695 102289 6 VPWR
port 613 nsew power input
rlabel viali s 1317 102255 1340 102289 6 VPWR
port 613 nsew power input
rlabel viali s 1225 102255 1259 102289 6 VPWR
port 613 nsew power input
rlabel viali s 1133 102255 1167 102289 6 VPWR
port 613 nsew power input
rlabel viali s 298753 103343 298787 103377 6 VPWR
port 613 nsew power input
rlabel viali s 298661 103343 298695 103377 6 VPWR
port 613 nsew power input
rlabel viali s 1317 103343 1340 103377 6 VPWR
port 613 nsew power input
rlabel viali s 1225 103343 1259 103377 6 VPWR
port 613 nsew power input
rlabel viali s 1133 103343 1167 103377 6 VPWR
port 613 nsew power input
rlabel viali s 298753 104431 298787 104465 6 VPWR
port 613 nsew power input
rlabel viali s 298661 104431 298695 104465 6 VPWR
port 613 nsew power input
rlabel viali s 1317 104431 1340 104465 6 VPWR
port 613 nsew power input
rlabel viali s 1225 104431 1259 104465 6 VPWR
port 613 nsew power input
rlabel viali s 1133 104431 1167 104465 6 VPWR
port 613 nsew power input
rlabel viali s 298753 105519 298787 105553 6 VPWR
port 613 nsew power input
rlabel viali s 298661 105519 298695 105553 6 VPWR
port 613 nsew power input
rlabel viali s 1317 105519 1340 105553 6 VPWR
port 613 nsew power input
rlabel viali s 1225 105519 1259 105553 6 VPWR
port 613 nsew power input
rlabel viali s 1133 105519 1167 105553 6 VPWR
port 613 nsew power input
rlabel viali s 298753 106607 298787 106641 6 VPWR
port 613 nsew power input
rlabel viali s 298661 106607 298695 106641 6 VPWR
port 613 nsew power input
rlabel viali s 1317 106607 1340 106641 6 VPWR
port 613 nsew power input
rlabel viali s 1225 106607 1259 106641 6 VPWR
port 613 nsew power input
rlabel viali s 1133 106607 1167 106641 6 VPWR
port 613 nsew power input
rlabel viali s 298753 107695 298787 107729 6 VPWR
port 613 nsew power input
rlabel viali s 298661 107695 298695 107729 6 VPWR
port 613 nsew power input
rlabel viali s 1317 107695 1340 107729 6 VPWR
port 613 nsew power input
rlabel viali s 1225 107695 1259 107729 6 VPWR
port 613 nsew power input
rlabel viali s 1133 107695 1167 107729 6 VPWR
port 613 nsew power input
rlabel viali s 298753 108783 298787 108817 6 VPWR
port 613 nsew power input
rlabel viali s 298661 108783 298695 108817 6 VPWR
port 613 nsew power input
rlabel viali s 1317 108783 1340 108817 6 VPWR
port 613 nsew power input
rlabel viali s 1225 108783 1259 108817 6 VPWR
port 613 nsew power input
rlabel viali s 1133 108783 1167 108817 6 VPWR
port 613 nsew power input
rlabel viali s 298753 109871 298787 109905 6 VPWR
port 613 nsew power input
rlabel viali s 298661 109871 298695 109905 6 VPWR
port 613 nsew power input
rlabel viali s 1317 109871 1340 109905 6 VPWR
port 613 nsew power input
rlabel viali s 1225 109871 1259 109905 6 VPWR
port 613 nsew power input
rlabel viali s 1133 109871 1167 109905 6 VPWR
port 613 nsew power input
rlabel viali s 298753 110959 298787 110993 6 VPWR
port 613 nsew power input
rlabel viali s 298661 110959 298695 110993 6 VPWR
port 613 nsew power input
rlabel viali s 1317 110959 1340 110993 6 VPWR
port 613 nsew power input
rlabel viali s 1225 110959 1259 110993 6 VPWR
port 613 nsew power input
rlabel viali s 1133 110959 1167 110993 6 VPWR
port 613 nsew power input
rlabel viali s 298753 112047 298787 112081 6 VPWR
port 613 nsew power input
rlabel viali s 298661 112047 298695 112081 6 VPWR
port 613 nsew power input
rlabel viali s 1317 112047 1340 112081 6 VPWR
port 613 nsew power input
rlabel viali s 1225 112047 1259 112081 6 VPWR
port 613 nsew power input
rlabel viali s 1133 112047 1167 112081 6 VPWR
port 613 nsew power input
rlabel viali s 298753 113135 298787 113169 6 VPWR
port 613 nsew power input
rlabel viali s 298661 113135 298695 113169 6 VPWR
port 613 nsew power input
rlabel viali s 1317 113135 1340 113169 6 VPWR
port 613 nsew power input
rlabel viali s 1225 113135 1259 113169 6 VPWR
port 613 nsew power input
rlabel viali s 1133 113135 1167 113169 6 VPWR
port 613 nsew power input
rlabel viali s 298753 114223 298787 114257 6 VPWR
port 613 nsew power input
rlabel viali s 298661 114223 298695 114257 6 VPWR
port 613 nsew power input
rlabel viali s 1317 114223 1340 114257 6 VPWR
port 613 nsew power input
rlabel viali s 1225 114223 1259 114257 6 VPWR
port 613 nsew power input
rlabel viali s 1133 114223 1167 114257 6 VPWR
port 613 nsew power input
rlabel viali s 298753 115311 298787 115345 6 VPWR
port 613 nsew power input
rlabel viali s 298661 115311 298695 115345 6 VPWR
port 613 nsew power input
rlabel viali s 1317 115311 1340 115345 6 VPWR
port 613 nsew power input
rlabel viali s 1225 115311 1259 115345 6 VPWR
port 613 nsew power input
rlabel viali s 1133 115311 1167 115345 6 VPWR
port 613 nsew power input
rlabel viali s 298753 116399 298787 116433 6 VPWR
port 613 nsew power input
rlabel viali s 298661 116399 298695 116433 6 VPWR
port 613 nsew power input
rlabel viali s 1317 116399 1340 116433 6 VPWR
port 613 nsew power input
rlabel viali s 1225 116399 1259 116433 6 VPWR
port 613 nsew power input
rlabel viali s 1133 116399 1167 116433 6 VPWR
port 613 nsew power input
rlabel viali s 298753 117487 298787 117521 6 VPWR
port 613 nsew power input
rlabel viali s 298661 117487 298695 117521 6 VPWR
port 613 nsew power input
rlabel viali s 1317 117487 1340 117521 6 VPWR
port 613 nsew power input
rlabel viali s 1225 117487 1259 117521 6 VPWR
port 613 nsew power input
rlabel viali s 1133 117487 1167 117521 6 VPWR
port 613 nsew power input
rlabel viali s 298753 118575 298787 118609 6 VPWR
port 613 nsew power input
rlabel viali s 298661 118575 298695 118609 6 VPWR
port 613 nsew power input
rlabel viali s 1317 118575 1340 118609 6 VPWR
port 613 nsew power input
rlabel viali s 1225 118575 1259 118609 6 VPWR
port 613 nsew power input
rlabel viali s 1133 118575 1167 118609 6 VPWR
port 613 nsew power input
rlabel viali s 298753 119663 298787 119697 6 VPWR
port 613 nsew power input
rlabel viali s 298661 119663 298695 119697 6 VPWR
port 613 nsew power input
rlabel viali s 1317 119663 1340 119697 6 VPWR
port 613 nsew power input
rlabel viali s 1225 119663 1259 119697 6 VPWR
port 613 nsew power input
rlabel viali s 1133 119663 1167 119697 6 VPWR
port 613 nsew power input
rlabel viali s 298753 120751 298787 120785 6 VPWR
port 613 nsew power input
rlabel viali s 298661 120751 298695 120785 6 VPWR
port 613 nsew power input
rlabel viali s 1317 120751 1340 120785 6 VPWR
port 613 nsew power input
rlabel viali s 1225 120751 1259 120785 6 VPWR
port 613 nsew power input
rlabel viali s 1133 120751 1167 120785 6 VPWR
port 613 nsew power input
rlabel viali s 298753 121839 298787 121873 6 VPWR
port 613 nsew power input
rlabel viali s 298661 121839 298695 121873 6 VPWR
port 613 nsew power input
rlabel viali s 1317 121839 1340 121873 6 VPWR
port 613 nsew power input
rlabel viali s 1225 121839 1259 121873 6 VPWR
port 613 nsew power input
rlabel viali s 1133 121839 1167 121873 6 VPWR
port 613 nsew power input
rlabel viali s 298753 122927 298787 122961 6 VPWR
port 613 nsew power input
rlabel viali s 298661 122927 298695 122961 6 VPWR
port 613 nsew power input
rlabel viali s 1317 122927 1340 122961 6 VPWR
port 613 nsew power input
rlabel viali s 1225 122927 1259 122961 6 VPWR
port 613 nsew power input
rlabel viali s 1133 122927 1167 122961 6 VPWR
port 613 nsew power input
rlabel viali s 298753 124015 298787 124049 6 VPWR
port 613 nsew power input
rlabel viali s 298661 124015 298695 124049 6 VPWR
port 613 nsew power input
rlabel viali s 1317 124015 1340 124049 6 VPWR
port 613 nsew power input
rlabel viali s 1225 124015 1259 124049 6 VPWR
port 613 nsew power input
rlabel viali s 1133 124015 1167 124049 6 VPWR
port 613 nsew power input
rlabel viali s 298753 125103 298787 125137 6 VPWR
port 613 nsew power input
rlabel viali s 298661 125103 298695 125137 6 VPWR
port 613 nsew power input
rlabel viali s 1317 125103 1340 125137 6 VPWR
port 613 nsew power input
rlabel viali s 1225 125103 1259 125137 6 VPWR
port 613 nsew power input
rlabel viali s 1133 125103 1167 125137 6 VPWR
port 613 nsew power input
rlabel viali s 298753 126191 298787 126225 6 VPWR
port 613 nsew power input
rlabel viali s 298661 126191 298695 126225 6 VPWR
port 613 nsew power input
rlabel viali s 1317 126191 1340 126225 6 VPWR
port 613 nsew power input
rlabel viali s 1225 126191 1259 126225 6 VPWR
port 613 nsew power input
rlabel viali s 1133 126191 1167 126225 6 VPWR
port 613 nsew power input
rlabel viali s 298753 127279 298787 127313 6 VPWR
port 613 nsew power input
rlabel viali s 298661 127279 298695 127313 6 VPWR
port 613 nsew power input
rlabel viali s 1317 127279 1340 127313 6 VPWR
port 613 nsew power input
rlabel viali s 1225 127279 1259 127313 6 VPWR
port 613 nsew power input
rlabel viali s 1133 127279 1167 127313 6 VPWR
port 613 nsew power input
rlabel viali s 298753 128367 298787 128401 6 VPWR
port 613 nsew power input
rlabel viali s 298661 128367 298695 128401 6 VPWR
port 613 nsew power input
rlabel viali s 1317 128367 1340 128401 6 VPWR
port 613 nsew power input
rlabel viali s 1225 128367 1259 128401 6 VPWR
port 613 nsew power input
rlabel viali s 1133 128367 1167 128401 6 VPWR
port 613 nsew power input
rlabel viali s 298753 129455 298787 129489 6 VPWR
port 613 nsew power input
rlabel viali s 298661 129455 298695 129489 6 VPWR
port 613 nsew power input
rlabel viali s 1317 129455 1340 129489 6 VPWR
port 613 nsew power input
rlabel viali s 1225 129455 1259 129489 6 VPWR
port 613 nsew power input
rlabel viali s 1133 129455 1167 129489 6 VPWR
port 613 nsew power input
rlabel viali s 298753 130543 298787 130577 6 VPWR
port 613 nsew power input
rlabel viali s 298661 130543 298695 130577 6 VPWR
port 613 nsew power input
rlabel viali s 1317 130543 1340 130577 6 VPWR
port 613 nsew power input
rlabel viali s 1225 130543 1259 130577 6 VPWR
port 613 nsew power input
rlabel viali s 1133 130543 1167 130577 6 VPWR
port 613 nsew power input
rlabel viali s 298753 131631 298787 131665 6 VPWR
port 613 nsew power input
rlabel viali s 298661 131631 298695 131665 6 VPWR
port 613 nsew power input
rlabel viali s 1317 131631 1340 131665 6 VPWR
port 613 nsew power input
rlabel viali s 1225 131631 1259 131665 6 VPWR
port 613 nsew power input
rlabel viali s 1133 131631 1167 131665 6 VPWR
port 613 nsew power input
rlabel viali s 298753 132719 298787 132753 6 VPWR
port 613 nsew power input
rlabel viali s 298661 132719 298695 132753 6 VPWR
port 613 nsew power input
rlabel viali s 1317 132719 1340 132753 6 VPWR
port 613 nsew power input
rlabel viali s 1225 132719 1259 132753 6 VPWR
port 613 nsew power input
rlabel viali s 1133 132719 1167 132753 6 VPWR
port 613 nsew power input
rlabel viali s 298753 133807 298787 133841 6 VPWR
port 613 nsew power input
rlabel viali s 298661 133807 298695 133841 6 VPWR
port 613 nsew power input
rlabel viali s 1317 133807 1340 133841 6 VPWR
port 613 nsew power input
rlabel viali s 1225 133807 1259 133841 6 VPWR
port 613 nsew power input
rlabel viali s 1133 133807 1167 133841 6 VPWR
port 613 nsew power input
rlabel viali s 298753 134895 298787 134929 6 VPWR
port 613 nsew power input
rlabel viali s 298661 134895 298695 134929 6 VPWR
port 613 nsew power input
rlabel viali s 1317 134895 1340 134929 6 VPWR
port 613 nsew power input
rlabel viali s 1225 134895 1259 134929 6 VPWR
port 613 nsew power input
rlabel viali s 1133 134895 1167 134929 6 VPWR
port 613 nsew power input
rlabel viali s 298753 135983 298787 136017 6 VPWR
port 613 nsew power input
rlabel viali s 298661 135983 298695 136017 6 VPWR
port 613 nsew power input
rlabel viali s 1317 135983 1340 136017 6 VPWR
port 613 nsew power input
rlabel viali s 1225 135983 1259 136017 6 VPWR
port 613 nsew power input
rlabel viali s 1133 135983 1167 136017 6 VPWR
port 613 nsew power input
rlabel viali s 298753 137071 298787 137105 6 VPWR
port 613 nsew power input
rlabel viali s 298661 137071 298695 137105 6 VPWR
port 613 nsew power input
rlabel viali s 1317 137071 1340 137105 6 VPWR
port 613 nsew power input
rlabel viali s 1225 137071 1259 137105 6 VPWR
port 613 nsew power input
rlabel viali s 1133 137071 1167 137105 6 VPWR
port 613 nsew power input
rlabel viali s 298753 138159 298787 138193 6 VPWR
port 613 nsew power input
rlabel viali s 298661 138159 298695 138193 6 VPWR
port 613 nsew power input
rlabel viali s 1317 138159 1340 138193 6 VPWR
port 613 nsew power input
rlabel viali s 1225 138159 1259 138193 6 VPWR
port 613 nsew power input
rlabel viali s 1133 138159 1167 138193 6 VPWR
port 613 nsew power input
rlabel viali s 298753 139247 298787 139281 6 VPWR
port 613 nsew power input
rlabel viali s 298661 139247 298695 139281 6 VPWR
port 613 nsew power input
rlabel viali s 1317 139247 1340 139281 6 VPWR
port 613 nsew power input
rlabel viali s 1225 139247 1259 139281 6 VPWR
port 613 nsew power input
rlabel viali s 1133 139247 1167 139281 6 VPWR
port 613 nsew power input
rlabel viali s 298753 140335 298787 140369 6 VPWR
port 613 nsew power input
rlabel viali s 298661 140335 298695 140369 6 VPWR
port 613 nsew power input
rlabel viali s 1317 140335 1340 140369 6 VPWR
port 613 nsew power input
rlabel viali s 1225 140335 1259 140369 6 VPWR
port 613 nsew power input
rlabel viali s 1133 140335 1167 140369 6 VPWR
port 613 nsew power input
rlabel viali s 298753 141423 298787 141457 6 VPWR
port 613 nsew power input
rlabel viali s 298661 141423 298695 141457 6 VPWR
port 613 nsew power input
rlabel viali s 1317 141423 1340 141457 6 VPWR
port 613 nsew power input
rlabel viali s 1225 141423 1259 141457 6 VPWR
port 613 nsew power input
rlabel viali s 1133 141423 1167 141457 6 VPWR
port 613 nsew power input
rlabel viali s 298753 142511 298787 142545 6 VPWR
port 613 nsew power input
rlabel viali s 298661 142511 298695 142545 6 VPWR
port 613 nsew power input
rlabel viali s 1317 142511 1340 142545 6 VPWR
port 613 nsew power input
rlabel viali s 1225 142511 1259 142545 6 VPWR
port 613 nsew power input
rlabel viali s 1133 142511 1167 142545 6 VPWR
port 613 nsew power input
rlabel viali s 298753 143599 298787 143633 6 VPWR
port 613 nsew power input
rlabel viali s 298661 143599 298695 143633 6 VPWR
port 613 nsew power input
rlabel viali s 1317 143599 1340 143633 6 VPWR
port 613 nsew power input
rlabel viali s 1225 143599 1259 143633 6 VPWR
port 613 nsew power input
rlabel viali s 1133 143599 1167 143633 6 VPWR
port 613 nsew power input
rlabel viali s 298753 144687 298787 144721 6 VPWR
port 613 nsew power input
rlabel viali s 298661 144687 298695 144721 6 VPWR
port 613 nsew power input
rlabel viali s 1317 144687 1340 144721 6 VPWR
port 613 nsew power input
rlabel viali s 1225 144687 1259 144721 6 VPWR
port 613 nsew power input
rlabel viali s 1133 144687 1167 144721 6 VPWR
port 613 nsew power input
rlabel viali s 298753 145775 298787 145809 6 VPWR
port 613 nsew power input
rlabel viali s 298661 145775 298695 145809 6 VPWR
port 613 nsew power input
rlabel viali s 1317 145775 1340 145809 6 VPWR
port 613 nsew power input
rlabel viali s 1225 145775 1259 145809 6 VPWR
port 613 nsew power input
rlabel viali s 1133 145775 1167 145809 6 VPWR
port 613 nsew power input
rlabel viali s 298753 146863 298787 146897 6 VPWR
port 613 nsew power input
rlabel viali s 298661 146863 298695 146897 6 VPWR
port 613 nsew power input
rlabel viali s 1317 146863 1340 146897 6 VPWR
port 613 nsew power input
rlabel viali s 1225 146863 1259 146897 6 VPWR
port 613 nsew power input
rlabel viali s 1133 146863 1167 146897 6 VPWR
port 613 nsew power input
rlabel viali s 298753 147951 298787 147985 6 VPWR
port 613 nsew power input
rlabel viali s 298661 147951 298695 147985 6 VPWR
port 613 nsew power input
rlabel viali s 1317 147951 1340 147985 6 VPWR
port 613 nsew power input
rlabel viali s 1225 147951 1259 147985 6 VPWR
port 613 nsew power input
rlabel viali s 1133 147951 1167 147985 6 VPWR
port 613 nsew power input
rlabel viali s 298753 149039 298787 149073 6 VPWR
port 613 nsew power input
rlabel viali s 298661 149039 298695 149073 6 VPWR
port 613 nsew power input
rlabel viali s 1317 149039 1340 149073 6 VPWR
port 613 nsew power input
rlabel viali s 1225 149039 1259 149073 6 VPWR
port 613 nsew power input
rlabel viali s 1133 149039 1167 149073 6 VPWR
port 613 nsew power input
rlabel viali s 298753 150127 298787 150161 6 VPWR
port 613 nsew power input
rlabel viali s 298661 150127 298695 150161 6 VPWR
port 613 nsew power input
rlabel viali s 1317 150127 1340 150161 6 VPWR
port 613 nsew power input
rlabel viali s 1225 150127 1259 150161 6 VPWR
port 613 nsew power input
rlabel viali s 1133 150127 1167 150161 6 VPWR
port 613 nsew power input
rlabel viali s 298753 151215 298787 151249 6 VPWR
port 613 nsew power input
rlabel viali s 298661 151215 298695 151249 6 VPWR
port 613 nsew power input
rlabel viali s 1317 151215 1340 151249 6 VPWR
port 613 nsew power input
rlabel viali s 1225 151215 1259 151249 6 VPWR
port 613 nsew power input
rlabel viali s 1133 151215 1167 151249 6 VPWR
port 613 nsew power input
rlabel viali s 298753 152303 298787 152337 6 VPWR
port 613 nsew power input
rlabel viali s 298661 152303 298695 152337 6 VPWR
port 613 nsew power input
rlabel viali s 1317 152303 1340 152337 6 VPWR
port 613 nsew power input
rlabel viali s 1225 152303 1259 152337 6 VPWR
port 613 nsew power input
rlabel viali s 1133 152303 1167 152337 6 VPWR
port 613 nsew power input
rlabel viali s 298753 153391 298787 153425 6 VPWR
port 613 nsew power input
rlabel viali s 298661 153391 298695 153425 6 VPWR
port 613 nsew power input
rlabel viali s 1317 153391 1340 153425 6 VPWR
port 613 nsew power input
rlabel viali s 1225 153391 1259 153425 6 VPWR
port 613 nsew power input
rlabel viali s 1133 153391 1167 153425 6 VPWR
port 613 nsew power input
rlabel viali s 298753 154479 298787 154513 6 VPWR
port 613 nsew power input
rlabel viali s 298661 154479 298695 154513 6 VPWR
port 613 nsew power input
rlabel viali s 1317 154479 1340 154513 6 VPWR
port 613 nsew power input
rlabel viali s 1225 154479 1259 154513 6 VPWR
port 613 nsew power input
rlabel viali s 1133 154479 1167 154513 6 VPWR
port 613 nsew power input
rlabel viali s 298753 155567 298787 155601 6 VPWR
port 613 nsew power input
rlabel viali s 298661 155567 298695 155601 6 VPWR
port 613 nsew power input
rlabel viali s 1317 155567 1340 155601 6 VPWR
port 613 nsew power input
rlabel viali s 1225 155567 1259 155601 6 VPWR
port 613 nsew power input
rlabel viali s 1133 155567 1167 155601 6 VPWR
port 613 nsew power input
rlabel viali s 298753 156655 298787 156689 6 VPWR
port 613 nsew power input
rlabel viali s 298661 156655 298695 156689 6 VPWR
port 613 nsew power input
rlabel viali s 1317 156655 1340 156689 6 VPWR
port 613 nsew power input
rlabel viali s 1225 156655 1259 156689 6 VPWR
port 613 nsew power input
rlabel viali s 1133 156655 1167 156689 6 VPWR
port 613 nsew power input
rlabel viali s 298753 157743 298787 157777 6 VPWR
port 613 nsew power input
rlabel viali s 298661 157743 298695 157777 6 VPWR
port 613 nsew power input
rlabel viali s 1317 157743 1340 157777 6 VPWR
port 613 nsew power input
rlabel viali s 1225 157743 1259 157777 6 VPWR
port 613 nsew power input
rlabel viali s 1133 157743 1167 157777 6 VPWR
port 613 nsew power input
rlabel viali s 298753 158831 298787 158865 6 VPWR
port 613 nsew power input
rlabel viali s 298661 158831 298695 158865 6 VPWR
port 613 nsew power input
rlabel viali s 1317 158831 1340 158865 6 VPWR
port 613 nsew power input
rlabel viali s 1225 158831 1259 158865 6 VPWR
port 613 nsew power input
rlabel viali s 1133 158831 1167 158865 6 VPWR
port 613 nsew power input
rlabel viali s 298753 159919 298787 159953 6 VPWR
port 613 nsew power input
rlabel viali s 298661 159919 298695 159953 6 VPWR
port 613 nsew power input
rlabel viali s 1317 159919 1340 159953 6 VPWR
port 613 nsew power input
rlabel viali s 1225 159919 1259 159953 6 VPWR
port 613 nsew power input
rlabel viali s 1133 159919 1167 159953 6 VPWR
port 613 nsew power input
rlabel viali s 298753 161007 298787 161041 6 VPWR
port 613 nsew power input
rlabel viali s 298661 161007 298695 161041 6 VPWR
port 613 nsew power input
rlabel viali s 1317 161007 1340 161041 6 VPWR
port 613 nsew power input
rlabel viali s 1225 161007 1259 161041 6 VPWR
port 613 nsew power input
rlabel viali s 1133 161007 1167 161041 6 VPWR
port 613 nsew power input
rlabel viali s 298753 162095 298787 162129 6 VPWR
port 613 nsew power input
rlabel viali s 298661 162095 298695 162129 6 VPWR
port 613 nsew power input
rlabel viali s 1317 162095 1340 162129 6 VPWR
port 613 nsew power input
rlabel viali s 1225 162095 1259 162129 6 VPWR
port 613 nsew power input
rlabel viali s 1133 162095 1167 162129 6 VPWR
port 613 nsew power input
rlabel viali s 298753 163183 298787 163217 6 VPWR
port 613 nsew power input
rlabel viali s 298661 163183 298695 163217 6 VPWR
port 613 nsew power input
rlabel viali s 1317 163183 1340 163217 6 VPWR
port 613 nsew power input
rlabel viali s 1225 163183 1259 163217 6 VPWR
port 613 nsew power input
rlabel viali s 1133 163183 1167 163217 6 VPWR
port 613 nsew power input
rlabel viali s 298753 164271 298787 164305 6 VPWR
port 613 nsew power input
rlabel viali s 298661 164271 298695 164305 6 VPWR
port 613 nsew power input
rlabel viali s 1317 164271 1340 164305 6 VPWR
port 613 nsew power input
rlabel viali s 1225 164271 1259 164305 6 VPWR
port 613 nsew power input
rlabel viali s 1133 164271 1167 164305 6 VPWR
port 613 nsew power input
rlabel viali s 298753 165359 298787 165393 6 VPWR
port 613 nsew power input
rlabel viali s 298661 165359 298695 165393 6 VPWR
port 613 nsew power input
rlabel viali s 1317 165359 1340 165393 6 VPWR
port 613 nsew power input
rlabel viali s 1225 165359 1259 165393 6 VPWR
port 613 nsew power input
rlabel viali s 1133 165359 1167 165393 6 VPWR
port 613 nsew power input
rlabel viali s 298753 166447 298787 166481 6 VPWR
port 613 nsew power input
rlabel viali s 298661 166447 298695 166481 6 VPWR
port 613 nsew power input
rlabel viali s 1317 166447 1340 166481 6 VPWR
port 613 nsew power input
rlabel viali s 1225 166447 1259 166481 6 VPWR
port 613 nsew power input
rlabel viali s 1133 166447 1167 166481 6 VPWR
port 613 nsew power input
rlabel viali s 298753 167535 298787 167569 6 VPWR
port 613 nsew power input
rlabel viali s 298661 167535 298695 167569 6 VPWR
port 613 nsew power input
rlabel viali s 1317 167535 1340 167569 6 VPWR
port 613 nsew power input
rlabel viali s 1225 167535 1259 167569 6 VPWR
port 613 nsew power input
rlabel viali s 1133 167535 1167 167569 6 VPWR
port 613 nsew power input
rlabel viali s 298753 168623 298787 168657 6 VPWR
port 613 nsew power input
rlabel viali s 298661 168623 298695 168657 6 VPWR
port 613 nsew power input
rlabel viali s 1317 168623 1340 168657 6 VPWR
port 613 nsew power input
rlabel viali s 1225 168623 1259 168657 6 VPWR
port 613 nsew power input
rlabel viali s 1133 168623 1167 168657 6 VPWR
port 613 nsew power input
rlabel viali s 298753 169711 298787 169745 6 VPWR
port 613 nsew power input
rlabel viali s 298661 169711 298695 169745 6 VPWR
port 613 nsew power input
rlabel viali s 1317 169711 1340 169745 6 VPWR
port 613 nsew power input
rlabel viali s 1225 169711 1259 169745 6 VPWR
port 613 nsew power input
rlabel viali s 1133 169711 1167 169745 6 VPWR
port 613 nsew power input
rlabel viali s 298753 170799 298787 170833 6 VPWR
port 613 nsew power input
rlabel viali s 298661 170799 298695 170833 6 VPWR
port 613 nsew power input
rlabel viali s 1317 170799 1340 170833 6 VPWR
port 613 nsew power input
rlabel viali s 1225 170799 1259 170833 6 VPWR
port 613 nsew power input
rlabel viali s 1133 170799 1167 170833 6 VPWR
port 613 nsew power input
rlabel viali s 298753 171887 298787 171921 6 VPWR
port 613 nsew power input
rlabel viali s 298661 171887 298695 171921 6 VPWR
port 613 nsew power input
rlabel viali s 1317 171887 1340 171921 6 VPWR
port 613 nsew power input
rlabel viali s 1225 171887 1259 171921 6 VPWR
port 613 nsew power input
rlabel viali s 1133 171887 1167 171921 6 VPWR
port 613 nsew power input
rlabel viali s 298753 172975 298787 173009 6 VPWR
port 613 nsew power input
rlabel viali s 298661 172975 298695 173009 6 VPWR
port 613 nsew power input
rlabel viali s 1317 172975 1340 173009 6 VPWR
port 613 nsew power input
rlabel viali s 1225 172975 1259 173009 6 VPWR
port 613 nsew power input
rlabel viali s 1133 172975 1167 173009 6 VPWR
port 613 nsew power input
rlabel viali s 298753 174063 298787 174097 6 VPWR
port 613 nsew power input
rlabel viali s 298661 174063 298695 174097 6 VPWR
port 613 nsew power input
rlabel viali s 1317 174063 1340 174097 6 VPWR
port 613 nsew power input
rlabel viali s 1225 174063 1259 174097 6 VPWR
port 613 nsew power input
rlabel viali s 1133 174063 1167 174097 6 VPWR
port 613 nsew power input
rlabel viali s 298753 175151 298787 175185 6 VPWR
port 613 nsew power input
rlabel viali s 298661 175151 298695 175185 6 VPWR
port 613 nsew power input
rlabel viali s 1317 175151 1340 175185 6 VPWR
port 613 nsew power input
rlabel viali s 1225 175151 1259 175185 6 VPWR
port 613 nsew power input
rlabel viali s 1133 175151 1167 175185 6 VPWR
port 613 nsew power input
rlabel viali s 298753 176239 298787 176273 6 VPWR
port 613 nsew power input
rlabel viali s 298661 176239 298695 176273 6 VPWR
port 613 nsew power input
rlabel viali s 1317 176239 1340 176273 6 VPWR
port 613 nsew power input
rlabel viali s 1225 176239 1259 176273 6 VPWR
port 613 nsew power input
rlabel viali s 1133 176239 1167 176273 6 VPWR
port 613 nsew power input
rlabel viali s 298753 177327 298787 177361 6 VPWR
port 613 nsew power input
rlabel viali s 298661 177327 298695 177361 6 VPWR
port 613 nsew power input
rlabel viali s 1317 177327 1340 177361 6 VPWR
port 613 nsew power input
rlabel viali s 1225 177327 1259 177361 6 VPWR
port 613 nsew power input
rlabel viali s 1133 177327 1167 177361 6 VPWR
port 613 nsew power input
rlabel viali s 298753 178415 298787 178449 6 VPWR
port 613 nsew power input
rlabel viali s 298661 178415 298695 178449 6 VPWR
port 613 nsew power input
rlabel viali s 1317 178415 1340 178449 6 VPWR
port 613 nsew power input
rlabel viali s 1225 178415 1259 178449 6 VPWR
port 613 nsew power input
rlabel viali s 1133 178415 1167 178449 6 VPWR
port 613 nsew power input
rlabel viali s 298753 179503 298787 179537 6 VPWR
port 613 nsew power input
rlabel viali s 298661 179503 298695 179537 6 VPWR
port 613 nsew power input
rlabel viali s 1317 179503 1340 179537 6 VPWR
port 613 nsew power input
rlabel viali s 1225 179503 1259 179537 6 VPWR
port 613 nsew power input
rlabel viali s 1133 179503 1167 179537 6 VPWR
port 613 nsew power input
rlabel viali s 298753 180591 298787 180625 6 VPWR
port 613 nsew power input
rlabel viali s 298661 180591 298695 180625 6 VPWR
port 613 nsew power input
rlabel viali s 1317 180591 1340 180625 6 VPWR
port 613 nsew power input
rlabel viali s 1225 180591 1259 180625 6 VPWR
port 613 nsew power input
rlabel viali s 1133 180591 1167 180625 6 VPWR
port 613 nsew power input
rlabel viali s 298753 181679 298787 181713 6 VPWR
port 613 nsew power input
rlabel viali s 298661 181679 298695 181713 6 VPWR
port 613 nsew power input
rlabel viali s 1317 181679 1340 181713 6 VPWR
port 613 nsew power input
rlabel viali s 1225 181679 1259 181713 6 VPWR
port 613 nsew power input
rlabel viali s 1133 181679 1167 181713 6 VPWR
port 613 nsew power input
rlabel viali s 298753 182767 298787 182801 6 VPWR
port 613 nsew power input
rlabel viali s 298661 182767 298695 182801 6 VPWR
port 613 nsew power input
rlabel viali s 1317 182767 1340 182801 6 VPWR
port 613 nsew power input
rlabel viali s 1225 182767 1259 182801 6 VPWR
port 613 nsew power input
rlabel viali s 1133 182767 1167 182801 6 VPWR
port 613 nsew power input
rlabel viali s 298753 183855 298787 183889 6 VPWR
port 613 nsew power input
rlabel viali s 298661 183855 298695 183889 6 VPWR
port 613 nsew power input
rlabel viali s 1317 183855 1340 183889 6 VPWR
port 613 nsew power input
rlabel viali s 1225 183855 1259 183889 6 VPWR
port 613 nsew power input
rlabel viali s 1133 183855 1167 183889 6 VPWR
port 613 nsew power input
rlabel viali s 298753 184943 298787 184977 6 VPWR
port 613 nsew power input
rlabel viali s 298661 184943 298695 184977 6 VPWR
port 613 nsew power input
rlabel viali s 1317 184943 1340 184977 6 VPWR
port 613 nsew power input
rlabel viali s 1225 184943 1259 184977 6 VPWR
port 613 nsew power input
rlabel viali s 1133 184943 1167 184977 6 VPWR
port 613 nsew power input
rlabel viali s 298753 186031 298787 186065 6 VPWR
port 613 nsew power input
rlabel viali s 298661 186031 298695 186065 6 VPWR
port 613 nsew power input
rlabel viali s 1317 186031 1340 186065 6 VPWR
port 613 nsew power input
rlabel viali s 1225 186031 1259 186065 6 VPWR
port 613 nsew power input
rlabel viali s 1133 186031 1167 186065 6 VPWR
port 613 nsew power input
rlabel viali s 298753 187119 298787 187153 6 VPWR
port 613 nsew power input
rlabel viali s 298661 187119 298695 187153 6 VPWR
port 613 nsew power input
rlabel viali s 1317 187119 1340 187153 6 VPWR
port 613 nsew power input
rlabel viali s 1225 187119 1259 187153 6 VPWR
port 613 nsew power input
rlabel viali s 1133 187119 1167 187153 6 VPWR
port 613 nsew power input
rlabel viali s 298753 188207 298787 188241 6 VPWR
port 613 nsew power input
rlabel viali s 298661 188207 298695 188241 6 VPWR
port 613 nsew power input
rlabel viali s 1317 188207 1340 188241 6 VPWR
port 613 nsew power input
rlabel viali s 1225 188207 1259 188241 6 VPWR
port 613 nsew power input
rlabel viali s 1133 188207 1167 188241 6 VPWR
port 613 nsew power input
rlabel viali s 298753 189295 298787 189329 6 VPWR
port 613 nsew power input
rlabel viali s 298661 189295 298695 189329 6 VPWR
port 613 nsew power input
rlabel viali s 1317 189295 1340 189329 6 VPWR
port 613 nsew power input
rlabel viali s 1225 189295 1259 189329 6 VPWR
port 613 nsew power input
rlabel viali s 1133 189295 1167 189329 6 VPWR
port 613 nsew power input
rlabel viali s 298753 190383 298787 190417 6 VPWR
port 613 nsew power input
rlabel viali s 298661 190383 298695 190417 6 VPWR
port 613 nsew power input
rlabel viali s 1317 190383 1340 190417 6 VPWR
port 613 nsew power input
rlabel viali s 1225 190383 1259 190417 6 VPWR
port 613 nsew power input
rlabel viali s 1133 190383 1167 190417 6 VPWR
port 613 nsew power input
rlabel viali s 298753 191471 298787 191505 6 VPWR
port 613 nsew power input
rlabel viali s 298661 191471 298695 191505 6 VPWR
port 613 nsew power input
rlabel viali s 1317 191471 1340 191505 6 VPWR
port 613 nsew power input
rlabel viali s 1225 191471 1259 191505 6 VPWR
port 613 nsew power input
rlabel viali s 1133 191471 1167 191505 6 VPWR
port 613 nsew power input
rlabel viali s 298753 192559 298787 192593 6 VPWR
port 613 nsew power input
rlabel viali s 298661 192559 298695 192593 6 VPWR
port 613 nsew power input
rlabel viali s 1317 192559 1340 192593 6 VPWR
port 613 nsew power input
rlabel viali s 1225 192559 1259 192593 6 VPWR
port 613 nsew power input
rlabel viali s 1133 192559 1167 192593 6 VPWR
port 613 nsew power input
rlabel viali s 298753 193647 298787 193681 6 VPWR
port 613 nsew power input
rlabel viali s 298661 193647 298695 193681 6 VPWR
port 613 nsew power input
rlabel viali s 1317 193647 1340 193681 6 VPWR
port 613 nsew power input
rlabel viali s 1225 193647 1259 193681 6 VPWR
port 613 nsew power input
rlabel viali s 1133 193647 1167 193681 6 VPWR
port 613 nsew power input
rlabel viali s 298753 194735 298787 194769 6 VPWR
port 613 nsew power input
rlabel viali s 298661 194735 298695 194769 6 VPWR
port 613 nsew power input
rlabel viali s 1317 194735 1340 194769 6 VPWR
port 613 nsew power input
rlabel viali s 1225 194735 1259 194769 6 VPWR
port 613 nsew power input
rlabel viali s 1133 194735 1167 194769 6 VPWR
port 613 nsew power input
rlabel viali s 298753 195823 298787 195857 6 VPWR
port 613 nsew power input
rlabel viali s 298661 195823 298695 195857 6 VPWR
port 613 nsew power input
rlabel viali s 1317 195823 1340 195857 6 VPWR
port 613 nsew power input
rlabel viali s 1225 195823 1259 195857 6 VPWR
port 613 nsew power input
rlabel viali s 1133 195823 1167 195857 6 VPWR
port 613 nsew power input
rlabel viali s 298753 196911 298787 196945 6 VPWR
port 613 nsew power input
rlabel viali s 298661 196911 298695 196945 6 VPWR
port 613 nsew power input
rlabel viali s 1317 196911 1340 196945 6 VPWR
port 613 nsew power input
rlabel viali s 1225 196911 1259 196945 6 VPWR
port 613 nsew power input
rlabel viali s 1133 196911 1167 196945 6 VPWR
port 613 nsew power input
rlabel viali s 298753 197999 298787 198033 6 VPWR
port 613 nsew power input
rlabel viali s 298661 197999 298695 198033 6 VPWR
port 613 nsew power input
rlabel viali s 1317 197999 1340 198033 6 VPWR
port 613 nsew power input
rlabel viali s 1225 197999 1259 198033 6 VPWR
port 613 nsew power input
rlabel viali s 1133 197999 1167 198033 6 VPWR
port 613 nsew power input
rlabel viali s 298753 199087 298787 199121 6 VPWR
port 613 nsew power input
rlabel viali s 298661 199087 298695 199121 6 VPWR
port 613 nsew power input
rlabel viali s 1317 199087 1340 199121 6 VPWR
port 613 nsew power input
rlabel viali s 1225 199087 1259 199121 6 VPWR
port 613 nsew power input
rlabel viali s 1133 199087 1167 199121 6 VPWR
port 613 nsew power input
rlabel viali s 298753 200175 298787 200209 6 VPWR
port 613 nsew power input
rlabel viali s 298661 200175 298695 200209 6 VPWR
port 613 nsew power input
rlabel viali s 1317 200175 1340 200209 6 VPWR
port 613 nsew power input
rlabel viali s 1225 200175 1259 200209 6 VPWR
port 613 nsew power input
rlabel viali s 1133 200175 1167 200209 6 VPWR
port 613 nsew power input
rlabel viali s 298753 201263 298787 201297 6 VPWR
port 613 nsew power input
rlabel viali s 298661 201263 298695 201297 6 VPWR
port 613 nsew power input
rlabel viali s 1317 201263 1340 201297 6 VPWR
port 613 nsew power input
rlabel viali s 1225 201263 1259 201297 6 VPWR
port 613 nsew power input
rlabel viali s 1133 201263 1167 201297 6 VPWR
port 613 nsew power input
rlabel viali s 298753 202351 298787 202385 6 VPWR
port 613 nsew power input
rlabel viali s 298661 202351 298695 202385 6 VPWR
port 613 nsew power input
rlabel viali s 1317 202351 1340 202385 6 VPWR
port 613 nsew power input
rlabel viali s 1225 202351 1259 202385 6 VPWR
port 613 nsew power input
rlabel viali s 1133 202351 1167 202385 6 VPWR
port 613 nsew power input
rlabel viali s 298753 203439 298787 203473 6 VPWR
port 613 nsew power input
rlabel viali s 298661 203439 298695 203473 6 VPWR
port 613 nsew power input
rlabel viali s 1317 203439 1340 203473 6 VPWR
port 613 nsew power input
rlabel viali s 1225 203439 1259 203473 6 VPWR
port 613 nsew power input
rlabel viali s 1133 203439 1167 203473 6 VPWR
port 613 nsew power input
rlabel viali s 298753 204527 298787 204561 6 VPWR
port 613 nsew power input
rlabel viali s 298661 204527 298695 204561 6 VPWR
port 613 nsew power input
rlabel viali s 1317 204527 1340 204561 6 VPWR
port 613 nsew power input
rlabel viali s 1225 204527 1259 204561 6 VPWR
port 613 nsew power input
rlabel viali s 1133 204527 1167 204561 6 VPWR
port 613 nsew power input
rlabel viali s 298753 205615 298787 205649 6 VPWR
port 613 nsew power input
rlabel viali s 298661 205615 298695 205649 6 VPWR
port 613 nsew power input
rlabel viali s 1317 205615 1340 205649 6 VPWR
port 613 nsew power input
rlabel viali s 1225 205615 1259 205649 6 VPWR
port 613 nsew power input
rlabel viali s 1133 205615 1167 205649 6 VPWR
port 613 nsew power input
rlabel viali s 298753 206703 298787 206737 6 VPWR
port 613 nsew power input
rlabel viali s 298661 206703 298695 206737 6 VPWR
port 613 nsew power input
rlabel viali s 1317 206703 1340 206737 6 VPWR
port 613 nsew power input
rlabel viali s 1225 206703 1259 206737 6 VPWR
port 613 nsew power input
rlabel viali s 1133 206703 1167 206737 6 VPWR
port 613 nsew power input
rlabel viali s 298753 207791 298787 207825 6 VPWR
port 613 nsew power input
rlabel viali s 298661 207791 298695 207825 6 VPWR
port 613 nsew power input
rlabel viali s 1317 207791 1340 207825 6 VPWR
port 613 nsew power input
rlabel viali s 1225 207791 1259 207825 6 VPWR
port 613 nsew power input
rlabel viali s 1133 207791 1167 207825 6 VPWR
port 613 nsew power input
rlabel viali s 298753 208879 298787 208913 6 VPWR
port 613 nsew power input
rlabel viali s 298661 208879 298695 208913 6 VPWR
port 613 nsew power input
rlabel viali s 1317 208879 1340 208913 6 VPWR
port 613 nsew power input
rlabel viali s 1225 208879 1259 208913 6 VPWR
port 613 nsew power input
rlabel viali s 1133 208879 1167 208913 6 VPWR
port 613 nsew power input
rlabel viali s 298753 209967 298787 210001 6 VPWR
port 613 nsew power input
rlabel viali s 298661 209967 298695 210001 6 VPWR
port 613 nsew power input
rlabel viali s 1317 209967 1340 210001 6 VPWR
port 613 nsew power input
rlabel viali s 1225 209967 1259 210001 6 VPWR
port 613 nsew power input
rlabel viali s 1133 209967 1167 210001 6 VPWR
port 613 nsew power input
rlabel viali s 298753 211055 298787 211089 6 VPWR
port 613 nsew power input
rlabel viali s 298661 211055 298695 211089 6 VPWR
port 613 nsew power input
rlabel viali s 1317 211055 1340 211089 6 VPWR
port 613 nsew power input
rlabel viali s 1225 211055 1259 211089 6 VPWR
port 613 nsew power input
rlabel viali s 1133 211055 1167 211089 6 VPWR
port 613 nsew power input
rlabel viali s 298753 212143 298787 212177 6 VPWR
port 613 nsew power input
rlabel viali s 298661 212143 298695 212177 6 VPWR
port 613 nsew power input
rlabel viali s 1317 212143 1340 212177 6 VPWR
port 613 nsew power input
rlabel viali s 1225 212143 1259 212177 6 VPWR
port 613 nsew power input
rlabel viali s 1133 212143 1167 212177 6 VPWR
port 613 nsew power input
rlabel viali s 298753 213231 298787 213265 6 VPWR
port 613 nsew power input
rlabel viali s 298661 213231 298695 213265 6 VPWR
port 613 nsew power input
rlabel viali s 1317 213231 1340 213265 6 VPWR
port 613 nsew power input
rlabel viali s 1225 213231 1259 213265 6 VPWR
port 613 nsew power input
rlabel viali s 1133 213231 1167 213265 6 VPWR
port 613 nsew power input
rlabel viali s 298753 214319 298787 214353 6 VPWR
port 613 nsew power input
rlabel viali s 298661 214319 298695 214353 6 VPWR
port 613 nsew power input
rlabel viali s 1317 214319 1340 214353 6 VPWR
port 613 nsew power input
rlabel viali s 1225 214319 1259 214353 6 VPWR
port 613 nsew power input
rlabel viali s 1133 214319 1167 214353 6 VPWR
port 613 nsew power input
rlabel viali s 298753 215407 298787 215441 6 VPWR
port 613 nsew power input
rlabel viali s 298661 215407 298695 215441 6 VPWR
port 613 nsew power input
rlabel viali s 1317 215407 1340 215441 6 VPWR
port 613 nsew power input
rlabel viali s 1225 215407 1259 215441 6 VPWR
port 613 nsew power input
rlabel viali s 1133 215407 1167 215441 6 VPWR
port 613 nsew power input
rlabel viali s 298753 216495 298787 216529 6 VPWR
port 613 nsew power input
rlabel viali s 298661 216495 298695 216529 6 VPWR
port 613 nsew power input
rlabel viali s 1317 216495 1340 216529 6 VPWR
port 613 nsew power input
rlabel viali s 1225 216495 1259 216529 6 VPWR
port 613 nsew power input
rlabel viali s 1133 216495 1167 216529 6 VPWR
port 613 nsew power input
rlabel viali s 298753 217583 298787 217617 6 VPWR
port 613 nsew power input
rlabel viali s 298661 217583 298695 217617 6 VPWR
port 613 nsew power input
rlabel viali s 1317 217583 1340 217617 6 VPWR
port 613 nsew power input
rlabel viali s 1225 217583 1259 217617 6 VPWR
port 613 nsew power input
rlabel viali s 1133 217583 1167 217617 6 VPWR
port 613 nsew power input
rlabel viali s 298753 218671 298787 218705 6 VPWR
port 613 nsew power input
rlabel viali s 298661 218671 298695 218705 6 VPWR
port 613 nsew power input
rlabel viali s 1317 218671 1340 218705 6 VPWR
port 613 nsew power input
rlabel viali s 1225 218671 1259 218705 6 VPWR
port 613 nsew power input
rlabel viali s 1133 218671 1167 218705 6 VPWR
port 613 nsew power input
rlabel viali s 298753 219759 298787 219793 6 VPWR
port 613 nsew power input
rlabel viali s 298661 219759 298695 219793 6 VPWR
port 613 nsew power input
rlabel viali s 1317 219759 1340 219793 6 VPWR
port 613 nsew power input
rlabel viali s 1225 219759 1259 219793 6 VPWR
port 613 nsew power input
rlabel viali s 1133 219759 1167 219793 6 VPWR
port 613 nsew power input
rlabel viali s 298753 220847 298787 220881 6 VPWR
port 613 nsew power input
rlabel viali s 298661 220847 298695 220881 6 VPWR
port 613 nsew power input
rlabel viali s 1317 220847 1340 220881 6 VPWR
port 613 nsew power input
rlabel viali s 1225 220847 1259 220881 6 VPWR
port 613 nsew power input
rlabel viali s 1133 220847 1167 220881 6 VPWR
port 613 nsew power input
rlabel viali s 298753 221935 298787 221969 6 VPWR
port 613 nsew power input
rlabel viali s 298661 221935 298695 221969 6 VPWR
port 613 nsew power input
rlabel viali s 1317 221935 1340 221969 6 VPWR
port 613 nsew power input
rlabel viali s 1225 221935 1259 221969 6 VPWR
port 613 nsew power input
rlabel viali s 1133 221935 1167 221969 6 VPWR
port 613 nsew power input
rlabel viali s 298753 223023 298787 223057 6 VPWR
port 613 nsew power input
rlabel viali s 298661 223023 298695 223057 6 VPWR
port 613 nsew power input
rlabel viali s 1317 223023 1340 223057 6 VPWR
port 613 nsew power input
rlabel viali s 1225 223023 1259 223057 6 VPWR
port 613 nsew power input
rlabel viali s 1133 223023 1167 223057 6 VPWR
port 613 nsew power input
rlabel viali s 298753 224111 298787 224145 6 VPWR
port 613 nsew power input
rlabel viali s 298661 224111 298695 224145 6 VPWR
port 613 nsew power input
rlabel viali s 1317 224111 1340 224145 6 VPWR
port 613 nsew power input
rlabel viali s 1225 224111 1259 224145 6 VPWR
port 613 nsew power input
rlabel viali s 1133 224111 1167 224145 6 VPWR
port 613 nsew power input
rlabel viali s 298753 225199 298787 225233 6 VPWR
port 613 nsew power input
rlabel viali s 298661 225199 298695 225233 6 VPWR
port 613 nsew power input
rlabel viali s 1317 225199 1340 225233 6 VPWR
port 613 nsew power input
rlabel viali s 1225 225199 1259 225233 6 VPWR
port 613 nsew power input
rlabel viali s 1133 225199 1167 225233 6 VPWR
port 613 nsew power input
rlabel viali s 298753 226287 298787 226321 6 VPWR
port 613 nsew power input
rlabel viali s 298661 226287 298695 226321 6 VPWR
port 613 nsew power input
rlabel viali s 1317 226287 1340 226321 6 VPWR
port 613 nsew power input
rlabel viali s 1225 226287 1259 226321 6 VPWR
port 613 nsew power input
rlabel viali s 1133 226287 1167 226321 6 VPWR
port 613 nsew power input
rlabel viali s 298753 227375 298787 227409 6 VPWR
port 613 nsew power input
rlabel viali s 298661 227375 298695 227409 6 VPWR
port 613 nsew power input
rlabel viali s 1317 227375 1340 227409 6 VPWR
port 613 nsew power input
rlabel viali s 1225 227375 1259 227409 6 VPWR
port 613 nsew power input
rlabel viali s 1133 227375 1167 227409 6 VPWR
port 613 nsew power input
rlabel viali s 298753 228463 298787 228497 6 VPWR
port 613 nsew power input
rlabel viali s 298661 228463 298695 228497 6 VPWR
port 613 nsew power input
rlabel viali s 1317 228463 1340 228497 6 VPWR
port 613 nsew power input
rlabel viali s 1225 228463 1259 228497 6 VPWR
port 613 nsew power input
rlabel viali s 1133 228463 1167 228497 6 VPWR
port 613 nsew power input
rlabel viali s 298753 229551 298787 229585 6 VPWR
port 613 nsew power input
rlabel viali s 298661 229551 298695 229585 6 VPWR
port 613 nsew power input
rlabel viali s 1317 229551 1340 229585 6 VPWR
port 613 nsew power input
rlabel viali s 1225 229551 1259 229585 6 VPWR
port 613 nsew power input
rlabel viali s 1133 229551 1167 229585 6 VPWR
port 613 nsew power input
rlabel viali s 298753 230639 298787 230673 6 VPWR
port 613 nsew power input
rlabel viali s 298661 230639 298695 230673 6 VPWR
port 613 nsew power input
rlabel viali s 1317 230639 1340 230673 6 VPWR
port 613 nsew power input
rlabel viali s 1225 230639 1259 230673 6 VPWR
port 613 nsew power input
rlabel viali s 1133 230639 1167 230673 6 VPWR
port 613 nsew power input
rlabel viali s 298753 231727 298787 231761 6 VPWR
port 613 nsew power input
rlabel viali s 298661 231727 298695 231761 6 VPWR
port 613 nsew power input
rlabel viali s 1317 231727 1340 231761 6 VPWR
port 613 nsew power input
rlabel viali s 1225 231727 1259 231761 6 VPWR
port 613 nsew power input
rlabel viali s 1133 231727 1167 231761 6 VPWR
port 613 nsew power input
rlabel viali s 298753 232815 298787 232849 6 VPWR
port 613 nsew power input
rlabel viali s 298661 232815 298695 232849 6 VPWR
port 613 nsew power input
rlabel viali s 1317 232815 1340 232849 6 VPWR
port 613 nsew power input
rlabel viali s 1225 232815 1259 232849 6 VPWR
port 613 nsew power input
rlabel viali s 1133 232815 1167 232849 6 VPWR
port 613 nsew power input
rlabel viali s 298753 233903 298787 233937 6 VPWR
port 613 nsew power input
rlabel viali s 298661 233903 298695 233937 6 VPWR
port 613 nsew power input
rlabel viali s 1317 233903 1340 233937 6 VPWR
port 613 nsew power input
rlabel viali s 1225 233903 1259 233937 6 VPWR
port 613 nsew power input
rlabel viali s 1133 233903 1167 233937 6 VPWR
port 613 nsew power input
rlabel viali s 298753 234991 298787 235025 6 VPWR
port 613 nsew power input
rlabel viali s 298661 234991 298695 235025 6 VPWR
port 613 nsew power input
rlabel viali s 1317 234991 1340 235025 6 VPWR
port 613 nsew power input
rlabel viali s 1225 234991 1259 235025 6 VPWR
port 613 nsew power input
rlabel viali s 1133 234991 1167 235025 6 VPWR
port 613 nsew power input
rlabel viali s 298753 236079 298787 236113 6 VPWR
port 613 nsew power input
rlabel viali s 298661 236079 298695 236113 6 VPWR
port 613 nsew power input
rlabel viali s 1317 236079 1340 236113 6 VPWR
port 613 nsew power input
rlabel viali s 1225 236079 1259 236113 6 VPWR
port 613 nsew power input
rlabel viali s 1133 236079 1167 236113 6 VPWR
port 613 nsew power input
rlabel viali s 298753 237167 298787 237201 6 VPWR
port 613 nsew power input
rlabel viali s 298661 237167 298695 237201 6 VPWR
port 613 nsew power input
rlabel viali s 1317 237167 1340 237201 6 VPWR
port 613 nsew power input
rlabel viali s 1225 237167 1259 237201 6 VPWR
port 613 nsew power input
rlabel viali s 1133 237167 1167 237201 6 VPWR
port 613 nsew power input
rlabel viali s 298753 238255 298787 238289 6 VPWR
port 613 nsew power input
rlabel viali s 298661 238255 298695 238289 6 VPWR
port 613 nsew power input
rlabel viali s 1317 238255 1340 238289 6 VPWR
port 613 nsew power input
rlabel viali s 1225 238255 1259 238289 6 VPWR
port 613 nsew power input
rlabel viali s 1133 238255 1167 238289 6 VPWR
port 613 nsew power input
rlabel viali s 298753 239343 298787 239377 6 VPWR
port 613 nsew power input
rlabel viali s 298661 239343 298695 239377 6 VPWR
port 613 nsew power input
rlabel viali s 1317 239343 1340 239377 6 VPWR
port 613 nsew power input
rlabel viali s 1225 239343 1259 239377 6 VPWR
port 613 nsew power input
rlabel viali s 1133 239343 1167 239377 6 VPWR
port 613 nsew power input
rlabel viali s 298753 240431 298787 240465 6 VPWR
port 613 nsew power input
rlabel viali s 298661 240431 298695 240465 6 VPWR
port 613 nsew power input
rlabel viali s 1317 240431 1340 240465 6 VPWR
port 613 nsew power input
rlabel viali s 1225 240431 1259 240465 6 VPWR
port 613 nsew power input
rlabel viali s 1133 240431 1167 240465 6 VPWR
port 613 nsew power input
rlabel viali s 298753 241519 298787 241553 6 VPWR
port 613 nsew power input
rlabel viali s 298661 241519 298695 241553 6 VPWR
port 613 nsew power input
rlabel viali s 1317 241519 1340 241553 6 VPWR
port 613 nsew power input
rlabel viali s 1225 241519 1259 241553 6 VPWR
port 613 nsew power input
rlabel viali s 1133 241519 1167 241553 6 VPWR
port 613 nsew power input
rlabel viali s 298753 242607 298787 242641 6 VPWR
port 613 nsew power input
rlabel viali s 298661 242607 298695 242641 6 VPWR
port 613 nsew power input
rlabel viali s 1317 242607 1340 242641 6 VPWR
port 613 nsew power input
rlabel viali s 1225 242607 1259 242641 6 VPWR
port 613 nsew power input
rlabel viali s 1133 242607 1167 242641 6 VPWR
port 613 nsew power input
rlabel viali s 298753 243695 298787 243729 6 VPWR
port 613 nsew power input
rlabel viali s 298661 243695 298695 243729 6 VPWR
port 613 nsew power input
rlabel viali s 1317 243695 1340 243729 6 VPWR
port 613 nsew power input
rlabel viali s 1225 243695 1259 243729 6 VPWR
port 613 nsew power input
rlabel viali s 1133 243695 1167 243729 6 VPWR
port 613 nsew power input
rlabel viali s 298753 244783 298787 244817 6 VPWR
port 613 nsew power input
rlabel viali s 298661 244783 298695 244817 6 VPWR
port 613 nsew power input
rlabel viali s 1317 244783 1340 244817 6 VPWR
port 613 nsew power input
rlabel viali s 1225 244783 1259 244817 6 VPWR
port 613 nsew power input
rlabel viali s 1133 244783 1167 244817 6 VPWR
port 613 nsew power input
rlabel viali s 298753 245871 298787 245905 6 VPWR
port 613 nsew power input
rlabel viali s 298661 245871 298695 245905 6 VPWR
port 613 nsew power input
rlabel viali s 1317 245871 1340 245905 6 VPWR
port 613 nsew power input
rlabel viali s 1225 245871 1259 245905 6 VPWR
port 613 nsew power input
rlabel viali s 1133 245871 1167 245905 6 VPWR
port 613 nsew power input
rlabel viali s 298753 246959 298787 246993 6 VPWR
port 613 nsew power input
rlabel viali s 298661 246959 298695 246993 6 VPWR
port 613 nsew power input
rlabel viali s 1317 246959 1340 246993 6 VPWR
port 613 nsew power input
rlabel viali s 1225 246959 1259 246993 6 VPWR
port 613 nsew power input
rlabel viali s 1133 246959 1167 246993 6 VPWR
port 613 nsew power input
rlabel viali s 298753 248047 298787 248081 6 VPWR
port 613 nsew power input
rlabel viali s 298661 248047 298695 248081 6 VPWR
port 613 nsew power input
rlabel viali s 1317 248047 1340 248081 6 VPWR
port 613 nsew power input
rlabel viali s 1225 248047 1259 248081 6 VPWR
port 613 nsew power input
rlabel viali s 1133 248047 1167 248081 6 VPWR
port 613 nsew power input
rlabel viali s 298753 249135 298787 249169 6 VPWR
port 613 nsew power input
rlabel viali s 298661 249135 298695 249169 6 VPWR
port 613 nsew power input
rlabel viali s 1317 249135 1340 249169 6 VPWR
port 613 nsew power input
rlabel viali s 1225 249135 1259 249169 6 VPWR
port 613 nsew power input
rlabel viali s 1133 249135 1167 249169 6 VPWR
port 613 nsew power input
rlabel viali s 298753 250223 298787 250257 6 VPWR
port 613 nsew power input
rlabel viali s 298661 250223 298695 250257 6 VPWR
port 613 nsew power input
rlabel viali s 1317 250223 1340 250257 6 VPWR
port 613 nsew power input
rlabel viali s 1225 250223 1259 250257 6 VPWR
port 613 nsew power input
rlabel viali s 1133 250223 1167 250257 6 VPWR
port 613 nsew power input
rlabel viali s 298753 251311 298787 251345 6 VPWR
port 613 nsew power input
rlabel viali s 298661 251311 298695 251345 6 VPWR
port 613 nsew power input
rlabel viali s 1317 251311 1340 251345 6 VPWR
port 613 nsew power input
rlabel viali s 1225 251311 1259 251345 6 VPWR
port 613 nsew power input
rlabel viali s 1133 251311 1167 251345 6 VPWR
port 613 nsew power input
rlabel viali s 298753 252399 298787 252433 6 VPWR
port 613 nsew power input
rlabel viali s 298661 252399 298695 252433 6 VPWR
port 613 nsew power input
rlabel viali s 1317 252399 1340 252433 6 VPWR
port 613 nsew power input
rlabel viali s 1225 252399 1259 252433 6 VPWR
port 613 nsew power input
rlabel viali s 1133 252399 1167 252433 6 VPWR
port 613 nsew power input
rlabel viali s 298753 253487 298787 253521 6 VPWR
port 613 nsew power input
rlabel viali s 298661 253487 298695 253521 6 VPWR
port 613 nsew power input
rlabel viali s 1317 253487 1340 253521 6 VPWR
port 613 nsew power input
rlabel viali s 1225 253487 1259 253521 6 VPWR
port 613 nsew power input
rlabel viali s 1133 253487 1167 253521 6 VPWR
port 613 nsew power input
rlabel viali s 298753 254575 298787 254609 6 VPWR
port 613 nsew power input
rlabel viali s 298661 254575 298695 254609 6 VPWR
port 613 nsew power input
rlabel viali s 1317 254575 1340 254609 6 VPWR
port 613 nsew power input
rlabel viali s 1225 254575 1259 254609 6 VPWR
port 613 nsew power input
rlabel viali s 1133 254575 1167 254609 6 VPWR
port 613 nsew power input
rlabel viali s 298753 255663 298787 255697 6 VPWR
port 613 nsew power input
rlabel viali s 298661 255663 298695 255697 6 VPWR
port 613 nsew power input
rlabel viali s 1317 255663 1340 255697 6 VPWR
port 613 nsew power input
rlabel viali s 1225 255663 1259 255697 6 VPWR
port 613 nsew power input
rlabel viali s 1133 255663 1167 255697 6 VPWR
port 613 nsew power input
rlabel viali s 298753 256751 298787 256785 6 VPWR
port 613 nsew power input
rlabel viali s 298661 256751 298695 256785 6 VPWR
port 613 nsew power input
rlabel viali s 1317 256751 1340 256785 6 VPWR
port 613 nsew power input
rlabel viali s 1225 256751 1259 256785 6 VPWR
port 613 nsew power input
rlabel viali s 1133 256751 1167 256785 6 VPWR
port 613 nsew power input
rlabel viali s 298753 257839 298787 257873 6 VPWR
port 613 nsew power input
rlabel viali s 298661 257839 298695 257873 6 VPWR
port 613 nsew power input
rlabel viali s 1317 257839 1340 257873 6 VPWR
port 613 nsew power input
rlabel viali s 1225 257839 1259 257873 6 VPWR
port 613 nsew power input
rlabel viali s 1133 257839 1167 257873 6 VPWR
port 613 nsew power input
rlabel viali s 298753 258927 298787 258961 6 VPWR
port 613 nsew power input
rlabel viali s 298661 258927 298695 258961 6 VPWR
port 613 nsew power input
rlabel viali s 1317 258927 1340 258961 6 VPWR
port 613 nsew power input
rlabel viali s 1225 258927 1259 258961 6 VPWR
port 613 nsew power input
rlabel viali s 1133 258927 1167 258961 6 VPWR
port 613 nsew power input
rlabel viali s 298753 260015 298787 260049 6 VPWR
port 613 nsew power input
rlabel viali s 298661 260015 298695 260049 6 VPWR
port 613 nsew power input
rlabel viali s 1317 260015 1340 260049 6 VPWR
port 613 nsew power input
rlabel viali s 1225 260015 1259 260049 6 VPWR
port 613 nsew power input
rlabel viali s 1133 260015 1167 260049 6 VPWR
port 613 nsew power input
rlabel viali s 298753 261103 298787 261137 6 VPWR
port 613 nsew power input
rlabel viali s 298661 261103 298695 261137 6 VPWR
port 613 nsew power input
rlabel viali s 1317 261103 1340 261137 6 VPWR
port 613 nsew power input
rlabel viali s 1225 261103 1259 261137 6 VPWR
port 613 nsew power input
rlabel viali s 1133 261103 1167 261137 6 VPWR
port 613 nsew power input
rlabel viali s 298753 262191 298787 262225 6 VPWR
port 613 nsew power input
rlabel viali s 298661 262191 298695 262225 6 VPWR
port 613 nsew power input
rlabel viali s 1317 262191 1340 262225 6 VPWR
port 613 nsew power input
rlabel viali s 1225 262191 1259 262225 6 VPWR
port 613 nsew power input
rlabel viali s 1133 262191 1167 262225 6 VPWR
port 613 nsew power input
rlabel viali s 298753 263279 298787 263313 6 VPWR
port 613 nsew power input
rlabel viali s 298661 263279 298695 263313 6 VPWR
port 613 nsew power input
rlabel viali s 1317 263279 1340 263313 6 VPWR
port 613 nsew power input
rlabel viali s 1225 263279 1259 263313 6 VPWR
port 613 nsew power input
rlabel viali s 1133 263279 1167 263313 6 VPWR
port 613 nsew power input
rlabel viali s 298753 264367 298787 264401 6 VPWR
port 613 nsew power input
rlabel viali s 298661 264367 298695 264401 6 VPWR
port 613 nsew power input
rlabel viali s 1317 264367 1340 264401 6 VPWR
port 613 nsew power input
rlabel viali s 1225 264367 1259 264401 6 VPWR
port 613 nsew power input
rlabel viali s 1133 264367 1167 264401 6 VPWR
port 613 nsew power input
rlabel viali s 298753 265455 298787 265489 6 VPWR
port 613 nsew power input
rlabel viali s 298661 265455 298695 265489 6 VPWR
port 613 nsew power input
rlabel viali s 1317 265455 1340 265489 6 VPWR
port 613 nsew power input
rlabel viali s 1225 265455 1259 265489 6 VPWR
port 613 nsew power input
rlabel viali s 1133 265455 1167 265489 6 VPWR
port 613 nsew power input
rlabel viali s 298753 266543 298787 266577 6 VPWR
port 613 nsew power input
rlabel viali s 298661 266543 298695 266577 6 VPWR
port 613 nsew power input
rlabel viali s 1317 266543 1340 266577 6 VPWR
port 613 nsew power input
rlabel viali s 1225 266543 1259 266577 6 VPWR
port 613 nsew power input
rlabel viali s 1133 266543 1167 266577 6 VPWR
port 613 nsew power input
rlabel viali s 298753 267631 298787 267665 6 VPWR
port 613 nsew power input
rlabel viali s 298661 267631 298695 267665 6 VPWR
port 613 nsew power input
rlabel viali s 1317 267631 1340 267665 6 VPWR
port 613 nsew power input
rlabel viali s 1225 267631 1259 267665 6 VPWR
port 613 nsew power input
rlabel viali s 1133 267631 1167 267665 6 VPWR
port 613 nsew power input
rlabel viali s 298753 268719 298787 268753 6 VPWR
port 613 nsew power input
rlabel viali s 298661 268719 298695 268753 6 VPWR
port 613 nsew power input
rlabel viali s 1317 268719 1340 268753 6 VPWR
port 613 nsew power input
rlabel viali s 1225 268719 1259 268753 6 VPWR
port 613 nsew power input
rlabel viali s 1133 268719 1167 268753 6 VPWR
port 613 nsew power input
rlabel viali s 298753 269807 298787 269841 6 VPWR
port 613 nsew power input
rlabel viali s 298661 269807 298695 269841 6 VPWR
port 613 nsew power input
rlabel viali s 1317 269807 1340 269841 6 VPWR
port 613 nsew power input
rlabel viali s 1225 269807 1259 269841 6 VPWR
port 613 nsew power input
rlabel viali s 1133 269807 1167 269841 6 VPWR
port 613 nsew power input
rlabel viali s 298753 270895 298787 270929 6 VPWR
port 613 nsew power input
rlabel viali s 298661 270895 298695 270929 6 VPWR
port 613 nsew power input
rlabel viali s 1317 270895 1340 270929 6 VPWR
port 613 nsew power input
rlabel viali s 1225 270895 1259 270929 6 VPWR
port 613 nsew power input
rlabel viali s 1133 270895 1167 270929 6 VPWR
port 613 nsew power input
rlabel viali s 298753 271983 298787 272017 6 VPWR
port 613 nsew power input
rlabel viali s 298661 271983 298695 272017 6 VPWR
port 613 nsew power input
rlabel viali s 1317 271983 1340 272017 6 VPWR
port 613 nsew power input
rlabel viali s 1225 271983 1259 272017 6 VPWR
port 613 nsew power input
rlabel viali s 1133 271983 1167 272017 6 VPWR
port 613 nsew power input
rlabel viali s 298753 273071 298787 273105 6 VPWR
port 613 nsew power input
rlabel viali s 298661 273071 298695 273105 6 VPWR
port 613 nsew power input
rlabel viali s 1317 273071 1340 273105 6 VPWR
port 613 nsew power input
rlabel viali s 1225 273071 1259 273105 6 VPWR
port 613 nsew power input
rlabel viali s 1133 273071 1167 273105 6 VPWR
port 613 nsew power input
rlabel viali s 298753 274159 298787 274193 6 VPWR
port 613 nsew power input
rlabel viali s 298661 274159 298695 274193 6 VPWR
port 613 nsew power input
rlabel viali s 1317 274159 1340 274193 6 VPWR
port 613 nsew power input
rlabel viali s 1225 274159 1259 274193 6 VPWR
port 613 nsew power input
rlabel viali s 1133 274159 1167 274193 6 VPWR
port 613 nsew power input
rlabel viali s 298753 275247 298787 275281 6 VPWR
port 613 nsew power input
rlabel viali s 298661 275247 298695 275281 6 VPWR
port 613 nsew power input
rlabel viali s 1317 275247 1340 275281 6 VPWR
port 613 nsew power input
rlabel viali s 1225 275247 1259 275281 6 VPWR
port 613 nsew power input
rlabel viali s 1133 275247 1167 275281 6 VPWR
port 613 nsew power input
rlabel viali s 298753 276335 298787 276369 6 VPWR
port 613 nsew power input
rlabel viali s 298661 276335 298695 276369 6 VPWR
port 613 nsew power input
rlabel viali s 1317 276335 1340 276369 6 VPWR
port 613 nsew power input
rlabel viali s 1225 276335 1259 276369 6 VPWR
port 613 nsew power input
rlabel viali s 1133 276335 1167 276369 6 VPWR
port 613 nsew power input
rlabel viali s 298753 277423 298787 277457 6 VPWR
port 613 nsew power input
rlabel viali s 298661 277423 298695 277457 6 VPWR
port 613 nsew power input
rlabel viali s 1317 277423 1340 277457 6 VPWR
port 613 nsew power input
rlabel viali s 1225 277423 1259 277457 6 VPWR
port 613 nsew power input
rlabel viali s 1133 277423 1167 277457 6 VPWR
port 613 nsew power input
rlabel viali s 298753 278511 298787 278545 6 VPWR
port 613 nsew power input
rlabel viali s 298661 278511 298695 278545 6 VPWR
port 613 nsew power input
rlabel viali s 1317 278511 1340 278545 6 VPWR
port 613 nsew power input
rlabel viali s 1225 278511 1259 278545 6 VPWR
port 613 nsew power input
rlabel viali s 1133 278511 1167 278545 6 VPWR
port 613 nsew power input
rlabel viali s 298753 279599 298787 279633 6 VPWR
port 613 nsew power input
rlabel viali s 298661 279599 298695 279633 6 VPWR
port 613 nsew power input
rlabel viali s 1317 279599 1340 279633 6 VPWR
port 613 nsew power input
rlabel viali s 1225 279599 1259 279633 6 VPWR
port 613 nsew power input
rlabel viali s 1133 279599 1167 279633 6 VPWR
port 613 nsew power input
rlabel viali s 298753 280687 298787 280721 6 VPWR
port 613 nsew power input
rlabel viali s 298661 280687 298695 280721 6 VPWR
port 613 nsew power input
rlabel viali s 1317 280687 1340 280721 6 VPWR
port 613 nsew power input
rlabel viali s 1225 280687 1259 280721 6 VPWR
port 613 nsew power input
rlabel viali s 1133 280687 1167 280721 6 VPWR
port 613 nsew power input
rlabel viali s 298753 281775 298787 281809 6 VPWR
port 613 nsew power input
rlabel viali s 298661 281775 298695 281809 6 VPWR
port 613 nsew power input
rlabel viali s 1317 281775 1340 281809 6 VPWR
port 613 nsew power input
rlabel viali s 1225 281775 1259 281809 6 VPWR
port 613 nsew power input
rlabel viali s 1133 281775 1167 281809 6 VPWR
port 613 nsew power input
rlabel viali s 298753 282863 298787 282897 6 VPWR
port 613 nsew power input
rlabel viali s 298661 282863 298695 282897 6 VPWR
port 613 nsew power input
rlabel viali s 1317 282863 1340 282897 6 VPWR
port 613 nsew power input
rlabel viali s 1225 282863 1259 282897 6 VPWR
port 613 nsew power input
rlabel viali s 1133 282863 1167 282897 6 VPWR
port 613 nsew power input
rlabel viali s 298753 283951 298787 283985 6 VPWR
port 613 nsew power input
rlabel viali s 298661 283951 298695 283985 6 VPWR
port 613 nsew power input
rlabel viali s 1317 283951 1340 283985 6 VPWR
port 613 nsew power input
rlabel viali s 1225 283951 1259 283985 6 VPWR
port 613 nsew power input
rlabel viali s 1133 283951 1167 283985 6 VPWR
port 613 nsew power input
rlabel viali s 298753 285039 298787 285073 6 VPWR
port 613 nsew power input
rlabel viali s 298661 285039 298695 285073 6 VPWR
port 613 nsew power input
rlabel viali s 1317 285039 1340 285073 6 VPWR
port 613 nsew power input
rlabel viali s 1225 285039 1259 285073 6 VPWR
port 613 nsew power input
rlabel viali s 1133 285039 1167 285073 6 VPWR
port 613 nsew power input
rlabel viali s 298753 286127 298787 286161 6 VPWR
port 613 nsew power input
rlabel viali s 298661 286127 298695 286161 6 VPWR
port 613 nsew power input
rlabel viali s 1317 286127 1340 286161 6 VPWR
port 613 nsew power input
rlabel viali s 1225 286127 1259 286161 6 VPWR
port 613 nsew power input
rlabel viali s 1133 286127 1167 286161 6 VPWR
port 613 nsew power input
rlabel viali s 298753 287215 298787 287249 6 VPWR
port 613 nsew power input
rlabel viali s 298661 287215 298695 287249 6 VPWR
port 613 nsew power input
rlabel viali s 1317 287215 1340 287249 6 VPWR
port 613 nsew power input
rlabel viali s 1225 287215 1259 287249 6 VPWR
port 613 nsew power input
rlabel viali s 1133 287215 1167 287249 6 VPWR
port 613 nsew power input
rlabel viali s 298753 288303 298787 288337 6 VPWR
port 613 nsew power input
rlabel viali s 298661 288303 298695 288337 6 VPWR
port 613 nsew power input
rlabel viali s 1317 288303 1340 288337 6 VPWR
port 613 nsew power input
rlabel viali s 1225 288303 1259 288337 6 VPWR
port 613 nsew power input
rlabel viali s 1133 288303 1167 288337 6 VPWR
port 613 nsew power input
rlabel viali s 298753 289391 298787 289425 6 VPWR
port 613 nsew power input
rlabel viali s 298661 289391 298695 289425 6 VPWR
port 613 nsew power input
rlabel viali s 1317 289391 1340 289425 6 VPWR
port 613 nsew power input
rlabel viali s 1225 289391 1259 289425 6 VPWR
port 613 nsew power input
rlabel viali s 1133 289391 1167 289425 6 VPWR
port 613 nsew power input
rlabel viali s 298753 290479 298787 290513 6 VPWR
port 613 nsew power input
rlabel viali s 298661 290479 298695 290513 6 VPWR
port 613 nsew power input
rlabel viali s 1317 290479 1340 290513 6 VPWR
port 613 nsew power input
rlabel viali s 1225 290479 1259 290513 6 VPWR
port 613 nsew power input
rlabel viali s 1133 290479 1167 290513 6 VPWR
port 613 nsew power input
rlabel viali s 298753 291567 298787 291601 6 VPWR
port 613 nsew power input
rlabel viali s 298661 291567 298695 291601 6 VPWR
port 613 nsew power input
rlabel viali s 1317 291567 1340 291601 6 VPWR
port 613 nsew power input
rlabel viali s 1225 291567 1259 291601 6 VPWR
port 613 nsew power input
rlabel viali s 1133 291567 1167 291601 6 VPWR
port 613 nsew power input
rlabel viali s 298753 292655 298787 292689 6 VPWR
port 613 nsew power input
rlabel viali s 298661 292655 298695 292689 6 VPWR
port 613 nsew power input
rlabel viali s 1317 292655 1340 292689 6 VPWR
port 613 nsew power input
rlabel viali s 1225 292655 1259 292689 6 VPWR
port 613 nsew power input
rlabel viali s 1133 292655 1167 292689 6 VPWR
port 613 nsew power input
rlabel viali s 298753 293743 298787 293777 6 VPWR
port 613 nsew power input
rlabel viali s 298661 293743 298695 293777 6 VPWR
port 613 nsew power input
rlabel viali s 1317 293743 1340 293777 6 VPWR
port 613 nsew power input
rlabel viali s 1225 293743 1259 293777 6 VPWR
port 613 nsew power input
rlabel viali s 1133 293743 1167 293777 6 VPWR
port 613 nsew power input
rlabel viali s 298753 294831 298787 294865 6 VPWR
port 613 nsew power input
rlabel viali s 298661 294831 298695 294865 6 VPWR
port 613 nsew power input
rlabel viali s 1317 294831 1340 294865 6 VPWR
port 613 nsew power input
rlabel viali s 1225 294831 1259 294865 6 VPWR
port 613 nsew power input
rlabel viali s 1133 294831 1167 294865 6 VPWR
port 613 nsew power input
rlabel viali s 298753 295919 298787 295953 6 VPWR
port 613 nsew power input
rlabel viali s 298661 295919 298695 295953 6 VPWR
port 613 nsew power input
rlabel viali s 1317 295919 1340 295953 6 VPWR
port 613 nsew power input
rlabel viali s 1225 295919 1259 295953 6 VPWR
port 613 nsew power input
rlabel viali s 1133 295919 1167 295953 6 VPWR
port 613 nsew power input
rlabel viali s 298753 297007 298787 297041 6 VPWR
port 613 nsew power input
rlabel viali s 298661 297007 298695 297041 6 VPWR
port 613 nsew power input
rlabel viali s 1317 297007 1340 297041 6 VPWR
port 613 nsew power input
rlabel viali s 1225 297007 1259 297041 6 VPWR
port 613 nsew power input
rlabel viali s 1133 297007 1167 297041 6 VPWR
port 613 nsew power input
rlabel locali s 298660 2159 298816 2193 6 VPWR
port 613 nsew power input
rlabel locali s 298660 2193 298799 2411 6 VPWR
port 613 nsew power input
rlabel locali s 298660 2411 298661 2519 6 VPWR
port 613 nsew power input
rlabel locali s 1104 2159 1340 2193 6 VPWR
port 613 nsew power input
rlabel locali s 1121 2193 1340 2411 6 VPWR
port 613 nsew power input
rlabel locali s 1259 2411 1340 2519 6 VPWR
port 613 nsew power input
rlabel locali s 298660 2921 298661 3029 6 VPWR
port 613 nsew power input
rlabel locali s 298660 3029 298799 3247 6 VPWR
port 613 nsew power input
rlabel locali s 298660 3247 298816 3281 6 VPWR
port 613 nsew power input
rlabel locali s 298660 3281 298799 3499 6 VPWR
port 613 nsew power input
rlabel locali s 298660 3499 298661 3607 6 VPWR
port 613 nsew power input
rlabel locali s 1259 2921 1340 3029 6 VPWR
port 613 nsew power input
rlabel locali s 1121 3029 1340 3247 6 VPWR
port 613 nsew power input
rlabel locali s 1104 3247 1340 3281 6 VPWR
port 613 nsew power input
rlabel locali s 1121 3281 1340 3499 6 VPWR
port 613 nsew power input
rlabel locali s 1259 3499 1340 3607 6 VPWR
port 613 nsew power input
rlabel locali s 298660 4009 298661 4117 6 VPWR
port 613 nsew power input
rlabel locali s 298660 4117 298799 4335 6 VPWR
port 613 nsew power input
rlabel locali s 298660 4335 298816 4369 6 VPWR
port 613 nsew power input
rlabel locali s 298660 4369 298799 4587 6 VPWR
port 613 nsew power input
rlabel locali s 298660 4587 298661 4695 6 VPWR
port 613 nsew power input
rlabel locali s 1259 4009 1340 4117 6 VPWR
port 613 nsew power input
rlabel locali s 1121 4117 1340 4335 6 VPWR
port 613 nsew power input
rlabel locali s 1104 4335 1340 4369 6 VPWR
port 613 nsew power input
rlabel locali s 1121 4369 1340 4587 6 VPWR
port 613 nsew power input
rlabel locali s 1259 4587 1340 4695 6 VPWR
port 613 nsew power input
rlabel locali s 298660 5097 298661 5205 6 VPWR
port 613 nsew power input
rlabel locali s 298660 5205 298799 5423 6 VPWR
port 613 nsew power input
rlabel locali s 298660 5423 298816 5457 6 VPWR
port 613 nsew power input
rlabel locali s 298660 5457 298799 5675 6 VPWR
port 613 nsew power input
rlabel locali s 298660 5675 298661 5783 6 VPWR
port 613 nsew power input
rlabel locali s 1259 5097 1340 5205 6 VPWR
port 613 nsew power input
rlabel locali s 1121 5205 1340 5423 6 VPWR
port 613 nsew power input
rlabel locali s 1104 5423 1340 5457 6 VPWR
port 613 nsew power input
rlabel locali s 1121 5457 1340 5675 6 VPWR
port 613 nsew power input
rlabel locali s 1259 5675 1340 5783 6 VPWR
port 613 nsew power input
rlabel locali s 298660 6185 298661 6293 6 VPWR
port 613 nsew power input
rlabel locali s 298660 6293 298799 6511 6 VPWR
port 613 nsew power input
rlabel locali s 298660 6511 298816 6545 6 VPWR
port 613 nsew power input
rlabel locali s 298660 6545 298799 6763 6 VPWR
port 613 nsew power input
rlabel locali s 298660 6763 298661 6871 6 VPWR
port 613 nsew power input
rlabel locali s 1259 6185 1340 6293 6 VPWR
port 613 nsew power input
rlabel locali s 1121 6293 1340 6511 6 VPWR
port 613 nsew power input
rlabel locali s 1104 6511 1340 6545 6 VPWR
port 613 nsew power input
rlabel locali s 1121 6545 1340 6763 6 VPWR
port 613 nsew power input
rlabel locali s 1259 6763 1340 6871 6 VPWR
port 613 nsew power input
rlabel locali s 298660 7273 298661 7381 6 VPWR
port 613 nsew power input
rlabel locali s 298660 7381 298799 7599 6 VPWR
port 613 nsew power input
rlabel locali s 298660 7599 298816 7633 6 VPWR
port 613 nsew power input
rlabel locali s 298660 7633 298799 7851 6 VPWR
port 613 nsew power input
rlabel locali s 298660 7851 298661 7959 6 VPWR
port 613 nsew power input
rlabel locali s 1259 7273 1340 7381 6 VPWR
port 613 nsew power input
rlabel locali s 1121 7381 1340 7599 6 VPWR
port 613 nsew power input
rlabel locali s 1104 7599 1340 7633 6 VPWR
port 613 nsew power input
rlabel locali s 1121 7633 1340 7851 6 VPWR
port 613 nsew power input
rlabel locali s 1259 7851 1340 7959 6 VPWR
port 613 nsew power input
rlabel locali s 298660 8361 298661 8469 6 VPWR
port 613 nsew power input
rlabel locali s 298660 8469 298799 8687 6 VPWR
port 613 nsew power input
rlabel locali s 298660 8687 298816 8721 6 VPWR
port 613 nsew power input
rlabel locali s 298660 8721 298799 8939 6 VPWR
port 613 nsew power input
rlabel locali s 298660 8939 298661 9047 6 VPWR
port 613 nsew power input
rlabel locali s 1259 8361 1340 8469 6 VPWR
port 613 nsew power input
rlabel locali s 1121 8469 1340 8687 6 VPWR
port 613 nsew power input
rlabel locali s 1104 8687 1340 8721 6 VPWR
port 613 nsew power input
rlabel locali s 1121 8721 1340 8939 6 VPWR
port 613 nsew power input
rlabel locali s 1259 8939 1340 9047 6 VPWR
port 613 nsew power input
rlabel locali s 298660 9449 298661 9557 6 VPWR
port 613 nsew power input
rlabel locali s 298660 9557 298799 9775 6 VPWR
port 613 nsew power input
rlabel locali s 298660 9775 298816 9809 6 VPWR
port 613 nsew power input
rlabel locali s 298660 9809 298799 10027 6 VPWR
port 613 nsew power input
rlabel locali s 298660 10027 298661 10135 6 VPWR
port 613 nsew power input
rlabel locali s 1259 9449 1340 9557 6 VPWR
port 613 nsew power input
rlabel locali s 1121 9557 1340 9775 6 VPWR
port 613 nsew power input
rlabel locali s 1104 9775 1340 9809 6 VPWR
port 613 nsew power input
rlabel locali s 1121 9809 1340 10027 6 VPWR
port 613 nsew power input
rlabel locali s 1259 10027 1340 10135 6 VPWR
port 613 nsew power input
rlabel locali s 298660 10537 298661 10645 6 VPWR
port 613 nsew power input
rlabel locali s 298660 10645 298799 10863 6 VPWR
port 613 nsew power input
rlabel locali s 298660 10863 298816 10897 6 VPWR
port 613 nsew power input
rlabel locali s 298660 10897 298799 11115 6 VPWR
port 613 nsew power input
rlabel locali s 298660 11115 298661 11223 6 VPWR
port 613 nsew power input
rlabel locali s 1259 10537 1340 10645 6 VPWR
port 613 nsew power input
rlabel locali s 1121 10645 1340 10863 6 VPWR
port 613 nsew power input
rlabel locali s 1104 10863 1340 10897 6 VPWR
port 613 nsew power input
rlabel locali s 1121 10897 1340 11115 6 VPWR
port 613 nsew power input
rlabel locali s 1259 11115 1340 11223 6 VPWR
port 613 nsew power input
rlabel locali s 298660 11625 298661 11733 6 VPWR
port 613 nsew power input
rlabel locali s 298660 11733 298799 11951 6 VPWR
port 613 nsew power input
rlabel locali s 298660 11951 298816 11985 6 VPWR
port 613 nsew power input
rlabel locali s 298660 11985 298799 12203 6 VPWR
port 613 nsew power input
rlabel locali s 298660 12203 298661 12311 6 VPWR
port 613 nsew power input
rlabel locali s 1259 11625 1340 11733 6 VPWR
port 613 nsew power input
rlabel locali s 1121 11733 1340 11951 6 VPWR
port 613 nsew power input
rlabel locali s 1104 11951 1340 11985 6 VPWR
port 613 nsew power input
rlabel locali s 1121 11985 1340 12203 6 VPWR
port 613 nsew power input
rlabel locali s 1259 12203 1340 12311 6 VPWR
port 613 nsew power input
rlabel locali s 298660 12713 298661 12821 6 VPWR
port 613 nsew power input
rlabel locali s 298660 12821 298799 13039 6 VPWR
port 613 nsew power input
rlabel locali s 298660 13039 298816 13073 6 VPWR
port 613 nsew power input
rlabel locali s 298660 13073 298799 13291 6 VPWR
port 613 nsew power input
rlabel locali s 298660 13291 298661 13399 6 VPWR
port 613 nsew power input
rlabel locali s 1259 12713 1340 12821 6 VPWR
port 613 nsew power input
rlabel locali s 1121 12821 1340 13039 6 VPWR
port 613 nsew power input
rlabel locali s 1104 13039 1340 13073 6 VPWR
port 613 nsew power input
rlabel locali s 1121 13073 1340 13291 6 VPWR
port 613 nsew power input
rlabel locali s 1259 13291 1340 13399 6 VPWR
port 613 nsew power input
rlabel locali s 298660 13801 298661 13909 6 VPWR
port 613 nsew power input
rlabel locali s 298660 13909 298799 14127 6 VPWR
port 613 nsew power input
rlabel locali s 298660 14127 298816 14161 6 VPWR
port 613 nsew power input
rlabel locali s 298660 14161 298799 14379 6 VPWR
port 613 nsew power input
rlabel locali s 298660 14379 298661 14487 6 VPWR
port 613 nsew power input
rlabel locali s 1259 13801 1340 13909 6 VPWR
port 613 nsew power input
rlabel locali s 1121 13909 1340 14127 6 VPWR
port 613 nsew power input
rlabel locali s 1104 14127 1340 14161 6 VPWR
port 613 nsew power input
rlabel locali s 1121 14161 1340 14379 6 VPWR
port 613 nsew power input
rlabel locali s 1259 14379 1340 14487 6 VPWR
port 613 nsew power input
rlabel locali s 298660 14889 298661 14997 6 VPWR
port 613 nsew power input
rlabel locali s 298660 14997 298799 15215 6 VPWR
port 613 nsew power input
rlabel locali s 298660 15215 298816 15249 6 VPWR
port 613 nsew power input
rlabel locali s 298660 15249 298799 15467 6 VPWR
port 613 nsew power input
rlabel locali s 298660 15467 298661 15575 6 VPWR
port 613 nsew power input
rlabel locali s 1259 14889 1340 14997 6 VPWR
port 613 nsew power input
rlabel locali s 1121 14997 1340 15215 6 VPWR
port 613 nsew power input
rlabel locali s 1104 15215 1340 15249 6 VPWR
port 613 nsew power input
rlabel locali s 1121 15249 1340 15467 6 VPWR
port 613 nsew power input
rlabel locali s 1259 15467 1340 15575 6 VPWR
port 613 nsew power input
rlabel locali s 298660 15977 298661 16085 6 VPWR
port 613 nsew power input
rlabel locali s 298660 16085 298799 16303 6 VPWR
port 613 nsew power input
rlabel locali s 298660 16303 298816 16337 6 VPWR
port 613 nsew power input
rlabel locali s 298660 16337 298799 16555 6 VPWR
port 613 nsew power input
rlabel locali s 298660 16555 298661 16663 6 VPWR
port 613 nsew power input
rlabel locali s 1259 15977 1340 16085 6 VPWR
port 613 nsew power input
rlabel locali s 1121 16085 1340 16303 6 VPWR
port 613 nsew power input
rlabel locali s 1104 16303 1340 16337 6 VPWR
port 613 nsew power input
rlabel locali s 1121 16337 1340 16555 6 VPWR
port 613 nsew power input
rlabel locali s 1259 16555 1340 16663 6 VPWR
port 613 nsew power input
rlabel locali s 298660 17065 298661 17173 6 VPWR
port 613 nsew power input
rlabel locali s 298660 17173 298799 17391 6 VPWR
port 613 nsew power input
rlabel locali s 298660 17391 298816 17425 6 VPWR
port 613 nsew power input
rlabel locali s 298660 17425 298799 17643 6 VPWR
port 613 nsew power input
rlabel locali s 298660 17643 298661 17751 6 VPWR
port 613 nsew power input
rlabel locali s 1259 17065 1340 17173 6 VPWR
port 613 nsew power input
rlabel locali s 1121 17173 1340 17391 6 VPWR
port 613 nsew power input
rlabel locali s 1104 17391 1340 17425 6 VPWR
port 613 nsew power input
rlabel locali s 1121 17425 1340 17643 6 VPWR
port 613 nsew power input
rlabel locali s 1259 17643 1340 17751 6 VPWR
port 613 nsew power input
rlabel locali s 298660 18153 298661 18261 6 VPWR
port 613 nsew power input
rlabel locali s 298660 18261 298799 18479 6 VPWR
port 613 nsew power input
rlabel locali s 298660 18479 298816 18513 6 VPWR
port 613 nsew power input
rlabel locali s 298660 18513 298799 18731 6 VPWR
port 613 nsew power input
rlabel locali s 298660 18731 298661 18839 6 VPWR
port 613 nsew power input
rlabel locali s 1259 18153 1340 18261 6 VPWR
port 613 nsew power input
rlabel locali s 1121 18261 1340 18479 6 VPWR
port 613 nsew power input
rlabel locali s 1104 18479 1340 18513 6 VPWR
port 613 nsew power input
rlabel locali s 1121 18513 1340 18731 6 VPWR
port 613 nsew power input
rlabel locali s 1259 18731 1340 18839 6 VPWR
port 613 nsew power input
rlabel locali s 298660 19241 298661 19349 6 VPWR
port 613 nsew power input
rlabel locali s 298660 19349 298799 19567 6 VPWR
port 613 nsew power input
rlabel locali s 298660 19567 298816 19601 6 VPWR
port 613 nsew power input
rlabel locali s 298660 19601 298799 19819 6 VPWR
port 613 nsew power input
rlabel locali s 298660 19819 298661 19927 6 VPWR
port 613 nsew power input
rlabel locali s 1259 19241 1340 19349 6 VPWR
port 613 nsew power input
rlabel locali s 1121 19349 1340 19567 6 VPWR
port 613 nsew power input
rlabel locali s 1104 19567 1340 19601 6 VPWR
port 613 nsew power input
rlabel locali s 1121 19601 1340 19819 6 VPWR
port 613 nsew power input
rlabel locali s 1259 19819 1340 19927 6 VPWR
port 613 nsew power input
rlabel locali s 298660 20329 298661 20437 6 VPWR
port 613 nsew power input
rlabel locali s 298660 20437 298799 20655 6 VPWR
port 613 nsew power input
rlabel locali s 298660 20655 298816 20689 6 VPWR
port 613 nsew power input
rlabel locali s 298660 20689 298799 20907 6 VPWR
port 613 nsew power input
rlabel locali s 298660 20907 298661 21015 6 VPWR
port 613 nsew power input
rlabel locali s 1259 20329 1340 20437 6 VPWR
port 613 nsew power input
rlabel locali s 1121 20437 1340 20655 6 VPWR
port 613 nsew power input
rlabel locali s 1104 20655 1340 20689 6 VPWR
port 613 nsew power input
rlabel locali s 1121 20689 1340 20907 6 VPWR
port 613 nsew power input
rlabel locali s 1259 20907 1340 21015 6 VPWR
port 613 nsew power input
rlabel locali s 298660 21417 298661 21525 6 VPWR
port 613 nsew power input
rlabel locali s 298660 21525 298799 21743 6 VPWR
port 613 nsew power input
rlabel locali s 298660 21743 298816 21777 6 VPWR
port 613 nsew power input
rlabel locali s 298660 21777 298799 21995 6 VPWR
port 613 nsew power input
rlabel locali s 298660 21995 298661 22103 6 VPWR
port 613 nsew power input
rlabel locali s 1259 21417 1340 21525 6 VPWR
port 613 nsew power input
rlabel locali s 1121 21525 1340 21743 6 VPWR
port 613 nsew power input
rlabel locali s 1104 21743 1340 21777 6 VPWR
port 613 nsew power input
rlabel locali s 1121 21777 1340 21995 6 VPWR
port 613 nsew power input
rlabel locali s 1259 21995 1340 22103 6 VPWR
port 613 nsew power input
rlabel locali s 298660 22505 298661 22613 6 VPWR
port 613 nsew power input
rlabel locali s 298660 22613 298799 22831 6 VPWR
port 613 nsew power input
rlabel locali s 298660 22831 298816 22865 6 VPWR
port 613 nsew power input
rlabel locali s 298660 22865 298799 23083 6 VPWR
port 613 nsew power input
rlabel locali s 298660 23083 298661 23191 6 VPWR
port 613 nsew power input
rlabel locali s 1259 22505 1340 22613 6 VPWR
port 613 nsew power input
rlabel locali s 1121 22613 1340 22831 6 VPWR
port 613 nsew power input
rlabel locali s 1104 22831 1340 22865 6 VPWR
port 613 nsew power input
rlabel locali s 1121 22865 1340 23083 6 VPWR
port 613 nsew power input
rlabel locali s 1259 23083 1340 23191 6 VPWR
port 613 nsew power input
rlabel locali s 298660 23593 298661 23701 6 VPWR
port 613 nsew power input
rlabel locali s 298660 23701 298799 23919 6 VPWR
port 613 nsew power input
rlabel locali s 298660 23919 298816 23953 6 VPWR
port 613 nsew power input
rlabel locali s 298660 23953 298799 24171 6 VPWR
port 613 nsew power input
rlabel locali s 298660 24171 298661 24279 6 VPWR
port 613 nsew power input
rlabel locali s 1259 23593 1340 23701 6 VPWR
port 613 nsew power input
rlabel locali s 1121 23701 1340 23919 6 VPWR
port 613 nsew power input
rlabel locali s 1104 23919 1340 23953 6 VPWR
port 613 nsew power input
rlabel locali s 1121 23953 1340 24171 6 VPWR
port 613 nsew power input
rlabel locali s 1259 24171 1340 24279 6 VPWR
port 613 nsew power input
rlabel locali s 298660 24681 298661 24789 6 VPWR
port 613 nsew power input
rlabel locali s 298660 24789 298799 25007 6 VPWR
port 613 nsew power input
rlabel locali s 298660 25007 298816 25041 6 VPWR
port 613 nsew power input
rlabel locali s 298660 25041 298799 25259 6 VPWR
port 613 nsew power input
rlabel locali s 298660 25259 298661 25367 6 VPWR
port 613 nsew power input
rlabel locali s 1259 24681 1340 24789 6 VPWR
port 613 nsew power input
rlabel locali s 1121 24789 1340 25007 6 VPWR
port 613 nsew power input
rlabel locali s 1104 25007 1340 25041 6 VPWR
port 613 nsew power input
rlabel locali s 1121 25041 1340 25259 6 VPWR
port 613 nsew power input
rlabel locali s 1259 25259 1340 25367 6 VPWR
port 613 nsew power input
rlabel locali s 298660 25769 298661 25877 6 VPWR
port 613 nsew power input
rlabel locali s 298660 25877 298799 26095 6 VPWR
port 613 nsew power input
rlabel locali s 298660 26095 298816 26129 6 VPWR
port 613 nsew power input
rlabel locali s 298660 26129 298799 26347 6 VPWR
port 613 nsew power input
rlabel locali s 298660 26347 298661 26455 6 VPWR
port 613 nsew power input
rlabel locali s 1259 25769 1340 25877 6 VPWR
port 613 nsew power input
rlabel locali s 1121 25877 1340 26095 6 VPWR
port 613 nsew power input
rlabel locali s 1104 26095 1340 26129 6 VPWR
port 613 nsew power input
rlabel locali s 1121 26129 1340 26347 6 VPWR
port 613 nsew power input
rlabel locali s 1259 26347 1340 26455 6 VPWR
port 613 nsew power input
rlabel locali s 298660 26857 298661 26965 6 VPWR
port 613 nsew power input
rlabel locali s 298660 26965 298799 27183 6 VPWR
port 613 nsew power input
rlabel locali s 298660 27183 298816 27217 6 VPWR
port 613 nsew power input
rlabel locali s 298660 27217 298799 27435 6 VPWR
port 613 nsew power input
rlabel locali s 298660 27435 298661 27543 6 VPWR
port 613 nsew power input
rlabel locali s 1259 26857 1340 26965 6 VPWR
port 613 nsew power input
rlabel locali s 1121 26965 1340 27183 6 VPWR
port 613 nsew power input
rlabel locali s 1104 27183 1340 27217 6 VPWR
port 613 nsew power input
rlabel locali s 1121 27217 1340 27435 6 VPWR
port 613 nsew power input
rlabel locali s 1259 27435 1340 27543 6 VPWR
port 613 nsew power input
rlabel locali s 298660 27945 298661 28053 6 VPWR
port 613 nsew power input
rlabel locali s 298660 28053 298799 28271 6 VPWR
port 613 nsew power input
rlabel locali s 298660 28271 298816 28305 6 VPWR
port 613 nsew power input
rlabel locali s 298660 28305 298799 28523 6 VPWR
port 613 nsew power input
rlabel locali s 298660 28523 298661 28631 6 VPWR
port 613 nsew power input
rlabel locali s 1259 27945 1340 28053 6 VPWR
port 613 nsew power input
rlabel locali s 1121 28053 1340 28271 6 VPWR
port 613 nsew power input
rlabel locali s 1104 28271 1340 28305 6 VPWR
port 613 nsew power input
rlabel locali s 1121 28305 1340 28523 6 VPWR
port 613 nsew power input
rlabel locali s 1259 28523 1340 28631 6 VPWR
port 613 nsew power input
rlabel locali s 298660 29033 298661 29141 6 VPWR
port 613 nsew power input
rlabel locali s 298660 29141 298799 29359 6 VPWR
port 613 nsew power input
rlabel locali s 298660 29359 298816 29393 6 VPWR
port 613 nsew power input
rlabel locali s 298660 29393 298799 29611 6 VPWR
port 613 nsew power input
rlabel locali s 298660 29611 298661 29719 6 VPWR
port 613 nsew power input
rlabel locali s 1259 29033 1340 29141 6 VPWR
port 613 nsew power input
rlabel locali s 1121 29141 1340 29359 6 VPWR
port 613 nsew power input
rlabel locali s 1104 29359 1340 29393 6 VPWR
port 613 nsew power input
rlabel locali s 1121 29393 1340 29611 6 VPWR
port 613 nsew power input
rlabel locali s 1259 29611 1340 29719 6 VPWR
port 613 nsew power input
rlabel locali s 298660 30121 298661 30229 6 VPWR
port 613 nsew power input
rlabel locali s 298660 30229 298799 30447 6 VPWR
port 613 nsew power input
rlabel locali s 298660 30447 298816 30481 6 VPWR
port 613 nsew power input
rlabel locali s 298660 30481 298799 30699 6 VPWR
port 613 nsew power input
rlabel locali s 298660 30699 298661 30807 6 VPWR
port 613 nsew power input
rlabel locali s 1259 30121 1340 30229 6 VPWR
port 613 nsew power input
rlabel locali s 1121 30229 1340 30447 6 VPWR
port 613 nsew power input
rlabel locali s 1104 30447 1340 30481 6 VPWR
port 613 nsew power input
rlabel locali s 1121 30481 1340 30699 6 VPWR
port 613 nsew power input
rlabel locali s 1259 30699 1340 30807 6 VPWR
port 613 nsew power input
rlabel locali s 298660 31209 298661 31317 6 VPWR
port 613 nsew power input
rlabel locali s 298660 31317 298799 31535 6 VPWR
port 613 nsew power input
rlabel locali s 298660 31535 298816 31569 6 VPWR
port 613 nsew power input
rlabel locali s 298660 31569 298799 31787 6 VPWR
port 613 nsew power input
rlabel locali s 298660 31787 298661 31895 6 VPWR
port 613 nsew power input
rlabel locali s 1259 31209 1340 31317 6 VPWR
port 613 nsew power input
rlabel locali s 1121 31317 1340 31535 6 VPWR
port 613 nsew power input
rlabel locali s 1104 31535 1340 31569 6 VPWR
port 613 nsew power input
rlabel locali s 1121 31569 1340 31787 6 VPWR
port 613 nsew power input
rlabel locali s 1259 31787 1340 31895 6 VPWR
port 613 nsew power input
rlabel locali s 298660 32297 298661 32405 6 VPWR
port 613 nsew power input
rlabel locali s 298660 32405 298799 32623 6 VPWR
port 613 nsew power input
rlabel locali s 298660 32623 298816 32657 6 VPWR
port 613 nsew power input
rlabel locali s 298660 32657 298799 32875 6 VPWR
port 613 nsew power input
rlabel locali s 298660 32875 298661 32983 6 VPWR
port 613 nsew power input
rlabel locali s 1259 32297 1340 32405 6 VPWR
port 613 nsew power input
rlabel locali s 1121 32405 1340 32623 6 VPWR
port 613 nsew power input
rlabel locali s 1104 32623 1340 32657 6 VPWR
port 613 nsew power input
rlabel locali s 1121 32657 1340 32875 6 VPWR
port 613 nsew power input
rlabel locali s 1259 32875 1340 32983 6 VPWR
port 613 nsew power input
rlabel locali s 298660 33385 298661 33493 6 VPWR
port 613 nsew power input
rlabel locali s 298660 33493 298799 33711 6 VPWR
port 613 nsew power input
rlabel locali s 298660 33711 298816 33745 6 VPWR
port 613 nsew power input
rlabel locali s 298660 33745 298799 33963 6 VPWR
port 613 nsew power input
rlabel locali s 298660 33963 298661 34071 6 VPWR
port 613 nsew power input
rlabel locali s 1259 33385 1340 33493 6 VPWR
port 613 nsew power input
rlabel locali s 1121 33493 1340 33711 6 VPWR
port 613 nsew power input
rlabel locali s 1104 33711 1340 33745 6 VPWR
port 613 nsew power input
rlabel locali s 1121 33745 1340 33963 6 VPWR
port 613 nsew power input
rlabel locali s 1259 33963 1340 34071 6 VPWR
port 613 nsew power input
rlabel locali s 298660 34473 298661 34581 6 VPWR
port 613 nsew power input
rlabel locali s 298660 34581 298799 34799 6 VPWR
port 613 nsew power input
rlabel locali s 298660 34799 298816 34833 6 VPWR
port 613 nsew power input
rlabel locali s 298660 34833 298799 35051 6 VPWR
port 613 nsew power input
rlabel locali s 298660 35051 298661 35159 6 VPWR
port 613 nsew power input
rlabel locali s 1259 34473 1340 34581 6 VPWR
port 613 nsew power input
rlabel locali s 1121 34581 1340 34799 6 VPWR
port 613 nsew power input
rlabel locali s 1104 34799 1340 34833 6 VPWR
port 613 nsew power input
rlabel locali s 1121 34833 1340 35051 6 VPWR
port 613 nsew power input
rlabel locali s 1259 35051 1340 35159 6 VPWR
port 613 nsew power input
rlabel locali s 298660 35561 298661 35669 6 VPWR
port 613 nsew power input
rlabel locali s 298660 35669 298799 35887 6 VPWR
port 613 nsew power input
rlabel locali s 298660 35887 298816 35921 6 VPWR
port 613 nsew power input
rlabel locali s 298660 35921 298799 36139 6 VPWR
port 613 nsew power input
rlabel locali s 298660 36139 298661 36247 6 VPWR
port 613 nsew power input
rlabel locali s 1259 35561 1340 35669 6 VPWR
port 613 nsew power input
rlabel locali s 1121 35669 1340 35887 6 VPWR
port 613 nsew power input
rlabel locali s 1104 35887 1340 35921 6 VPWR
port 613 nsew power input
rlabel locali s 1121 35921 1340 36139 6 VPWR
port 613 nsew power input
rlabel locali s 1259 36139 1340 36247 6 VPWR
port 613 nsew power input
rlabel locali s 298660 36649 298661 36757 6 VPWR
port 613 nsew power input
rlabel locali s 298660 36757 298799 36975 6 VPWR
port 613 nsew power input
rlabel locali s 298660 36975 298816 37009 6 VPWR
port 613 nsew power input
rlabel locali s 298660 37009 298799 37227 6 VPWR
port 613 nsew power input
rlabel locali s 298660 37227 298661 37335 6 VPWR
port 613 nsew power input
rlabel locali s 1259 36649 1340 36757 6 VPWR
port 613 nsew power input
rlabel locali s 1121 36757 1340 36975 6 VPWR
port 613 nsew power input
rlabel locali s 1104 36975 1340 37009 6 VPWR
port 613 nsew power input
rlabel locali s 1121 37009 1340 37227 6 VPWR
port 613 nsew power input
rlabel locali s 1259 37227 1340 37335 6 VPWR
port 613 nsew power input
rlabel locali s 298660 37737 298661 37845 6 VPWR
port 613 nsew power input
rlabel locali s 298660 37845 298799 38063 6 VPWR
port 613 nsew power input
rlabel locali s 298660 38063 298816 38097 6 VPWR
port 613 nsew power input
rlabel locali s 298660 38097 298799 38315 6 VPWR
port 613 nsew power input
rlabel locali s 298660 38315 298661 38423 6 VPWR
port 613 nsew power input
rlabel locali s 1259 37737 1340 37845 6 VPWR
port 613 nsew power input
rlabel locali s 1121 37845 1340 38063 6 VPWR
port 613 nsew power input
rlabel locali s 1104 38063 1340 38097 6 VPWR
port 613 nsew power input
rlabel locali s 1121 38097 1340 38315 6 VPWR
port 613 nsew power input
rlabel locali s 1259 38315 1340 38423 6 VPWR
port 613 nsew power input
rlabel locali s 298660 38825 298661 38933 6 VPWR
port 613 nsew power input
rlabel locali s 298660 38933 298799 39151 6 VPWR
port 613 nsew power input
rlabel locali s 298660 39151 298816 39185 6 VPWR
port 613 nsew power input
rlabel locali s 298660 39185 298799 39403 6 VPWR
port 613 nsew power input
rlabel locali s 298660 39403 298661 39511 6 VPWR
port 613 nsew power input
rlabel locali s 1259 38825 1340 38933 6 VPWR
port 613 nsew power input
rlabel locali s 1121 38933 1340 39151 6 VPWR
port 613 nsew power input
rlabel locali s 1104 39151 1340 39185 6 VPWR
port 613 nsew power input
rlabel locali s 1121 39185 1340 39403 6 VPWR
port 613 nsew power input
rlabel locali s 1259 39403 1340 39511 6 VPWR
port 613 nsew power input
rlabel locali s 298660 39913 298661 40021 6 VPWR
port 613 nsew power input
rlabel locali s 298660 40021 298799 40239 6 VPWR
port 613 nsew power input
rlabel locali s 298660 40239 298816 40273 6 VPWR
port 613 nsew power input
rlabel locali s 298660 40273 298799 40491 6 VPWR
port 613 nsew power input
rlabel locali s 298660 40491 298661 40599 6 VPWR
port 613 nsew power input
rlabel locali s 1259 39913 1340 40021 6 VPWR
port 613 nsew power input
rlabel locali s 1121 40021 1340 40239 6 VPWR
port 613 nsew power input
rlabel locali s 1104 40239 1340 40273 6 VPWR
port 613 nsew power input
rlabel locali s 1121 40273 1340 40491 6 VPWR
port 613 nsew power input
rlabel locali s 1259 40491 1340 40599 6 VPWR
port 613 nsew power input
rlabel locali s 298660 41001 298661 41109 6 VPWR
port 613 nsew power input
rlabel locali s 298660 41109 298799 41327 6 VPWR
port 613 nsew power input
rlabel locali s 298660 41327 298816 41361 6 VPWR
port 613 nsew power input
rlabel locali s 298660 41361 298799 41579 6 VPWR
port 613 nsew power input
rlabel locali s 298660 41579 298661 41687 6 VPWR
port 613 nsew power input
rlabel locali s 1259 41001 1340 41109 6 VPWR
port 613 nsew power input
rlabel locali s 1121 41109 1340 41327 6 VPWR
port 613 nsew power input
rlabel locali s 1104 41327 1340 41361 6 VPWR
port 613 nsew power input
rlabel locali s 1121 41361 1340 41579 6 VPWR
port 613 nsew power input
rlabel locali s 1259 41579 1340 41687 6 VPWR
port 613 nsew power input
rlabel locali s 298660 42089 298661 42197 6 VPWR
port 613 nsew power input
rlabel locali s 298660 42197 298799 42415 6 VPWR
port 613 nsew power input
rlabel locali s 298660 42415 298816 42449 6 VPWR
port 613 nsew power input
rlabel locali s 298660 42449 298799 42667 6 VPWR
port 613 nsew power input
rlabel locali s 298660 42667 298661 42775 6 VPWR
port 613 nsew power input
rlabel locali s 1259 42089 1340 42197 6 VPWR
port 613 nsew power input
rlabel locali s 1121 42197 1340 42415 6 VPWR
port 613 nsew power input
rlabel locali s 1104 42415 1340 42449 6 VPWR
port 613 nsew power input
rlabel locali s 1121 42449 1340 42667 6 VPWR
port 613 nsew power input
rlabel locali s 1259 42667 1340 42775 6 VPWR
port 613 nsew power input
rlabel locali s 298660 43177 298661 43285 6 VPWR
port 613 nsew power input
rlabel locali s 298660 43285 298799 43503 6 VPWR
port 613 nsew power input
rlabel locali s 298660 43503 298816 43537 6 VPWR
port 613 nsew power input
rlabel locali s 298660 43537 298799 43755 6 VPWR
port 613 nsew power input
rlabel locali s 298660 43755 298661 43863 6 VPWR
port 613 nsew power input
rlabel locali s 1259 43177 1340 43285 6 VPWR
port 613 nsew power input
rlabel locali s 1121 43285 1340 43503 6 VPWR
port 613 nsew power input
rlabel locali s 1104 43503 1340 43537 6 VPWR
port 613 nsew power input
rlabel locali s 1121 43537 1340 43755 6 VPWR
port 613 nsew power input
rlabel locali s 1259 43755 1340 43863 6 VPWR
port 613 nsew power input
rlabel locali s 298660 44265 298661 44373 6 VPWR
port 613 nsew power input
rlabel locali s 298660 44373 298799 44591 6 VPWR
port 613 nsew power input
rlabel locali s 298660 44591 298816 44625 6 VPWR
port 613 nsew power input
rlabel locali s 298660 44625 298799 44843 6 VPWR
port 613 nsew power input
rlabel locali s 298660 44843 298661 44951 6 VPWR
port 613 nsew power input
rlabel locali s 1259 44265 1340 44373 6 VPWR
port 613 nsew power input
rlabel locali s 1121 44373 1340 44591 6 VPWR
port 613 nsew power input
rlabel locali s 1104 44591 1340 44625 6 VPWR
port 613 nsew power input
rlabel locali s 1121 44625 1340 44843 6 VPWR
port 613 nsew power input
rlabel locali s 1259 44843 1340 44951 6 VPWR
port 613 nsew power input
rlabel locali s 298660 45353 298661 45461 6 VPWR
port 613 nsew power input
rlabel locali s 298660 45461 298799 45679 6 VPWR
port 613 nsew power input
rlabel locali s 298660 45679 298816 45713 6 VPWR
port 613 nsew power input
rlabel locali s 298660 45713 298799 45931 6 VPWR
port 613 nsew power input
rlabel locali s 298660 45931 298661 46039 6 VPWR
port 613 nsew power input
rlabel locali s 1259 45353 1340 45461 6 VPWR
port 613 nsew power input
rlabel locali s 1121 45461 1340 45679 6 VPWR
port 613 nsew power input
rlabel locali s 1104 45679 1340 45713 6 VPWR
port 613 nsew power input
rlabel locali s 1121 45713 1340 45931 6 VPWR
port 613 nsew power input
rlabel locali s 1259 45931 1340 46039 6 VPWR
port 613 nsew power input
rlabel locali s 298660 46441 298661 46549 6 VPWR
port 613 nsew power input
rlabel locali s 298660 46549 298799 46767 6 VPWR
port 613 nsew power input
rlabel locali s 298660 46767 298816 46801 6 VPWR
port 613 nsew power input
rlabel locali s 298660 46801 298799 47019 6 VPWR
port 613 nsew power input
rlabel locali s 298660 47019 298661 47127 6 VPWR
port 613 nsew power input
rlabel locali s 1259 46441 1340 46549 6 VPWR
port 613 nsew power input
rlabel locali s 1121 46549 1340 46767 6 VPWR
port 613 nsew power input
rlabel locali s 1104 46767 1340 46801 6 VPWR
port 613 nsew power input
rlabel locali s 1121 46801 1340 47019 6 VPWR
port 613 nsew power input
rlabel locali s 1259 47019 1340 47127 6 VPWR
port 613 nsew power input
rlabel locali s 298660 47529 298661 47637 6 VPWR
port 613 nsew power input
rlabel locali s 298660 47637 298799 47855 6 VPWR
port 613 nsew power input
rlabel locali s 298660 47855 298816 47889 6 VPWR
port 613 nsew power input
rlabel locali s 298660 47889 298799 48107 6 VPWR
port 613 nsew power input
rlabel locali s 298660 48107 298661 48215 6 VPWR
port 613 nsew power input
rlabel locali s 1259 47529 1340 47637 6 VPWR
port 613 nsew power input
rlabel locali s 1121 47637 1340 47855 6 VPWR
port 613 nsew power input
rlabel locali s 1104 47855 1340 47889 6 VPWR
port 613 nsew power input
rlabel locali s 1121 47889 1340 48107 6 VPWR
port 613 nsew power input
rlabel locali s 1259 48107 1340 48215 6 VPWR
port 613 nsew power input
rlabel locali s 298660 48617 298661 48725 6 VPWR
port 613 nsew power input
rlabel locali s 298660 48725 298799 48943 6 VPWR
port 613 nsew power input
rlabel locali s 298660 48943 298816 48977 6 VPWR
port 613 nsew power input
rlabel locali s 298660 48977 298799 49195 6 VPWR
port 613 nsew power input
rlabel locali s 298660 49195 298661 49303 6 VPWR
port 613 nsew power input
rlabel locali s 1259 48617 1340 48725 6 VPWR
port 613 nsew power input
rlabel locali s 1121 48725 1340 48943 6 VPWR
port 613 nsew power input
rlabel locali s 1104 48943 1340 48977 6 VPWR
port 613 nsew power input
rlabel locali s 1121 48977 1340 49195 6 VPWR
port 613 nsew power input
rlabel locali s 1259 49195 1340 49303 6 VPWR
port 613 nsew power input
rlabel locali s 298660 49705 298661 49813 6 VPWR
port 613 nsew power input
rlabel locali s 298660 49813 298799 50031 6 VPWR
port 613 nsew power input
rlabel locali s 298660 50031 298816 50065 6 VPWR
port 613 nsew power input
rlabel locali s 298660 50065 298799 50283 6 VPWR
port 613 nsew power input
rlabel locali s 298660 50283 298661 50391 6 VPWR
port 613 nsew power input
rlabel locali s 1259 49705 1340 49813 6 VPWR
port 613 nsew power input
rlabel locali s 1121 49813 1340 50031 6 VPWR
port 613 nsew power input
rlabel locali s 1104 50031 1340 50065 6 VPWR
port 613 nsew power input
rlabel locali s 1121 50065 1340 50283 6 VPWR
port 613 nsew power input
rlabel locali s 1259 50283 1340 50391 6 VPWR
port 613 nsew power input
rlabel locali s 298660 50793 298661 50901 6 VPWR
port 613 nsew power input
rlabel locali s 298660 50901 298799 51119 6 VPWR
port 613 nsew power input
rlabel locali s 298660 51119 298816 51153 6 VPWR
port 613 nsew power input
rlabel locali s 298660 51153 298799 51371 6 VPWR
port 613 nsew power input
rlabel locali s 298660 51371 298661 51479 6 VPWR
port 613 nsew power input
rlabel locali s 1259 50793 1340 50901 6 VPWR
port 613 nsew power input
rlabel locali s 1121 50901 1340 51119 6 VPWR
port 613 nsew power input
rlabel locali s 1104 51119 1340 51153 6 VPWR
port 613 nsew power input
rlabel locali s 1121 51153 1340 51371 6 VPWR
port 613 nsew power input
rlabel locali s 1259 51371 1340 51479 6 VPWR
port 613 nsew power input
rlabel locali s 298660 51881 298661 51989 6 VPWR
port 613 nsew power input
rlabel locali s 298660 51989 298799 52207 6 VPWR
port 613 nsew power input
rlabel locali s 298660 52207 298816 52241 6 VPWR
port 613 nsew power input
rlabel locali s 298660 52241 298799 52459 6 VPWR
port 613 nsew power input
rlabel locali s 298660 52459 298661 52567 6 VPWR
port 613 nsew power input
rlabel locali s 1259 51881 1340 51989 6 VPWR
port 613 nsew power input
rlabel locali s 1121 51989 1340 52207 6 VPWR
port 613 nsew power input
rlabel locali s 1104 52207 1340 52241 6 VPWR
port 613 nsew power input
rlabel locali s 1121 52241 1340 52459 6 VPWR
port 613 nsew power input
rlabel locali s 1259 52459 1340 52567 6 VPWR
port 613 nsew power input
rlabel locali s 298660 52969 298661 53077 6 VPWR
port 613 nsew power input
rlabel locali s 298660 53077 298799 53295 6 VPWR
port 613 nsew power input
rlabel locali s 298660 53295 298816 53329 6 VPWR
port 613 nsew power input
rlabel locali s 298660 53329 298799 53547 6 VPWR
port 613 nsew power input
rlabel locali s 298660 53547 298661 53655 6 VPWR
port 613 nsew power input
rlabel locali s 1259 52969 1340 53077 6 VPWR
port 613 nsew power input
rlabel locali s 1121 53077 1340 53295 6 VPWR
port 613 nsew power input
rlabel locali s 1104 53295 1340 53329 6 VPWR
port 613 nsew power input
rlabel locali s 1121 53329 1340 53547 6 VPWR
port 613 nsew power input
rlabel locali s 1259 53547 1340 53655 6 VPWR
port 613 nsew power input
rlabel locali s 298660 54057 298661 54165 6 VPWR
port 613 nsew power input
rlabel locali s 298660 54165 298799 54383 6 VPWR
port 613 nsew power input
rlabel locali s 298660 54383 298816 54417 6 VPWR
port 613 nsew power input
rlabel locali s 298660 54417 298799 54635 6 VPWR
port 613 nsew power input
rlabel locali s 298660 54635 298661 54743 6 VPWR
port 613 nsew power input
rlabel locali s 1259 54057 1340 54165 6 VPWR
port 613 nsew power input
rlabel locali s 1121 54165 1340 54383 6 VPWR
port 613 nsew power input
rlabel locali s 1104 54383 1340 54417 6 VPWR
port 613 nsew power input
rlabel locali s 1121 54417 1340 54635 6 VPWR
port 613 nsew power input
rlabel locali s 1259 54635 1340 54743 6 VPWR
port 613 nsew power input
rlabel locali s 298660 55145 298661 55253 6 VPWR
port 613 nsew power input
rlabel locali s 298660 55253 298799 55471 6 VPWR
port 613 nsew power input
rlabel locali s 298660 55471 298816 55505 6 VPWR
port 613 nsew power input
rlabel locali s 298660 55505 298799 55723 6 VPWR
port 613 nsew power input
rlabel locali s 298660 55723 298661 55831 6 VPWR
port 613 nsew power input
rlabel locali s 1259 55145 1340 55253 6 VPWR
port 613 nsew power input
rlabel locali s 1121 55253 1340 55471 6 VPWR
port 613 nsew power input
rlabel locali s 1104 55471 1340 55505 6 VPWR
port 613 nsew power input
rlabel locali s 1121 55505 1340 55723 6 VPWR
port 613 nsew power input
rlabel locali s 1259 55723 1340 55831 6 VPWR
port 613 nsew power input
rlabel locali s 298660 56233 298661 56341 6 VPWR
port 613 nsew power input
rlabel locali s 298660 56341 298799 56559 6 VPWR
port 613 nsew power input
rlabel locali s 298660 56559 298816 56593 6 VPWR
port 613 nsew power input
rlabel locali s 298660 56593 298799 56811 6 VPWR
port 613 nsew power input
rlabel locali s 298660 56811 298661 56919 6 VPWR
port 613 nsew power input
rlabel locali s 1259 56233 1340 56341 6 VPWR
port 613 nsew power input
rlabel locali s 1121 56341 1340 56559 6 VPWR
port 613 nsew power input
rlabel locali s 1104 56559 1340 56593 6 VPWR
port 613 nsew power input
rlabel locali s 1121 56593 1340 56811 6 VPWR
port 613 nsew power input
rlabel locali s 1259 56811 1340 56919 6 VPWR
port 613 nsew power input
rlabel locali s 298660 57321 298661 57429 6 VPWR
port 613 nsew power input
rlabel locali s 298660 57429 298799 57647 6 VPWR
port 613 nsew power input
rlabel locali s 298660 57647 298816 57681 6 VPWR
port 613 nsew power input
rlabel locali s 298660 57681 298799 57899 6 VPWR
port 613 nsew power input
rlabel locali s 298660 57899 298661 58007 6 VPWR
port 613 nsew power input
rlabel locali s 1259 57321 1340 57429 6 VPWR
port 613 nsew power input
rlabel locali s 1121 57429 1340 57647 6 VPWR
port 613 nsew power input
rlabel locali s 1104 57647 1340 57681 6 VPWR
port 613 nsew power input
rlabel locali s 1121 57681 1340 57899 6 VPWR
port 613 nsew power input
rlabel locali s 1259 57899 1340 58007 6 VPWR
port 613 nsew power input
rlabel locali s 298660 58409 298661 58517 6 VPWR
port 613 nsew power input
rlabel locali s 298660 58517 298799 58735 6 VPWR
port 613 nsew power input
rlabel locali s 298660 58735 298816 58769 6 VPWR
port 613 nsew power input
rlabel locali s 298660 58769 298799 58987 6 VPWR
port 613 nsew power input
rlabel locali s 298660 58987 298661 59095 6 VPWR
port 613 nsew power input
rlabel locali s 1259 58409 1340 58517 6 VPWR
port 613 nsew power input
rlabel locali s 1121 58517 1340 58735 6 VPWR
port 613 nsew power input
rlabel locali s 1104 58735 1340 58769 6 VPWR
port 613 nsew power input
rlabel locali s 1121 58769 1340 58987 6 VPWR
port 613 nsew power input
rlabel locali s 1259 58987 1340 59095 6 VPWR
port 613 nsew power input
rlabel locali s 298660 59497 298661 59605 6 VPWR
port 613 nsew power input
rlabel locali s 298660 59605 298799 59823 6 VPWR
port 613 nsew power input
rlabel locali s 298660 59823 298816 59857 6 VPWR
port 613 nsew power input
rlabel locali s 298660 59857 298799 60075 6 VPWR
port 613 nsew power input
rlabel locali s 298660 60075 298661 60183 6 VPWR
port 613 nsew power input
rlabel locali s 1259 59497 1340 59605 6 VPWR
port 613 nsew power input
rlabel locali s 1121 59605 1340 59823 6 VPWR
port 613 nsew power input
rlabel locali s 1104 59823 1340 59857 6 VPWR
port 613 nsew power input
rlabel locali s 1121 59857 1340 60075 6 VPWR
port 613 nsew power input
rlabel locali s 1259 60075 1340 60183 6 VPWR
port 613 nsew power input
rlabel locali s 298660 60585 298661 60693 6 VPWR
port 613 nsew power input
rlabel locali s 298660 60693 298799 60911 6 VPWR
port 613 nsew power input
rlabel locali s 298660 60911 298816 60945 6 VPWR
port 613 nsew power input
rlabel locali s 298660 60945 298799 61163 6 VPWR
port 613 nsew power input
rlabel locali s 298660 61163 298661 61271 6 VPWR
port 613 nsew power input
rlabel locali s 1259 60585 1340 60693 6 VPWR
port 613 nsew power input
rlabel locali s 1121 60693 1340 60911 6 VPWR
port 613 nsew power input
rlabel locali s 1104 60911 1340 60945 6 VPWR
port 613 nsew power input
rlabel locali s 1121 60945 1340 61163 6 VPWR
port 613 nsew power input
rlabel locali s 1259 61163 1340 61271 6 VPWR
port 613 nsew power input
rlabel locali s 298660 61673 298661 61781 6 VPWR
port 613 nsew power input
rlabel locali s 298660 61781 298799 61999 6 VPWR
port 613 nsew power input
rlabel locali s 298660 61999 298816 62033 6 VPWR
port 613 nsew power input
rlabel locali s 298660 62033 298799 62251 6 VPWR
port 613 nsew power input
rlabel locali s 298660 62251 298661 62359 6 VPWR
port 613 nsew power input
rlabel locali s 1259 61673 1340 61781 6 VPWR
port 613 nsew power input
rlabel locali s 1121 61781 1340 61999 6 VPWR
port 613 nsew power input
rlabel locali s 1104 61999 1340 62033 6 VPWR
port 613 nsew power input
rlabel locali s 1121 62033 1340 62251 6 VPWR
port 613 nsew power input
rlabel locali s 1259 62251 1340 62359 6 VPWR
port 613 nsew power input
rlabel locali s 298660 62761 298661 62869 6 VPWR
port 613 nsew power input
rlabel locali s 298660 62869 298799 63087 6 VPWR
port 613 nsew power input
rlabel locali s 298660 63087 298816 63121 6 VPWR
port 613 nsew power input
rlabel locali s 298660 63121 298799 63339 6 VPWR
port 613 nsew power input
rlabel locali s 298660 63339 298661 63447 6 VPWR
port 613 nsew power input
rlabel locali s 1259 62761 1340 62869 6 VPWR
port 613 nsew power input
rlabel locali s 1121 62869 1340 63087 6 VPWR
port 613 nsew power input
rlabel locali s 1104 63087 1340 63121 6 VPWR
port 613 nsew power input
rlabel locali s 1121 63121 1340 63339 6 VPWR
port 613 nsew power input
rlabel locali s 1259 63339 1340 63447 6 VPWR
port 613 nsew power input
rlabel locali s 298660 63849 298661 63957 6 VPWR
port 613 nsew power input
rlabel locali s 298660 63957 298799 64175 6 VPWR
port 613 nsew power input
rlabel locali s 298660 64175 298816 64209 6 VPWR
port 613 nsew power input
rlabel locali s 298660 64209 298799 64427 6 VPWR
port 613 nsew power input
rlabel locali s 298660 64427 298661 64535 6 VPWR
port 613 nsew power input
rlabel locali s 1259 63849 1340 63957 6 VPWR
port 613 nsew power input
rlabel locali s 1121 63957 1340 64175 6 VPWR
port 613 nsew power input
rlabel locali s 1104 64175 1340 64209 6 VPWR
port 613 nsew power input
rlabel locali s 1121 64209 1340 64427 6 VPWR
port 613 nsew power input
rlabel locali s 1259 64427 1340 64535 6 VPWR
port 613 nsew power input
rlabel locali s 298660 64937 298661 65045 6 VPWR
port 613 nsew power input
rlabel locali s 298660 65045 298799 65263 6 VPWR
port 613 nsew power input
rlabel locali s 298660 65263 298816 65297 6 VPWR
port 613 nsew power input
rlabel locali s 298660 65297 298799 65515 6 VPWR
port 613 nsew power input
rlabel locali s 298660 65515 298661 65623 6 VPWR
port 613 nsew power input
rlabel locali s 1259 64937 1340 65045 6 VPWR
port 613 nsew power input
rlabel locali s 1121 65045 1340 65263 6 VPWR
port 613 nsew power input
rlabel locali s 1104 65263 1340 65297 6 VPWR
port 613 nsew power input
rlabel locali s 1121 65297 1340 65515 6 VPWR
port 613 nsew power input
rlabel locali s 1259 65515 1340 65623 6 VPWR
port 613 nsew power input
rlabel locali s 298660 66025 298661 66133 6 VPWR
port 613 nsew power input
rlabel locali s 298660 66133 298799 66351 6 VPWR
port 613 nsew power input
rlabel locali s 298660 66351 298816 66385 6 VPWR
port 613 nsew power input
rlabel locali s 298660 66385 298799 66603 6 VPWR
port 613 nsew power input
rlabel locali s 298660 66603 298661 66711 6 VPWR
port 613 nsew power input
rlabel locali s 1259 66025 1340 66133 6 VPWR
port 613 nsew power input
rlabel locali s 1121 66133 1340 66351 6 VPWR
port 613 nsew power input
rlabel locali s 1104 66351 1340 66385 6 VPWR
port 613 nsew power input
rlabel locali s 1121 66385 1340 66603 6 VPWR
port 613 nsew power input
rlabel locali s 1259 66603 1340 66711 6 VPWR
port 613 nsew power input
rlabel locali s 298660 67113 298661 67221 6 VPWR
port 613 nsew power input
rlabel locali s 298660 67221 298799 67439 6 VPWR
port 613 nsew power input
rlabel locali s 298660 67439 298816 67473 6 VPWR
port 613 nsew power input
rlabel locali s 298660 67473 298799 67691 6 VPWR
port 613 nsew power input
rlabel locali s 298660 67691 298661 67799 6 VPWR
port 613 nsew power input
rlabel locali s 1259 67113 1340 67221 6 VPWR
port 613 nsew power input
rlabel locali s 1121 67221 1340 67439 6 VPWR
port 613 nsew power input
rlabel locali s 1104 67439 1340 67473 6 VPWR
port 613 nsew power input
rlabel locali s 1121 67473 1340 67691 6 VPWR
port 613 nsew power input
rlabel locali s 1259 67691 1340 67799 6 VPWR
port 613 nsew power input
rlabel locali s 298660 68201 298661 68309 6 VPWR
port 613 nsew power input
rlabel locali s 298660 68309 298799 68527 6 VPWR
port 613 nsew power input
rlabel locali s 298660 68527 298816 68561 6 VPWR
port 613 nsew power input
rlabel locali s 298660 68561 298799 68779 6 VPWR
port 613 nsew power input
rlabel locali s 298660 68779 298661 68887 6 VPWR
port 613 nsew power input
rlabel locali s 1259 68201 1340 68309 6 VPWR
port 613 nsew power input
rlabel locali s 1121 68309 1340 68527 6 VPWR
port 613 nsew power input
rlabel locali s 1104 68527 1340 68561 6 VPWR
port 613 nsew power input
rlabel locali s 1121 68561 1340 68779 6 VPWR
port 613 nsew power input
rlabel locali s 1259 68779 1340 68887 6 VPWR
port 613 nsew power input
rlabel locali s 298660 69289 298661 69397 6 VPWR
port 613 nsew power input
rlabel locali s 298660 69397 298799 69615 6 VPWR
port 613 nsew power input
rlabel locali s 298660 69615 298816 69649 6 VPWR
port 613 nsew power input
rlabel locali s 298660 69649 298799 69867 6 VPWR
port 613 nsew power input
rlabel locali s 298660 69867 298661 69975 6 VPWR
port 613 nsew power input
rlabel locali s 1259 69289 1340 69397 6 VPWR
port 613 nsew power input
rlabel locali s 1121 69397 1340 69615 6 VPWR
port 613 nsew power input
rlabel locali s 1104 69615 1340 69649 6 VPWR
port 613 nsew power input
rlabel locali s 1121 69649 1340 69867 6 VPWR
port 613 nsew power input
rlabel locali s 1259 69867 1340 69975 6 VPWR
port 613 nsew power input
rlabel locali s 298660 70377 298661 70485 6 VPWR
port 613 nsew power input
rlabel locali s 298660 70485 298799 70703 6 VPWR
port 613 nsew power input
rlabel locali s 298660 70703 298816 70737 6 VPWR
port 613 nsew power input
rlabel locali s 298660 70737 298799 70955 6 VPWR
port 613 nsew power input
rlabel locali s 298660 70955 298661 71063 6 VPWR
port 613 nsew power input
rlabel locali s 1259 70377 1340 70485 6 VPWR
port 613 nsew power input
rlabel locali s 1121 70485 1340 70703 6 VPWR
port 613 nsew power input
rlabel locali s 1104 70703 1340 70737 6 VPWR
port 613 nsew power input
rlabel locali s 1121 70737 1340 70955 6 VPWR
port 613 nsew power input
rlabel locali s 1259 70955 1340 71063 6 VPWR
port 613 nsew power input
rlabel locali s 298660 71465 298661 71573 6 VPWR
port 613 nsew power input
rlabel locali s 298660 71573 298799 71791 6 VPWR
port 613 nsew power input
rlabel locali s 298660 71791 298816 71825 6 VPWR
port 613 nsew power input
rlabel locali s 298660 71825 298799 72043 6 VPWR
port 613 nsew power input
rlabel locali s 298660 72043 298661 72151 6 VPWR
port 613 nsew power input
rlabel locali s 1259 71465 1340 71573 6 VPWR
port 613 nsew power input
rlabel locali s 1121 71573 1340 71791 6 VPWR
port 613 nsew power input
rlabel locali s 1104 71791 1340 71825 6 VPWR
port 613 nsew power input
rlabel locali s 1121 71825 1340 72043 6 VPWR
port 613 nsew power input
rlabel locali s 1259 72043 1340 72151 6 VPWR
port 613 nsew power input
rlabel locali s 298660 72553 298661 72661 6 VPWR
port 613 nsew power input
rlabel locali s 298660 72661 298799 72879 6 VPWR
port 613 nsew power input
rlabel locali s 298660 72879 298816 72913 6 VPWR
port 613 nsew power input
rlabel locali s 298660 72913 298799 73131 6 VPWR
port 613 nsew power input
rlabel locali s 298660 73131 298661 73239 6 VPWR
port 613 nsew power input
rlabel locali s 1259 72553 1340 72661 6 VPWR
port 613 nsew power input
rlabel locali s 1121 72661 1340 72879 6 VPWR
port 613 nsew power input
rlabel locali s 1104 72879 1340 72913 6 VPWR
port 613 nsew power input
rlabel locali s 1121 72913 1340 73131 6 VPWR
port 613 nsew power input
rlabel locali s 1259 73131 1340 73239 6 VPWR
port 613 nsew power input
rlabel locali s 298660 73641 298661 73749 6 VPWR
port 613 nsew power input
rlabel locali s 298660 73749 298799 73967 6 VPWR
port 613 nsew power input
rlabel locali s 298660 73967 298816 74001 6 VPWR
port 613 nsew power input
rlabel locali s 298660 74001 298799 74219 6 VPWR
port 613 nsew power input
rlabel locali s 298660 74219 298661 74327 6 VPWR
port 613 nsew power input
rlabel locali s 1259 73641 1340 73749 6 VPWR
port 613 nsew power input
rlabel locali s 1121 73749 1340 73967 6 VPWR
port 613 nsew power input
rlabel locali s 1104 73967 1340 74001 6 VPWR
port 613 nsew power input
rlabel locali s 1121 74001 1340 74219 6 VPWR
port 613 nsew power input
rlabel locali s 1259 74219 1340 74327 6 VPWR
port 613 nsew power input
rlabel locali s 298660 74729 298661 74837 6 VPWR
port 613 nsew power input
rlabel locali s 298660 74837 298799 75055 6 VPWR
port 613 nsew power input
rlabel locali s 298660 75055 298816 75089 6 VPWR
port 613 nsew power input
rlabel locali s 298660 75089 298799 75307 6 VPWR
port 613 nsew power input
rlabel locali s 298660 75307 298661 75415 6 VPWR
port 613 nsew power input
rlabel locali s 1259 74729 1340 74837 6 VPWR
port 613 nsew power input
rlabel locali s 1121 74837 1340 75055 6 VPWR
port 613 nsew power input
rlabel locali s 1104 75055 1340 75089 6 VPWR
port 613 nsew power input
rlabel locali s 1121 75089 1340 75307 6 VPWR
port 613 nsew power input
rlabel locali s 1259 75307 1340 75415 6 VPWR
port 613 nsew power input
rlabel locali s 298660 75817 298661 75925 6 VPWR
port 613 nsew power input
rlabel locali s 298660 75925 298799 76143 6 VPWR
port 613 nsew power input
rlabel locali s 298660 76143 298816 76177 6 VPWR
port 613 nsew power input
rlabel locali s 298660 76177 298799 76395 6 VPWR
port 613 nsew power input
rlabel locali s 298660 76395 298661 76503 6 VPWR
port 613 nsew power input
rlabel locali s 1259 75817 1340 75925 6 VPWR
port 613 nsew power input
rlabel locali s 1121 75925 1340 76143 6 VPWR
port 613 nsew power input
rlabel locali s 1104 76143 1340 76177 6 VPWR
port 613 nsew power input
rlabel locali s 1121 76177 1340 76395 6 VPWR
port 613 nsew power input
rlabel locali s 1259 76395 1340 76503 6 VPWR
port 613 nsew power input
rlabel locali s 298660 76905 298661 77013 6 VPWR
port 613 nsew power input
rlabel locali s 298660 77013 298799 77231 6 VPWR
port 613 nsew power input
rlabel locali s 298660 77231 298816 77265 6 VPWR
port 613 nsew power input
rlabel locali s 298660 77265 298799 77483 6 VPWR
port 613 nsew power input
rlabel locali s 298660 77483 298661 77591 6 VPWR
port 613 nsew power input
rlabel locali s 1259 76905 1340 77013 6 VPWR
port 613 nsew power input
rlabel locali s 1121 77013 1340 77231 6 VPWR
port 613 nsew power input
rlabel locali s 1104 77231 1340 77265 6 VPWR
port 613 nsew power input
rlabel locali s 1121 77265 1340 77483 6 VPWR
port 613 nsew power input
rlabel locali s 1259 77483 1340 77591 6 VPWR
port 613 nsew power input
rlabel locali s 298660 77993 298661 78101 6 VPWR
port 613 nsew power input
rlabel locali s 298660 78101 298799 78319 6 VPWR
port 613 nsew power input
rlabel locali s 298660 78319 298816 78353 6 VPWR
port 613 nsew power input
rlabel locali s 298660 78353 298799 78571 6 VPWR
port 613 nsew power input
rlabel locali s 298660 78571 298661 78679 6 VPWR
port 613 nsew power input
rlabel locali s 1259 77993 1340 78101 6 VPWR
port 613 nsew power input
rlabel locali s 1121 78101 1340 78319 6 VPWR
port 613 nsew power input
rlabel locali s 1104 78319 1340 78353 6 VPWR
port 613 nsew power input
rlabel locali s 1121 78353 1340 78571 6 VPWR
port 613 nsew power input
rlabel locali s 1259 78571 1340 78679 6 VPWR
port 613 nsew power input
rlabel locali s 298660 79081 298661 79189 6 VPWR
port 613 nsew power input
rlabel locali s 298660 79189 298799 79407 6 VPWR
port 613 nsew power input
rlabel locali s 298660 79407 298816 79441 6 VPWR
port 613 nsew power input
rlabel locali s 298660 79441 298799 79659 6 VPWR
port 613 nsew power input
rlabel locali s 298660 79659 298661 79767 6 VPWR
port 613 nsew power input
rlabel locali s 1259 79081 1340 79189 6 VPWR
port 613 nsew power input
rlabel locali s 1121 79189 1340 79407 6 VPWR
port 613 nsew power input
rlabel locali s 1104 79407 1340 79441 6 VPWR
port 613 nsew power input
rlabel locali s 1121 79441 1340 79659 6 VPWR
port 613 nsew power input
rlabel locali s 1259 79659 1340 79767 6 VPWR
port 613 nsew power input
rlabel locali s 298660 80169 298661 80277 6 VPWR
port 613 nsew power input
rlabel locali s 298660 80277 298799 80495 6 VPWR
port 613 nsew power input
rlabel locali s 298660 80495 298816 80529 6 VPWR
port 613 nsew power input
rlabel locali s 298660 80529 298799 80747 6 VPWR
port 613 nsew power input
rlabel locali s 298660 80747 298661 80855 6 VPWR
port 613 nsew power input
rlabel locali s 1259 80169 1340 80277 6 VPWR
port 613 nsew power input
rlabel locali s 1121 80277 1340 80495 6 VPWR
port 613 nsew power input
rlabel locali s 1104 80495 1340 80529 6 VPWR
port 613 nsew power input
rlabel locali s 1121 80529 1340 80747 6 VPWR
port 613 nsew power input
rlabel locali s 1259 80747 1340 80855 6 VPWR
port 613 nsew power input
rlabel locali s 298660 81257 298661 81365 6 VPWR
port 613 nsew power input
rlabel locali s 298660 81365 298799 81583 6 VPWR
port 613 nsew power input
rlabel locali s 298660 81583 298816 81617 6 VPWR
port 613 nsew power input
rlabel locali s 298660 81617 298799 81835 6 VPWR
port 613 nsew power input
rlabel locali s 298660 81835 298661 81943 6 VPWR
port 613 nsew power input
rlabel locali s 1259 81257 1340 81365 6 VPWR
port 613 nsew power input
rlabel locali s 1121 81365 1340 81583 6 VPWR
port 613 nsew power input
rlabel locali s 1104 81583 1340 81617 6 VPWR
port 613 nsew power input
rlabel locali s 1121 81617 1340 81835 6 VPWR
port 613 nsew power input
rlabel locali s 1259 81835 1340 81943 6 VPWR
port 613 nsew power input
rlabel locali s 298660 82345 298661 82453 6 VPWR
port 613 nsew power input
rlabel locali s 298660 82453 298799 82671 6 VPWR
port 613 nsew power input
rlabel locali s 298660 82671 298816 82705 6 VPWR
port 613 nsew power input
rlabel locali s 298660 82705 298799 82923 6 VPWR
port 613 nsew power input
rlabel locali s 298660 82923 298661 83031 6 VPWR
port 613 nsew power input
rlabel locali s 1259 82345 1340 82453 6 VPWR
port 613 nsew power input
rlabel locali s 1121 82453 1340 82671 6 VPWR
port 613 nsew power input
rlabel locali s 1104 82671 1340 82705 6 VPWR
port 613 nsew power input
rlabel locali s 1121 82705 1340 82923 6 VPWR
port 613 nsew power input
rlabel locali s 1259 82923 1340 83031 6 VPWR
port 613 nsew power input
rlabel locali s 298660 83433 298661 83541 6 VPWR
port 613 nsew power input
rlabel locali s 298660 83541 298799 83759 6 VPWR
port 613 nsew power input
rlabel locali s 298660 83759 298816 83793 6 VPWR
port 613 nsew power input
rlabel locali s 298660 83793 298799 84011 6 VPWR
port 613 nsew power input
rlabel locali s 298660 84011 298661 84119 6 VPWR
port 613 nsew power input
rlabel locali s 1259 83433 1340 83541 6 VPWR
port 613 nsew power input
rlabel locali s 1121 83541 1340 83759 6 VPWR
port 613 nsew power input
rlabel locali s 1104 83759 1340 83793 6 VPWR
port 613 nsew power input
rlabel locali s 1121 83793 1340 84011 6 VPWR
port 613 nsew power input
rlabel locali s 1259 84011 1340 84119 6 VPWR
port 613 nsew power input
rlabel locali s 298660 84521 298661 84629 6 VPWR
port 613 nsew power input
rlabel locali s 298660 84629 298799 84847 6 VPWR
port 613 nsew power input
rlabel locali s 298660 84847 298816 84881 6 VPWR
port 613 nsew power input
rlabel locali s 298660 84881 298799 85099 6 VPWR
port 613 nsew power input
rlabel locali s 298660 85099 298661 85207 6 VPWR
port 613 nsew power input
rlabel locali s 1259 84521 1340 84629 6 VPWR
port 613 nsew power input
rlabel locali s 1121 84629 1340 84847 6 VPWR
port 613 nsew power input
rlabel locali s 1104 84847 1340 84881 6 VPWR
port 613 nsew power input
rlabel locali s 1121 84881 1340 85099 6 VPWR
port 613 nsew power input
rlabel locali s 1259 85099 1340 85207 6 VPWR
port 613 nsew power input
rlabel locali s 298660 85609 298661 85717 6 VPWR
port 613 nsew power input
rlabel locali s 298660 85717 298799 85935 6 VPWR
port 613 nsew power input
rlabel locali s 298660 85935 298816 85969 6 VPWR
port 613 nsew power input
rlabel locali s 298660 85969 298799 86187 6 VPWR
port 613 nsew power input
rlabel locali s 298660 86187 298661 86295 6 VPWR
port 613 nsew power input
rlabel locali s 1259 85609 1340 85717 6 VPWR
port 613 nsew power input
rlabel locali s 1121 85717 1340 85935 6 VPWR
port 613 nsew power input
rlabel locali s 1104 85935 1340 85969 6 VPWR
port 613 nsew power input
rlabel locali s 1121 85969 1340 86187 6 VPWR
port 613 nsew power input
rlabel locali s 1259 86187 1340 86295 6 VPWR
port 613 nsew power input
rlabel locali s 298660 86697 298661 86805 6 VPWR
port 613 nsew power input
rlabel locali s 298660 86805 298799 87023 6 VPWR
port 613 nsew power input
rlabel locali s 298660 87023 298816 87057 6 VPWR
port 613 nsew power input
rlabel locali s 298660 87057 298799 87275 6 VPWR
port 613 nsew power input
rlabel locali s 298660 87275 298661 87383 6 VPWR
port 613 nsew power input
rlabel locali s 1259 86697 1340 86805 6 VPWR
port 613 nsew power input
rlabel locali s 1121 86805 1340 87023 6 VPWR
port 613 nsew power input
rlabel locali s 1104 87023 1340 87057 6 VPWR
port 613 nsew power input
rlabel locali s 1121 87057 1340 87275 6 VPWR
port 613 nsew power input
rlabel locali s 1259 87275 1340 87383 6 VPWR
port 613 nsew power input
rlabel locali s 298660 87785 298661 87893 6 VPWR
port 613 nsew power input
rlabel locali s 298660 87893 298799 88111 6 VPWR
port 613 nsew power input
rlabel locali s 298660 88111 298816 88145 6 VPWR
port 613 nsew power input
rlabel locali s 298660 88145 298799 88363 6 VPWR
port 613 nsew power input
rlabel locali s 298660 88363 298661 88471 6 VPWR
port 613 nsew power input
rlabel locali s 1259 87785 1340 87893 6 VPWR
port 613 nsew power input
rlabel locali s 1121 87893 1340 88111 6 VPWR
port 613 nsew power input
rlabel locali s 1104 88111 1340 88145 6 VPWR
port 613 nsew power input
rlabel locali s 1121 88145 1340 88363 6 VPWR
port 613 nsew power input
rlabel locali s 1259 88363 1340 88471 6 VPWR
port 613 nsew power input
rlabel locali s 298660 88873 298661 88981 6 VPWR
port 613 nsew power input
rlabel locali s 298660 88981 298799 89199 6 VPWR
port 613 nsew power input
rlabel locali s 298660 89199 298816 89233 6 VPWR
port 613 nsew power input
rlabel locali s 298660 89233 298799 89451 6 VPWR
port 613 nsew power input
rlabel locali s 298660 89451 298661 89559 6 VPWR
port 613 nsew power input
rlabel locali s 1259 88873 1340 88981 6 VPWR
port 613 nsew power input
rlabel locali s 1121 88981 1340 89199 6 VPWR
port 613 nsew power input
rlabel locali s 1104 89199 1340 89233 6 VPWR
port 613 nsew power input
rlabel locali s 1121 89233 1340 89451 6 VPWR
port 613 nsew power input
rlabel locali s 1259 89451 1340 89559 6 VPWR
port 613 nsew power input
rlabel locali s 298660 89961 298661 90069 6 VPWR
port 613 nsew power input
rlabel locali s 298660 90069 298799 90287 6 VPWR
port 613 nsew power input
rlabel locali s 298660 90287 298816 90321 6 VPWR
port 613 nsew power input
rlabel locali s 298660 90321 298799 90539 6 VPWR
port 613 nsew power input
rlabel locali s 298660 90539 298661 90647 6 VPWR
port 613 nsew power input
rlabel locali s 1259 89961 1340 90069 6 VPWR
port 613 nsew power input
rlabel locali s 1121 90069 1340 90287 6 VPWR
port 613 nsew power input
rlabel locali s 1104 90287 1340 90321 6 VPWR
port 613 nsew power input
rlabel locali s 1121 90321 1340 90539 6 VPWR
port 613 nsew power input
rlabel locali s 1259 90539 1340 90647 6 VPWR
port 613 nsew power input
rlabel locali s 298660 91049 298661 91157 6 VPWR
port 613 nsew power input
rlabel locali s 298660 91157 298799 91375 6 VPWR
port 613 nsew power input
rlabel locali s 298660 91375 298816 91409 6 VPWR
port 613 nsew power input
rlabel locali s 298660 91409 298799 91627 6 VPWR
port 613 nsew power input
rlabel locali s 298660 91627 298661 91735 6 VPWR
port 613 nsew power input
rlabel locali s 1259 91049 1340 91157 6 VPWR
port 613 nsew power input
rlabel locali s 1121 91157 1340 91375 6 VPWR
port 613 nsew power input
rlabel locali s 1104 91375 1340 91409 6 VPWR
port 613 nsew power input
rlabel locali s 1121 91409 1340 91627 6 VPWR
port 613 nsew power input
rlabel locali s 1259 91627 1340 91735 6 VPWR
port 613 nsew power input
rlabel locali s 298660 92137 298661 92245 6 VPWR
port 613 nsew power input
rlabel locali s 298660 92245 298799 92463 6 VPWR
port 613 nsew power input
rlabel locali s 298660 92463 298816 92497 6 VPWR
port 613 nsew power input
rlabel locali s 298660 92497 298799 92715 6 VPWR
port 613 nsew power input
rlabel locali s 298660 92715 298661 92823 6 VPWR
port 613 nsew power input
rlabel locali s 1259 92137 1340 92245 6 VPWR
port 613 nsew power input
rlabel locali s 1121 92245 1340 92463 6 VPWR
port 613 nsew power input
rlabel locali s 1104 92463 1340 92497 6 VPWR
port 613 nsew power input
rlabel locali s 1121 92497 1340 92715 6 VPWR
port 613 nsew power input
rlabel locali s 1259 92715 1340 92823 6 VPWR
port 613 nsew power input
rlabel locali s 298660 93225 298661 93333 6 VPWR
port 613 nsew power input
rlabel locali s 298660 93333 298799 93551 6 VPWR
port 613 nsew power input
rlabel locali s 298660 93551 298816 93585 6 VPWR
port 613 nsew power input
rlabel locali s 298660 93585 298799 93803 6 VPWR
port 613 nsew power input
rlabel locali s 298660 93803 298661 93911 6 VPWR
port 613 nsew power input
rlabel locali s 1259 93225 1340 93333 6 VPWR
port 613 nsew power input
rlabel locali s 1121 93333 1340 93551 6 VPWR
port 613 nsew power input
rlabel locali s 1104 93551 1340 93585 6 VPWR
port 613 nsew power input
rlabel locali s 1121 93585 1340 93803 6 VPWR
port 613 nsew power input
rlabel locali s 1259 93803 1340 93911 6 VPWR
port 613 nsew power input
rlabel locali s 298660 94313 298661 94421 6 VPWR
port 613 nsew power input
rlabel locali s 298660 94421 298799 94639 6 VPWR
port 613 nsew power input
rlabel locali s 298660 94639 298816 94673 6 VPWR
port 613 nsew power input
rlabel locali s 298660 94673 298799 94891 6 VPWR
port 613 nsew power input
rlabel locali s 298660 94891 298661 94999 6 VPWR
port 613 nsew power input
rlabel locali s 1259 94313 1340 94421 6 VPWR
port 613 nsew power input
rlabel locali s 1121 94421 1340 94639 6 VPWR
port 613 nsew power input
rlabel locali s 1104 94639 1340 94673 6 VPWR
port 613 nsew power input
rlabel locali s 1121 94673 1340 94891 6 VPWR
port 613 nsew power input
rlabel locali s 1259 94891 1340 94999 6 VPWR
port 613 nsew power input
rlabel locali s 298660 95401 298661 95509 6 VPWR
port 613 nsew power input
rlabel locali s 298660 95509 298799 95727 6 VPWR
port 613 nsew power input
rlabel locali s 298660 95727 298816 95761 6 VPWR
port 613 nsew power input
rlabel locali s 298660 95761 298799 95979 6 VPWR
port 613 nsew power input
rlabel locali s 298660 95979 298661 96087 6 VPWR
port 613 nsew power input
rlabel locali s 1259 95401 1340 95509 6 VPWR
port 613 nsew power input
rlabel locali s 1121 95509 1340 95727 6 VPWR
port 613 nsew power input
rlabel locali s 1104 95727 1340 95761 6 VPWR
port 613 nsew power input
rlabel locali s 1121 95761 1340 95979 6 VPWR
port 613 nsew power input
rlabel locali s 1259 95979 1340 96087 6 VPWR
port 613 nsew power input
rlabel locali s 298660 96489 298661 96597 6 VPWR
port 613 nsew power input
rlabel locali s 298660 96597 298799 96815 6 VPWR
port 613 nsew power input
rlabel locali s 298660 96815 298816 96849 6 VPWR
port 613 nsew power input
rlabel locali s 298660 96849 298799 97067 6 VPWR
port 613 nsew power input
rlabel locali s 298660 97067 298661 97175 6 VPWR
port 613 nsew power input
rlabel locali s 1259 96489 1340 96597 6 VPWR
port 613 nsew power input
rlabel locali s 1121 96597 1340 96815 6 VPWR
port 613 nsew power input
rlabel locali s 1104 96815 1340 96849 6 VPWR
port 613 nsew power input
rlabel locali s 1121 96849 1340 97067 6 VPWR
port 613 nsew power input
rlabel locali s 1259 97067 1340 97175 6 VPWR
port 613 nsew power input
rlabel locali s 298660 97577 298661 97685 6 VPWR
port 613 nsew power input
rlabel locali s 298660 97685 298799 97903 6 VPWR
port 613 nsew power input
rlabel locali s 298660 97903 298816 97937 6 VPWR
port 613 nsew power input
rlabel locali s 298660 97937 298799 98155 6 VPWR
port 613 nsew power input
rlabel locali s 298660 98155 298661 98263 6 VPWR
port 613 nsew power input
rlabel locali s 1259 97577 1340 97685 6 VPWR
port 613 nsew power input
rlabel locali s 1121 97685 1340 97903 6 VPWR
port 613 nsew power input
rlabel locali s 1104 97903 1340 97937 6 VPWR
port 613 nsew power input
rlabel locali s 1121 97937 1340 98155 6 VPWR
port 613 nsew power input
rlabel locali s 1259 98155 1340 98263 6 VPWR
port 613 nsew power input
rlabel locali s 298660 98665 298661 98773 6 VPWR
port 613 nsew power input
rlabel locali s 298660 98773 298799 98991 6 VPWR
port 613 nsew power input
rlabel locali s 298660 98991 298816 99025 6 VPWR
port 613 nsew power input
rlabel locali s 298660 99025 298799 99243 6 VPWR
port 613 nsew power input
rlabel locali s 298660 99243 298661 99351 6 VPWR
port 613 nsew power input
rlabel locali s 1259 98665 1340 98773 6 VPWR
port 613 nsew power input
rlabel locali s 1121 98773 1340 98991 6 VPWR
port 613 nsew power input
rlabel locali s 1104 98991 1340 99025 6 VPWR
port 613 nsew power input
rlabel locali s 1121 99025 1340 99243 6 VPWR
port 613 nsew power input
rlabel locali s 1259 99243 1340 99351 6 VPWR
port 613 nsew power input
rlabel locali s 298660 99753 298661 99861 6 VPWR
port 613 nsew power input
rlabel locali s 298660 99861 298799 100079 6 VPWR
port 613 nsew power input
rlabel locali s 298660 100079 298816 100113 6 VPWR
port 613 nsew power input
rlabel locali s 298660 100113 298799 100331 6 VPWR
port 613 nsew power input
rlabel locali s 298660 100331 298661 100439 6 VPWR
port 613 nsew power input
rlabel locali s 1259 99753 1340 99861 6 VPWR
port 613 nsew power input
rlabel locali s 1121 99861 1340 100079 6 VPWR
port 613 nsew power input
rlabel locali s 1104 100079 1340 100113 6 VPWR
port 613 nsew power input
rlabel locali s 1121 100113 1340 100331 6 VPWR
port 613 nsew power input
rlabel locali s 1259 100331 1340 100439 6 VPWR
port 613 nsew power input
rlabel locali s 298660 100841 298661 100949 6 VPWR
port 613 nsew power input
rlabel locali s 298660 100949 298799 101167 6 VPWR
port 613 nsew power input
rlabel locali s 298660 101167 298816 101201 6 VPWR
port 613 nsew power input
rlabel locali s 298660 101201 298799 101419 6 VPWR
port 613 nsew power input
rlabel locali s 298660 101419 298661 101527 6 VPWR
port 613 nsew power input
rlabel locali s 1259 100841 1340 100949 6 VPWR
port 613 nsew power input
rlabel locali s 1121 100949 1340 101167 6 VPWR
port 613 nsew power input
rlabel locali s 1104 101167 1340 101201 6 VPWR
port 613 nsew power input
rlabel locali s 1121 101201 1340 101419 6 VPWR
port 613 nsew power input
rlabel locali s 1259 101419 1340 101527 6 VPWR
port 613 nsew power input
rlabel locali s 298660 101929 298661 102037 6 VPWR
port 613 nsew power input
rlabel locali s 298660 102037 298799 102255 6 VPWR
port 613 nsew power input
rlabel locali s 298660 102255 298816 102289 6 VPWR
port 613 nsew power input
rlabel locali s 298660 102289 298799 102507 6 VPWR
port 613 nsew power input
rlabel locali s 298660 102507 298661 102615 6 VPWR
port 613 nsew power input
rlabel locali s 1259 101929 1340 102037 6 VPWR
port 613 nsew power input
rlabel locali s 1121 102037 1340 102255 6 VPWR
port 613 nsew power input
rlabel locali s 1104 102255 1340 102289 6 VPWR
port 613 nsew power input
rlabel locali s 1121 102289 1340 102507 6 VPWR
port 613 nsew power input
rlabel locali s 1259 102507 1340 102615 6 VPWR
port 613 nsew power input
rlabel locali s 298660 103017 298661 103125 6 VPWR
port 613 nsew power input
rlabel locali s 298660 103125 298799 103343 6 VPWR
port 613 nsew power input
rlabel locali s 298660 103343 298816 103377 6 VPWR
port 613 nsew power input
rlabel locali s 298660 103377 298799 103595 6 VPWR
port 613 nsew power input
rlabel locali s 298660 103595 298661 103703 6 VPWR
port 613 nsew power input
rlabel locali s 1259 103017 1340 103125 6 VPWR
port 613 nsew power input
rlabel locali s 1121 103125 1340 103343 6 VPWR
port 613 nsew power input
rlabel locali s 1104 103343 1340 103377 6 VPWR
port 613 nsew power input
rlabel locali s 1121 103377 1340 103595 6 VPWR
port 613 nsew power input
rlabel locali s 1259 103595 1340 103703 6 VPWR
port 613 nsew power input
rlabel locali s 298660 104105 298661 104213 6 VPWR
port 613 nsew power input
rlabel locali s 298660 104213 298799 104431 6 VPWR
port 613 nsew power input
rlabel locali s 298660 104431 298816 104465 6 VPWR
port 613 nsew power input
rlabel locali s 298660 104465 298799 104683 6 VPWR
port 613 nsew power input
rlabel locali s 298660 104683 298661 104791 6 VPWR
port 613 nsew power input
rlabel locali s 1259 104105 1340 104213 6 VPWR
port 613 nsew power input
rlabel locali s 1121 104213 1340 104431 6 VPWR
port 613 nsew power input
rlabel locali s 1104 104431 1340 104465 6 VPWR
port 613 nsew power input
rlabel locali s 1121 104465 1340 104683 6 VPWR
port 613 nsew power input
rlabel locali s 1259 104683 1340 104791 6 VPWR
port 613 nsew power input
rlabel locali s 298660 105193 298661 105301 6 VPWR
port 613 nsew power input
rlabel locali s 298660 105301 298799 105519 6 VPWR
port 613 nsew power input
rlabel locali s 298660 105519 298816 105553 6 VPWR
port 613 nsew power input
rlabel locali s 298660 105553 298799 105771 6 VPWR
port 613 nsew power input
rlabel locali s 298660 105771 298661 105879 6 VPWR
port 613 nsew power input
rlabel locali s 1259 105193 1340 105301 6 VPWR
port 613 nsew power input
rlabel locali s 1121 105301 1340 105519 6 VPWR
port 613 nsew power input
rlabel locali s 1104 105519 1340 105553 6 VPWR
port 613 nsew power input
rlabel locali s 1121 105553 1340 105771 6 VPWR
port 613 nsew power input
rlabel locali s 1259 105771 1340 105879 6 VPWR
port 613 nsew power input
rlabel locali s 298660 106281 298661 106389 6 VPWR
port 613 nsew power input
rlabel locali s 298660 106389 298799 106607 6 VPWR
port 613 nsew power input
rlabel locali s 298660 106607 298816 106641 6 VPWR
port 613 nsew power input
rlabel locali s 298660 106641 298799 106859 6 VPWR
port 613 nsew power input
rlabel locali s 298660 106859 298661 106967 6 VPWR
port 613 nsew power input
rlabel locali s 1259 106281 1340 106389 6 VPWR
port 613 nsew power input
rlabel locali s 1121 106389 1340 106607 6 VPWR
port 613 nsew power input
rlabel locali s 1104 106607 1340 106641 6 VPWR
port 613 nsew power input
rlabel locali s 1121 106641 1340 106859 6 VPWR
port 613 nsew power input
rlabel locali s 1259 106859 1340 106967 6 VPWR
port 613 nsew power input
rlabel locali s 298660 107369 298661 107477 6 VPWR
port 613 nsew power input
rlabel locali s 298660 107477 298799 107695 6 VPWR
port 613 nsew power input
rlabel locali s 298660 107695 298816 107729 6 VPWR
port 613 nsew power input
rlabel locali s 298660 107729 298799 107947 6 VPWR
port 613 nsew power input
rlabel locali s 298660 107947 298661 108055 6 VPWR
port 613 nsew power input
rlabel locali s 1259 107369 1340 107477 6 VPWR
port 613 nsew power input
rlabel locali s 1121 107477 1340 107695 6 VPWR
port 613 nsew power input
rlabel locali s 1104 107695 1340 107729 6 VPWR
port 613 nsew power input
rlabel locali s 1121 107729 1340 107947 6 VPWR
port 613 nsew power input
rlabel locali s 1259 107947 1340 108055 6 VPWR
port 613 nsew power input
rlabel locali s 298660 108457 298661 108565 6 VPWR
port 613 nsew power input
rlabel locali s 298660 108565 298799 108783 6 VPWR
port 613 nsew power input
rlabel locali s 298660 108783 298816 108817 6 VPWR
port 613 nsew power input
rlabel locali s 298660 108817 298799 109035 6 VPWR
port 613 nsew power input
rlabel locali s 298660 109035 298661 109143 6 VPWR
port 613 nsew power input
rlabel locali s 1259 108457 1340 108565 6 VPWR
port 613 nsew power input
rlabel locali s 1121 108565 1340 108783 6 VPWR
port 613 nsew power input
rlabel locali s 1104 108783 1340 108817 6 VPWR
port 613 nsew power input
rlabel locali s 1121 108817 1340 109035 6 VPWR
port 613 nsew power input
rlabel locali s 1259 109035 1340 109143 6 VPWR
port 613 nsew power input
rlabel locali s 298660 109545 298661 109653 6 VPWR
port 613 nsew power input
rlabel locali s 298660 109653 298799 109871 6 VPWR
port 613 nsew power input
rlabel locali s 298660 109871 298816 109905 6 VPWR
port 613 nsew power input
rlabel locali s 298660 109905 298799 110123 6 VPWR
port 613 nsew power input
rlabel locali s 298660 110123 298661 110231 6 VPWR
port 613 nsew power input
rlabel locali s 1259 109545 1340 109653 6 VPWR
port 613 nsew power input
rlabel locali s 1121 109653 1340 109871 6 VPWR
port 613 nsew power input
rlabel locali s 1104 109871 1340 109905 6 VPWR
port 613 nsew power input
rlabel locali s 1121 109905 1340 110123 6 VPWR
port 613 nsew power input
rlabel locali s 1259 110123 1340 110231 6 VPWR
port 613 nsew power input
rlabel locali s 298660 110633 298661 110741 6 VPWR
port 613 nsew power input
rlabel locali s 298660 110741 298799 110959 6 VPWR
port 613 nsew power input
rlabel locali s 298660 110959 298816 110993 6 VPWR
port 613 nsew power input
rlabel locali s 298660 110993 298799 111211 6 VPWR
port 613 nsew power input
rlabel locali s 298660 111211 298661 111319 6 VPWR
port 613 nsew power input
rlabel locali s 1259 110633 1340 110741 6 VPWR
port 613 nsew power input
rlabel locali s 1121 110741 1340 110959 6 VPWR
port 613 nsew power input
rlabel locali s 1104 110959 1340 110993 6 VPWR
port 613 nsew power input
rlabel locali s 1121 110993 1340 111211 6 VPWR
port 613 nsew power input
rlabel locali s 1259 111211 1340 111319 6 VPWR
port 613 nsew power input
rlabel locali s 298660 111721 298661 111829 6 VPWR
port 613 nsew power input
rlabel locali s 298660 111829 298799 112047 6 VPWR
port 613 nsew power input
rlabel locali s 298660 112047 298816 112081 6 VPWR
port 613 nsew power input
rlabel locali s 298660 112081 298799 112299 6 VPWR
port 613 nsew power input
rlabel locali s 298660 112299 298661 112407 6 VPWR
port 613 nsew power input
rlabel locali s 1259 111721 1340 111829 6 VPWR
port 613 nsew power input
rlabel locali s 1121 111829 1340 112047 6 VPWR
port 613 nsew power input
rlabel locali s 1104 112047 1340 112081 6 VPWR
port 613 nsew power input
rlabel locali s 1121 112081 1340 112299 6 VPWR
port 613 nsew power input
rlabel locali s 1259 112299 1340 112407 6 VPWR
port 613 nsew power input
rlabel locali s 298660 112809 298661 112917 6 VPWR
port 613 nsew power input
rlabel locali s 298660 112917 298799 113135 6 VPWR
port 613 nsew power input
rlabel locali s 298660 113135 298816 113169 6 VPWR
port 613 nsew power input
rlabel locali s 298660 113169 298799 113387 6 VPWR
port 613 nsew power input
rlabel locali s 298660 113387 298661 113495 6 VPWR
port 613 nsew power input
rlabel locali s 1259 112809 1340 112917 6 VPWR
port 613 nsew power input
rlabel locali s 1121 112917 1340 113135 6 VPWR
port 613 nsew power input
rlabel locali s 1104 113135 1340 113169 6 VPWR
port 613 nsew power input
rlabel locali s 1121 113169 1340 113387 6 VPWR
port 613 nsew power input
rlabel locali s 1259 113387 1340 113495 6 VPWR
port 613 nsew power input
rlabel locali s 298660 113897 298661 114005 6 VPWR
port 613 nsew power input
rlabel locali s 298660 114005 298799 114223 6 VPWR
port 613 nsew power input
rlabel locali s 298660 114223 298816 114257 6 VPWR
port 613 nsew power input
rlabel locali s 298660 114257 298799 114475 6 VPWR
port 613 nsew power input
rlabel locali s 298660 114475 298661 114583 6 VPWR
port 613 nsew power input
rlabel locali s 1259 113897 1340 114005 6 VPWR
port 613 nsew power input
rlabel locali s 1121 114005 1340 114223 6 VPWR
port 613 nsew power input
rlabel locali s 1104 114223 1340 114257 6 VPWR
port 613 nsew power input
rlabel locali s 1121 114257 1340 114475 6 VPWR
port 613 nsew power input
rlabel locali s 1259 114475 1340 114583 6 VPWR
port 613 nsew power input
rlabel locali s 298660 114985 298661 115093 6 VPWR
port 613 nsew power input
rlabel locali s 298660 115093 298799 115311 6 VPWR
port 613 nsew power input
rlabel locali s 298660 115311 298816 115345 6 VPWR
port 613 nsew power input
rlabel locali s 298660 115345 298799 115563 6 VPWR
port 613 nsew power input
rlabel locali s 298660 115563 298661 115671 6 VPWR
port 613 nsew power input
rlabel locali s 1259 114985 1340 115093 6 VPWR
port 613 nsew power input
rlabel locali s 1121 115093 1340 115311 6 VPWR
port 613 nsew power input
rlabel locali s 1104 115311 1340 115345 6 VPWR
port 613 nsew power input
rlabel locali s 1121 115345 1340 115563 6 VPWR
port 613 nsew power input
rlabel locali s 1259 115563 1340 115671 6 VPWR
port 613 nsew power input
rlabel locali s 298660 116073 298661 116181 6 VPWR
port 613 nsew power input
rlabel locali s 298660 116181 298799 116399 6 VPWR
port 613 nsew power input
rlabel locali s 298660 116399 298816 116433 6 VPWR
port 613 nsew power input
rlabel locali s 298660 116433 298799 116651 6 VPWR
port 613 nsew power input
rlabel locali s 298660 116651 298661 116759 6 VPWR
port 613 nsew power input
rlabel locali s 1259 116073 1340 116181 6 VPWR
port 613 nsew power input
rlabel locali s 1121 116181 1340 116399 6 VPWR
port 613 nsew power input
rlabel locali s 1104 116399 1340 116433 6 VPWR
port 613 nsew power input
rlabel locali s 1121 116433 1340 116651 6 VPWR
port 613 nsew power input
rlabel locali s 1259 116651 1340 116759 6 VPWR
port 613 nsew power input
rlabel locali s 298660 117161 298661 117269 6 VPWR
port 613 nsew power input
rlabel locali s 298660 117269 298799 117487 6 VPWR
port 613 nsew power input
rlabel locali s 298660 117487 298816 117521 6 VPWR
port 613 nsew power input
rlabel locali s 298660 117521 298799 117739 6 VPWR
port 613 nsew power input
rlabel locali s 298660 117739 298661 117847 6 VPWR
port 613 nsew power input
rlabel locali s 1259 117161 1340 117269 6 VPWR
port 613 nsew power input
rlabel locali s 1121 117269 1340 117487 6 VPWR
port 613 nsew power input
rlabel locali s 1104 117487 1340 117521 6 VPWR
port 613 nsew power input
rlabel locali s 1121 117521 1340 117739 6 VPWR
port 613 nsew power input
rlabel locali s 1259 117739 1340 117847 6 VPWR
port 613 nsew power input
rlabel locali s 298660 118249 298661 118357 6 VPWR
port 613 nsew power input
rlabel locali s 298660 118357 298799 118575 6 VPWR
port 613 nsew power input
rlabel locali s 298660 118575 298816 118609 6 VPWR
port 613 nsew power input
rlabel locali s 298660 118609 298799 118827 6 VPWR
port 613 nsew power input
rlabel locali s 298660 118827 298661 118935 6 VPWR
port 613 nsew power input
rlabel locali s 1259 118249 1340 118357 6 VPWR
port 613 nsew power input
rlabel locali s 1121 118357 1340 118575 6 VPWR
port 613 nsew power input
rlabel locali s 1104 118575 1340 118609 6 VPWR
port 613 nsew power input
rlabel locali s 1121 118609 1340 118827 6 VPWR
port 613 nsew power input
rlabel locali s 1259 118827 1340 118935 6 VPWR
port 613 nsew power input
rlabel locali s 298660 119337 298661 119445 6 VPWR
port 613 nsew power input
rlabel locali s 298660 119445 298799 119663 6 VPWR
port 613 nsew power input
rlabel locali s 298660 119663 298816 119697 6 VPWR
port 613 nsew power input
rlabel locali s 298660 119697 298799 119915 6 VPWR
port 613 nsew power input
rlabel locali s 298660 119915 298661 120023 6 VPWR
port 613 nsew power input
rlabel locali s 1259 119337 1340 119445 6 VPWR
port 613 nsew power input
rlabel locali s 1121 119445 1340 119663 6 VPWR
port 613 nsew power input
rlabel locali s 1104 119663 1340 119697 6 VPWR
port 613 nsew power input
rlabel locali s 1121 119697 1340 119915 6 VPWR
port 613 nsew power input
rlabel locali s 1259 119915 1340 120023 6 VPWR
port 613 nsew power input
rlabel locali s 298660 120425 298661 120533 6 VPWR
port 613 nsew power input
rlabel locali s 298660 120533 298799 120751 6 VPWR
port 613 nsew power input
rlabel locali s 298660 120751 298816 120785 6 VPWR
port 613 nsew power input
rlabel locali s 298660 120785 298799 121003 6 VPWR
port 613 nsew power input
rlabel locali s 298660 121003 298661 121111 6 VPWR
port 613 nsew power input
rlabel locali s 1259 120425 1340 120533 6 VPWR
port 613 nsew power input
rlabel locali s 1121 120533 1340 120751 6 VPWR
port 613 nsew power input
rlabel locali s 1104 120751 1340 120785 6 VPWR
port 613 nsew power input
rlabel locali s 1121 120785 1340 121003 6 VPWR
port 613 nsew power input
rlabel locali s 1259 121003 1340 121111 6 VPWR
port 613 nsew power input
rlabel locali s 298660 121513 298661 121621 6 VPWR
port 613 nsew power input
rlabel locali s 298660 121621 298799 121839 6 VPWR
port 613 nsew power input
rlabel locali s 298660 121839 298816 121873 6 VPWR
port 613 nsew power input
rlabel locali s 298660 121873 298799 122091 6 VPWR
port 613 nsew power input
rlabel locali s 298660 122091 298661 122199 6 VPWR
port 613 nsew power input
rlabel locali s 1259 121513 1340 121621 6 VPWR
port 613 nsew power input
rlabel locali s 1121 121621 1340 121839 6 VPWR
port 613 nsew power input
rlabel locali s 1104 121839 1340 121873 6 VPWR
port 613 nsew power input
rlabel locali s 1121 121873 1340 122091 6 VPWR
port 613 nsew power input
rlabel locali s 1259 122091 1340 122199 6 VPWR
port 613 nsew power input
rlabel locali s 298660 122601 298661 122709 6 VPWR
port 613 nsew power input
rlabel locali s 298660 122709 298799 122927 6 VPWR
port 613 nsew power input
rlabel locali s 298660 122927 298816 122961 6 VPWR
port 613 nsew power input
rlabel locali s 298660 122961 298799 123179 6 VPWR
port 613 nsew power input
rlabel locali s 298660 123179 298661 123287 6 VPWR
port 613 nsew power input
rlabel locali s 1259 122601 1340 122709 6 VPWR
port 613 nsew power input
rlabel locali s 1121 122709 1340 122927 6 VPWR
port 613 nsew power input
rlabel locali s 1104 122927 1340 122961 6 VPWR
port 613 nsew power input
rlabel locali s 1121 122961 1340 123179 6 VPWR
port 613 nsew power input
rlabel locali s 1259 123179 1340 123287 6 VPWR
port 613 nsew power input
rlabel locali s 298660 123689 298661 123797 6 VPWR
port 613 nsew power input
rlabel locali s 298660 123797 298799 124015 6 VPWR
port 613 nsew power input
rlabel locali s 298660 124015 298816 124049 6 VPWR
port 613 nsew power input
rlabel locali s 298660 124049 298799 124267 6 VPWR
port 613 nsew power input
rlabel locali s 298660 124267 298661 124375 6 VPWR
port 613 nsew power input
rlabel locali s 1259 123689 1340 123797 6 VPWR
port 613 nsew power input
rlabel locali s 1121 123797 1340 124015 6 VPWR
port 613 nsew power input
rlabel locali s 1104 124015 1340 124049 6 VPWR
port 613 nsew power input
rlabel locali s 1121 124049 1340 124267 6 VPWR
port 613 nsew power input
rlabel locali s 1259 124267 1340 124375 6 VPWR
port 613 nsew power input
rlabel locali s 298660 124777 298661 124885 6 VPWR
port 613 nsew power input
rlabel locali s 298660 124885 298799 125103 6 VPWR
port 613 nsew power input
rlabel locali s 298660 125103 298816 125137 6 VPWR
port 613 nsew power input
rlabel locali s 298660 125137 298799 125355 6 VPWR
port 613 nsew power input
rlabel locali s 298660 125355 298661 125463 6 VPWR
port 613 nsew power input
rlabel locali s 1259 124777 1340 124885 6 VPWR
port 613 nsew power input
rlabel locali s 1121 124885 1340 125103 6 VPWR
port 613 nsew power input
rlabel locali s 1104 125103 1340 125137 6 VPWR
port 613 nsew power input
rlabel locali s 1121 125137 1340 125355 6 VPWR
port 613 nsew power input
rlabel locali s 1259 125355 1340 125463 6 VPWR
port 613 nsew power input
rlabel locali s 298660 125865 298661 125973 6 VPWR
port 613 nsew power input
rlabel locali s 298660 125973 298799 126191 6 VPWR
port 613 nsew power input
rlabel locali s 298660 126191 298816 126225 6 VPWR
port 613 nsew power input
rlabel locali s 298660 126225 298799 126443 6 VPWR
port 613 nsew power input
rlabel locali s 298660 126443 298661 126551 6 VPWR
port 613 nsew power input
rlabel locali s 1259 125865 1340 125973 6 VPWR
port 613 nsew power input
rlabel locali s 1121 125973 1340 126191 6 VPWR
port 613 nsew power input
rlabel locali s 1104 126191 1340 126225 6 VPWR
port 613 nsew power input
rlabel locali s 1121 126225 1340 126443 6 VPWR
port 613 nsew power input
rlabel locali s 1259 126443 1340 126551 6 VPWR
port 613 nsew power input
rlabel locali s 298660 126953 298661 127061 6 VPWR
port 613 nsew power input
rlabel locali s 298660 127061 298799 127279 6 VPWR
port 613 nsew power input
rlabel locali s 298660 127279 298816 127313 6 VPWR
port 613 nsew power input
rlabel locali s 298660 127313 298799 127531 6 VPWR
port 613 nsew power input
rlabel locali s 298660 127531 298661 127639 6 VPWR
port 613 nsew power input
rlabel locali s 1259 126953 1340 127061 6 VPWR
port 613 nsew power input
rlabel locali s 1121 127061 1340 127279 6 VPWR
port 613 nsew power input
rlabel locali s 1104 127279 1340 127313 6 VPWR
port 613 nsew power input
rlabel locali s 1121 127313 1340 127531 6 VPWR
port 613 nsew power input
rlabel locali s 1259 127531 1340 127639 6 VPWR
port 613 nsew power input
rlabel locali s 298660 128041 298661 128149 6 VPWR
port 613 nsew power input
rlabel locali s 298660 128149 298799 128367 6 VPWR
port 613 nsew power input
rlabel locali s 298660 128367 298816 128401 6 VPWR
port 613 nsew power input
rlabel locali s 298660 128401 298799 128619 6 VPWR
port 613 nsew power input
rlabel locali s 298660 128619 298661 128727 6 VPWR
port 613 nsew power input
rlabel locali s 1259 128041 1340 128149 6 VPWR
port 613 nsew power input
rlabel locali s 1121 128149 1340 128367 6 VPWR
port 613 nsew power input
rlabel locali s 1104 128367 1340 128401 6 VPWR
port 613 nsew power input
rlabel locali s 1121 128401 1340 128619 6 VPWR
port 613 nsew power input
rlabel locali s 1259 128619 1340 128727 6 VPWR
port 613 nsew power input
rlabel locali s 298660 129129 298661 129237 6 VPWR
port 613 nsew power input
rlabel locali s 298660 129237 298799 129455 6 VPWR
port 613 nsew power input
rlabel locali s 298660 129455 298816 129489 6 VPWR
port 613 nsew power input
rlabel locali s 298660 129489 298799 129707 6 VPWR
port 613 nsew power input
rlabel locali s 298660 129707 298661 129815 6 VPWR
port 613 nsew power input
rlabel locali s 1259 129129 1340 129237 6 VPWR
port 613 nsew power input
rlabel locali s 1121 129237 1340 129455 6 VPWR
port 613 nsew power input
rlabel locali s 1104 129455 1340 129489 6 VPWR
port 613 nsew power input
rlabel locali s 1121 129489 1340 129707 6 VPWR
port 613 nsew power input
rlabel locali s 1259 129707 1340 129815 6 VPWR
port 613 nsew power input
rlabel locali s 298660 130217 298661 130325 6 VPWR
port 613 nsew power input
rlabel locali s 298660 130325 298799 130543 6 VPWR
port 613 nsew power input
rlabel locali s 298660 130543 298816 130577 6 VPWR
port 613 nsew power input
rlabel locali s 298660 130577 298799 130795 6 VPWR
port 613 nsew power input
rlabel locali s 298660 130795 298661 130903 6 VPWR
port 613 nsew power input
rlabel locali s 1259 130217 1340 130325 6 VPWR
port 613 nsew power input
rlabel locali s 1121 130325 1340 130543 6 VPWR
port 613 nsew power input
rlabel locali s 1104 130543 1340 130577 6 VPWR
port 613 nsew power input
rlabel locali s 1121 130577 1340 130795 6 VPWR
port 613 nsew power input
rlabel locali s 1259 130795 1340 130903 6 VPWR
port 613 nsew power input
rlabel locali s 298660 131305 298661 131413 6 VPWR
port 613 nsew power input
rlabel locali s 298660 131413 298799 131631 6 VPWR
port 613 nsew power input
rlabel locali s 298660 131631 298816 131665 6 VPWR
port 613 nsew power input
rlabel locali s 298660 131665 298799 131883 6 VPWR
port 613 nsew power input
rlabel locali s 298660 131883 298661 131991 6 VPWR
port 613 nsew power input
rlabel locali s 1259 131305 1340 131413 6 VPWR
port 613 nsew power input
rlabel locali s 1121 131413 1340 131631 6 VPWR
port 613 nsew power input
rlabel locali s 1104 131631 1340 131665 6 VPWR
port 613 nsew power input
rlabel locali s 1121 131665 1340 131883 6 VPWR
port 613 nsew power input
rlabel locali s 1259 131883 1340 131991 6 VPWR
port 613 nsew power input
rlabel locali s 298660 132393 298661 132501 6 VPWR
port 613 nsew power input
rlabel locali s 298660 132501 298799 132719 6 VPWR
port 613 nsew power input
rlabel locali s 298660 132719 298816 132753 6 VPWR
port 613 nsew power input
rlabel locali s 298660 132753 298799 132971 6 VPWR
port 613 nsew power input
rlabel locali s 298660 132971 298661 133079 6 VPWR
port 613 nsew power input
rlabel locali s 1259 132393 1340 132501 6 VPWR
port 613 nsew power input
rlabel locali s 1121 132501 1340 132719 6 VPWR
port 613 nsew power input
rlabel locali s 1104 132719 1340 132753 6 VPWR
port 613 nsew power input
rlabel locali s 1121 132753 1340 132971 6 VPWR
port 613 nsew power input
rlabel locali s 1259 132971 1340 133079 6 VPWR
port 613 nsew power input
rlabel locali s 298660 133481 298661 133589 6 VPWR
port 613 nsew power input
rlabel locali s 298660 133589 298799 133807 6 VPWR
port 613 nsew power input
rlabel locali s 298660 133807 298816 133841 6 VPWR
port 613 nsew power input
rlabel locali s 298660 133841 298799 134059 6 VPWR
port 613 nsew power input
rlabel locali s 298660 134059 298661 134167 6 VPWR
port 613 nsew power input
rlabel locali s 1259 133481 1340 133589 6 VPWR
port 613 nsew power input
rlabel locali s 1121 133589 1340 133807 6 VPWR
port 613 nsew power input
rlabel locali s 1104 133807 1340 133841 6 VPWR
port 613 nsew power input
rlabel locali s 1121 133841 1340 134059 6 VPWR
port 613 nsew power input
rlabel locali s 1259 134059 1340 134167 6 VPWR
port 613 nsew power input
rlabel locali s 298660 134569 298661 134677 6 VPWR
port 613 nsew power input
rlabel locali s 298660 134677 298799 134895 6 VPWR
port 613 nsew power input
rlabel locali s 298660 134895 298816 134929 6 VPWR
port 613 nsew power input
rlabel locali s 298660 134929 298799 135147 6 VPWR
port 613 nsew power input
rlabel locali s 298660 135147 298661 135255 6 VPWR
port 613 nsew power input
rlabel locali s 1259 134569 1340 134677 6 VPWR
port 613 nsew power input
rlabel locali s 1121 134677 1340 134895 6 VPWR
port 613 nsew power input
rlabel locali s 1104 134895 1340 134929 6 VPWR
port 613 nsew power input
rlabel locali s 1121 134929 1340 135147 6 VPWR
port 613 nsew power input
rlabel locali s 1259 135147 1340 135255 6 VPWR
port 613 nsew power input
rlabel locali s 298660 135657 298661 135765 6 VPWR
port 613 nsew power input
rlabel locali s 298660 135765 298799 135983 6 VPWR
port 613 nsew power input
rlabel locali s 298660 135983 298816 136017 6 VPWR
port 613 nsew power input
rlabel locali s 298660 136017 298799 136235 6 VPWR
port 613 nsew power input
rlabel locali s 298660 136235 298661 136343 6 VPWR
port 613 nsew power input
rlabel locali s 1259 135657 1340 135765 6 VPWR
port 613 nsew power input
rlabel locali s 1121 135765 1340 135983 6 VPWR
port 613 nsew power input
rlabel locali s 1104 135983 1340 136017 6 VPWR
port 613 nsew power input
rlabel locali s 1121 136017 1340 136235 6 VPWR
port 613 nsew power input
rlabel locali s 1259 136235 1340 136343 6 VPWR
port 613 nsew power input
rlabel locali s 298660 136745 298661 136853 6 VPWR
port 613 nsew power input
rlabel locali s 298660 136853 298799 137071 6 VPWR
port 613 nsew power input
rlabel locali s 298660 137071 298816 137105 6 VPWR
port 613 nsew power input
rlabel locali s 298660 137105 298799 137323 6 VPWR
port 613 nsew power input
rlabel locali s 298660 137323 298661 137431 6 VPWR
port 613 nsew power input
rlabel locali s 1259 136745 1340 136853 6 VPWR
port 613 nsew power input
rlabel locali s 1121 136853 1340 137071 6 VPWR
port 613 nsew power input
rlabel locali s 1104 137071 1340 137105 6 VPWR
port 613 nsew power input
rlabel locali s 1121 137105 1340 137323 6 VPWR
port 613 nsew power input
rlabel locali s 1259 137323 1340 137431 6 VPWR
port 613 nsew power input
rlabel locali s 298660 137833 298661 137941 6 VPWR
port 613 nsew power input
rlabel locali s 298660 137941 298799 138159 6 VPWR
port 613 nsew power input
rlabel locali s 298660 138159 298816 138193 6 VPWR
port 613 nsew power input
rlabel locali s 298660 138193 298799 138411 6 VPWR
port 613 nsew power input
rlabel locali s 298660 138411 298661 138519 6 VPWR
port 613 nsew power input
rlabel locali s 1259 137833 1340 137941 6 VPWR
port 613 nsew power input
rlabel locali s 1121 137941 1340 138159 6 VPWR
port 613 nsew power input
rlabel locali s 1104 138159 1340 138193 6 VPWR
port 613 nsew power input
rlabel locali s 1121 138193 1340 138411 6 VPWR
port 613 nsew power input
rlabel locali s 1259 138411 1340 138519 6 VPWR
port 613 nsew power input
rlabel locali s 298660 138921 298661 139029 6 VPWR
port 613 nsew power input
rlabel locali s 298660 139029 298799 139247 6 VPWR
port 613 nsew power input
rlabel locali s 298660 139247 298816 139281 6 VPWR
port 613 nsew power input
rlabel locali s 298660 139281 298799 139499 6 VPWR
port 613 nsew power input
rlabel locali s 298660 139499 298661 139607 6 VPWR
port 613 nsew power input
rlabel locali s 1259 138921 1340 139029 6 VPWR
port 613 nsew power input
rlabel locali s 1121 139029 1340 139247 6 VPWR
port 613 nsew power input
rlabel locali s 1104 139247 1340 139281 6 VPWR
port 613 nsew power input
rlabel locali s 1121 139281 1340 139499 6 VPWR
port 613 nsew power input
rlabel locali s 1259 139499 1340 139607 6 VPWR
port 613 nsew power input
rlabel locali s 298660 140009 298661 140117 6 VPWR
port 613 nsew power input
rlabel locali s 298660 140117 298799 140335 6 VPWR
port 613 nsew power input
rlabel locali s 298660 140335 298816 140369 6 VPWR
port 613 nsew power input
rlabel locali s 298660 140369 298799 140587 6 VPWR
port 613 nsew power input
rlabel locali s 298660 140587 298661 140695 6 VPWR
port 613 nsew power input
rlabel locali s 1259 140009 1340 140117 6 VPWR
port 613 nsew power input
rlabel locali s 1121 140117 1340 140335 6 VPWR
port 613 nsew power input
rlabel locali s 1104 140335 1340 140369 6 VPWR
port 613 nsew power input
rlabel locali s 1121 140369 1340 140587 6 VPWR
port 613 nsew power input
rlabel locali s 1259 140587 1340 140695 6 VPWR
port 613 nsew power input
rlabel locali s 298660 141097 298661 141205 6 VPWR
port 613 nsew power input
rlabel locali s 298660 141205 298799 141423 6 VPWR
port 613 nsew power input
rlabel locali s 298660 141423 298816 141457 6 VPWR
port 613 nsew power input
rlabel locali s 298660 141457 298799 141675 6 VPWR
port 613 nsew power input
rlabel locali s 298660 141675 298661 141783 6 VPWR
port 613 nsew power input
rlabel locali s 1259 141097 1340 141205 6 VPWR
port 613 nsew power input
rlabel locali s 1121 141205 1340 141423 6 VPWR
port 613 nsew power input
rlabel locali s 1104 141423 1340 141457 6 VPWR
port 613 nsew power input
rlabel locali s 1121 141457 1340 141675 6 VPWR
port 613 nsew power input
rlabel locali s 1259 141675 1340 141783 6 VPWR
port 613 nsew power input
rlabel locali s 298660 142185 298661 142293 6 VPWR
port 613 nsew power input
rlabel locali s 298660 142293 298799 142511 6 VPWR
port 613 nsew power input
rlabel locali s 298660 142511 298816 142545 6 VPWR
port 613 nsew power input
rlabel locali s 298660 142545 298799 142763 6 VPWR
port 613 nsew power input
rlabel locali s 298660 142763 298661 142871 6 VPWR
port 613 nsew power input
rlabel locali s 1259 142185 1340 142293 6 VPWR
port 613 nsew power input
rlabel locali s 1121 142293 1340 142511 6 VPWR
port 613 nsew power input
rlabel locali s 1104 142511 1340 142545 6 VPWR
port 613 nsew power input
rlabel locali s 1121 142545 1340 142763 6 VPWR
port 613 nsew power input
rlabel locali s 1259 142763 1340 142871 6 VPWR
port 613 nsew power input
rlabel locali s 298660 143273 298661 143381 6 VPWR
port 613 nsew power input
rlabel locali s 298660 143381 298799 143599 6 VPWR
port 613 nsew power input
rlabel locali s 298660 143599 298816 143633 6 VPWR
port 613 nsew power input
rlabel locali s 298660 143633 298799 143851 6 VPWR
port 613 nsew power input
rlabel locali s 298660 143851 298661 143959 6 VPWR
port 613 nsew power input
rlabel locali s 1259 143273 1340 143381 6 VPWR
port 613 nsew power input
rlabel locali s 1121 143381 1340 143599 6 VPWR
port 613 nsew power input
rlabel locali s 1104 143599 1340 143633 6 VPWR
port 613 nsew power input
rlabel locali s 1121 143633 1340 143851 6 VPWR
port 613 nsew power input
rlabel locali s 1259 143851 1340 143959 6 VPWR
port 613 nsew power input
rlabel locali s 298660 144361 298661 144469 6 VPWR
port 613 nsew power input
rlabel locali s 298660 144469 298799 144687 6 VPWR
port 613 nsew power input
rlabel locali s 298660 144687 298816 144721 6 VPWR
port 613 nsew power input
rlabel locali s 298660 144721 298799 144939 6 VPWR
port 613 nsew power input
rlabel locali s 298660 144939 298661 145047 6 VPWR
port 613 nsew power input
rlabel locali s 1259 144361 1340 144469 6 VPWR
port 613 nsew power input
rlabel locali s 1121 144469 1340 144687 6 VPWR
port 613 nsew power input
rlabel locali s 1104 144687 1340 144721 6 VPWR
port 613 nsew power input
rlabel locali s 1121 144721 1340 144939 6 VPWR
port 613 nsew power input
rlabel locali s 1259 144939 1340 145047 6 VPWR
port 613 nsew power input
rlabel locali s 298660 145449 298661 145557 6 VPWR
port 613 nsew power input
rlabel locali s 298660 145557 298799 145775 6 VPWR
port 613 nsew power input
rlabel locali s 298660 145775 298816 145809 6 VPWR
port 613 nsew power input
rlabel locali s 298660 145809 298799 146027 6 VPWR
port 613 nsew power input
rlabel locali s 298660 146027 298661 146135 6 VPWR
port 613 nsew power input
rlabel locali s 1259 145449 1340 145557 6 VPWR
port 613 nsew power input
rlabel locali s 1121 145557 1340 145775 6 VPWR
port 613 nsew power input
rlabel locali s 1104 145775 1340 145809 6 VPWR
port 613 nsew power input
rlabel locali s 1121 145809 1340 146027 6 VPWR
port 613 nsew power input
rlabel locali s 1259 146027 1340 146135 6 VPWR
port 613 nsew power input
rlabel locali s 298660 146537 298661 146645 6 VPWR
port 613 nsew power input
rlabel locali s 298660 146645 298799 146863 6 VPWR
port 613 nsew power input
rlabel locali s 298660 146863 298816 146897 6 VPWR
port 613 nsew power input
rlabel locali s 298660 146897 298799 147115 6 VPWR
port 613 nsew power input
rlabel locali s 298660 147115 298661 147223 6 VPWR
port 613 nsew power input
rlabel locali s 1259 146537 1340 146645 6 VPWR
port 613 nsew power input
rlabel locali s 1121 146645 1340 146863 6 VPWR
port 613 nsew power input
rlabel locali s 1104 146863 1340 146897 6 VPWR
port 613 nsew power input
rlabel locali s 1121 146897 1340 147115 6 VPWR
port 613 nsew power input
rlabel locali s 1259 147115 1340 147223 6 VPWR
port 613 nsew power input
rlabel locali s 298660 147625 298661 147733 6 VPWR
port 613 nsew power input
rlabel locali s 298660 147733 298799 147951 6 VPWR
port 613 nsew power input
rlabel locali s 298660 147951 298816 147985 6 VPWR
port 613 nsew power input
rlabel locali s 298660 147985 298799 148203 6 VPWR
port 613 nsew power input
rlabel locali s 298660 148203 298661 148311 6 VPWR
port 613 nsew power input
rlabel locali s 1259 147625 1340 147733 6 VPWR
port 613 nsew power input
rlabel locali s 1121 147733 1340 147951 6 VPWR
port 613 nsew power input
rlabel locali s 1104 147951 1340 147985 6 VPWR
port 613 nsew power input
rlabel locali s 1121 147985 1340 148203 6 VPWR
port 613 nsew power input
rlabel locali s 1259 148203 1340 148311 6 VPWR
port 613 nsew power input
rlabel locali s 298660 148713 298661 148821 6 VPWR
port 613 nsew power input
rlabel locali s 298660 148821 298799 149039 6 VPWR
port 613 nsew power input
rlabel locali s 298660 149039 298816 149073 6 VPWR
port 613 nsew power input
rlabel locali s 298660 149073 298799 149291 6 VPWR
port 613 nsew power input
rlabel locali s 298660 149291 298661 149399 6 VPWR
port 613 nsew power input
rlabel locali s 1259 148713 1340 148821 6 VPWR
port 613 nsew power input
rlabel locali s 1121 148821 1340 149039 6 VPWR
port 613 nsew power input
rlabel locali s 1104 149039 1340 149073 6 VPWR
port 613 nsew power input
rlabel locali s 1121 149073 1340 149291 6 VPWR
port 613 nsew power input
rlabel locali s 1259 149291 1340 149399 6 VPWR
port 613 nsew power input
rlabel locali s 298660 149801 298661 149909 6 VPWR
port 613 nsew power input
rlabel locali s 298660 149909 298799 150127 6 VPWR
port 613 nsew power input
rlabel locali s 298660 150127 298816 150161 6 VPWR
port 613 nsew power input
rlabel locali s 298660 150161 298799 150379 6 VPWR
port 613 nsew power input
rlabel locali s 298660 150379 298661 150487 6 VPWR
port 613 nsew power input
rlabel locali s 1259 149801 1340 149909 6 VPWR
port 613 nsew power input
rlabel locali s 1121 149909 1340 150127 6 VPWR
port 613 nsew power input
rlabel locali s 1104 150127 1340 150161 6 VPWR
port 613 nsew power input
rlabel locali s 1121 150161 1340 150379 6 VPWR
port 613 nsew power input
rlabel locali s 1259 150379 1340 150487 6 VPWR
port 613 nsew power input
rlabel locali s 298660 150889 298661 150997 6 VPWR
port 613 nsew power input
rlabel locali s 298660 150997 298799 151215 6 VPWR
port 613 nsew power input
rlabel locali s 298660 151215 298816 151249 6 VPWR
port 613 nsew power input
rlabel locali s 298660 151249 298799 151467 6 VPWR
port 613 nsew power input
rlabel locali s 298660 151467 298661 151575 6 VPWR
port 613 nsew power input
rlabel locali s 1259 150889 1340 150997 6 VPWR
port 613 nsew power input
rlabel locali s 1121 150997 1340 151215 6 VPWR
port 613 nsew power input
rlabel locali s 1104 151215 1340 151249 6 VPWR
port 613 nsew power input
rlabel locali s 1121 151249 1340 151467 6 VPWR
port 613 nsew power input
rlabel locali s 1259 151467 1340 151575 6 VPWR
port 613 nsew power input
rlabel locali s 298660 151977 298661 152085 6 VPWR
port 613 nsew power input
rlabel locali s 298660 152085 298799 152303 6 VPWR
port 613 nsew power input
rlabel locali s 298660 152303 298816 152337 6 VPWR
port 613 nsew power input
rlabel locali s 298660 152337 298799 152555 6 VPWR
port 613 nsew power input
rlabel locali s 298660 152555 298661 152663 6 VPWR
port 613 nsew power input
rlabel locali s 1259 151977 1340 152085 6 VPWR
port 613 nsew power input
rlabel locali s 1121 152085 1340 152303 6 VPWR
port 613 nsew power input
rlabel locali s 1104 152303 1340 152337 6 VPWR
port 613 nsew power input
rlabel locali s 1121 152337 1340 152555 6 VPWR
port 613 nsew power input
rlabel locali s 1259 152555 1340 152663 6 VPWR
port 613 nsew power input
rlabel locali s 298660 153065 298661 153173 6 VPWR
port 613 nsew power input
rlabel locali s 298660 153173 298799 153391 6 VPWR
port 613 nsew power input
rlabel locali s 298660 153391 298816 153425 6 VPWR
port 613 nsew power input
rlabel locali s 298660 153425 298799 153643 6 VPWR
port 613 nsew power input
rlabel locali s 298660 153643 298661 153751 6 VPWR
port 613 nsew power input
rlabel locali s 1259 153065 1340 153173 6 VPWR
port 613 nsew power input
rlabel locali s 1121 153173 1340 153391 6 VPWR
port 613 nsew power input
rlabel locali s 1104 153391 1340 153425 6 VPWR
port 613 nsew power input
rlabel locali s 1121 153425 1340 153643 6 VPWR
port 613 nsew power input
rlabel locali s 1259 153643 1340 153751 6 VPWR
port 613 nsew power input
rlabel locali s 298660 154153 298661 154261 6 VPWR
port 613 nsew power input
rlabel locali s 298660 154261 298799 154479 6 VPWR
port 613 nsew power input
rlabel locali s 298660 154479 298816 154513 6 VPWR
port 613 nsew power input
rlabel locali s 298660 154513 298799 154731 6 VPWR
port 613 nsew power input
rlabel locali s 298660 154731 298661 154839 6 VPWR
port 613 nsew power input
rlabel locali s 1259 154153 1340 154261 6 VPWR
port 613 nsew power input
rlabel locali s 1121 154261 1340 154479 6 VPWR
port 613 nsew power input
rlabel locali s 1104 154479 1340 154513 6 VPWR
port 613 nsew power input
rlabel locali s 1121 154513 1340 154731 6 VPWR
port 613 nsew power input
rlabel locali s 1259 154731 1340 154839 6 VPWR
port 613 nsew power input
rlabel locali s 298660 155241 298661 155349 6 VPWR
port 613 nsew power input
rlabel locali s 298660 155349 298799 155567 6 VPWR
port 613 nsew power input
rlabel locali s 298660 155567 298816 155601 6 VPWR
port 613 nsew power input
rlabel locali s 298660 155601 298799 155819 6 VPWR
port 613 nsew power input
rlabel locali s 298660 155819 298661 155927 6 VPWR
port 613 nsew power input
rlabel locali s 1259 155241 1340 155349 6 VPWR
port 613 nsew power input
rlabel locali s 1121 155349 1340 155567 6 VPWR
port 613 nsew power input
rlabel locali s 1104 155567 1340 155601 6 VPWR
port 613 nsew power input
rlabel locali s 1121 155601 1340 155819 6 VPWR
port 613 nsew power input
rlabel locali s 1259 155819 1340 155927 6 VPWR
port 613 nsew power input
rlabel locali s 298660 156329 298661 156437 6 VPWR
port 613 nsew power input
rlabel locali s 298660 156437 298799 156655 6 VPWR
port 613 nsew power input
rlabel locali s 298660 156655 298816 156689 6 VPWR
port 613 nsew power input
rlabel locali s 298660 156689 298799 156907 6 VPWR
port 613 nsew power input
rlabel locali s 298660 156907 298661 157015 6 VPWR
port 613 nsew power input
rlabel locali s 1259 156329 1340 156437 6 VPWR
port 613 nsew power input
rlabel locali s 1121 156437 1340 156655 6 VPWR
port 613 nsew power input
rlabel locali s 1104 156655 1340 156689 6 VPWR
port 613 nsew power input
rlabel locali s 1121 156689 1340 156907 6 VPWR
port 613 nsew power input
rlabel locali s 1259 156907 1340 157015 6 VPWR
port 613 nsew power input
rlabel locali s 298660 157417 298661 157525 6 VPWR
port 613 nsew power input
rlabel locali s 298660 157525 298799 157743 6 VPWR
port 613 nsew power input
rlabel locali s 298660 157743 298816 157777 6 VPWR
port 613 nsew power input
rlabel locali s 298660 157777 298799 157995 6 VPWR
port 613 nsew power input
rlabel locali s 298660 157995 298661 158103 6 VPWR
port 613 nsew power input
rlabel locali s 1259 157417 1340 157525 6 VPWR
port 613 nsew power input
rlabel locali s 1121 157525 1340 157743 6 VPWR
port 613 nsew power input
rlabel locali s 1104 157743 1340 157777 6 VPWR
port 613 nsew power input
rlabel locali s 1121 157777 1340 157995 6 VPWR
port 613 nsew power input
rlabel locali s 1259 157995 1340 158103 6 VPWR
port 613 nsew power input
rlabel locali s 298660 158505 298661 158613 6 VPWR
port 613 nsew power input
rlabel locali s 298660 158613 298799 158831 6 VPWR
port 613 nsew power input
rlabel locali s 298660 158831 298816 158865 6 VPWR
port 613 nsew power input
rlabel locali s 298660 158865 298799 159083 6 VPWR
port 613 nsew power input
rlabel locali s 298660 159083 298661 159191 6 VPWR
port 613 nsew power input
rlabel locali s 1259 158505 1340 158613 6 VPWR
port 613 nsew power input
rlabel locali s 1121 158613 1340 158831 6 VPWR
port 613 nsew power input
rlabel locali s 1104 158831 1340 158865 6 VPWR
port 613 nsew power input
rlabel locali s 1121 158865 1340 159083 6 VPWR
port 613 nsew power input
rlabel locali s 1259 159083 1340 159191 6 VPWR
port 613 nsew power input
rlabel locali s 298660 159593 298661 159701 6 VPWR
port 613 nsew power input
rlabel locali s 298660 159701 298799 159919 6 VPWR
port 613 nsew power input
rlabel locali s 298660 159919 298816 159953 6 VPWR
port 613 nsew power input
rlabel locali s 298660 159953 298799 160171 6 VPWR
port 613 nsew power input
rlabel locali s 298660 160171 298661 160279 6 VPWR
port 613 nsew power input
rlabel locali s 1259 159593 1340 159701 6 VPWR
port 613 nsew power input
rlabel locali s 1121 159701 1340 159919 6 VPWR
port 613 nsew power input
rlabel locali s 1104 159919 1340 159953 6 VPWR
port 613 nsew power input
rlabel locali s 1121 159953 1340 160171 6 VPWR
port 613 nsew power input
rlabel locali s 1259 160171 1340 160279 6 VPWR
port 613 nsew power input
rlabel locali s 298660 160681 298661 160789 6 VPWR
port 613 nsew power input
rlabel locali s 298660 160789 298799 161007 6 VPWR
port 613 nsew power input
rlabel locali s 298660 161007 298816 161041 6 VPWR
port 613 nsew power input
rlabel locali s 298660 161041 298799 161259 6 VPWR
port 613 nsew power input
rlabel locali s 298660 161259 298661 161367 6 VPWR
port 613 nsew power input
rlabel locali s 1259 160681 1340 160789 6 VPWR
port 613 nsew power input
rlabel locali s 1121 160789 1340 161007 6 VPWR
port 613 nsew power input
rlabel locali s 1104 161007 1340 161041 6 VPWR
port 613 nsew power input
rlabel locali s 1121 161041 1340 161259 6 VPWR
port 613 nsew power input
rlabel locali s 1259 161259 1340 161367 6 VPWR
port 613 nsew power input
rlabel locali s 298660 161769 298661 161877 6 VPWR
port 613 nsew power input
rlabel locali s 298660 161877 298799 162095 6 VPWR
port 613 nsew power input
rlabel locali s 298660 162095 298816 162129 6 VPWR
port 613 nsew power input
rlabel locali s 298660 162129 298799 162347 6 VPWR
port 613 nsew power input
rlabel locali s 298660 162347 298661 162455 6 VPWR
port 613 nsew power input
rlabel locali s 1259 161769 1340 161877 6 VPWR
port 613 nsew power input
rlabel locali s 1121 161877 1340 162095 6 VPWR
port 613 nsew power input
rlabel locali s 1104 162095 1340 162129 6 VPWR
port 613 nsew power input
rlabel locali s 1121 162129 1340 162347 6 VPWR
port 613 nsew power input
rlabel locali s 1259 162347 1340 162455 6 VPWR
port 613 nsew power input
rlabel locali s 298660 162857 298661 162965 6 VPWR
port 613 nsew power input
rlabel locali s 298660 162965 298799 163183 6 VPWR
port 613 nsew power input
rlabel locali s 298660 163183 298816 163217 6 VPWR
port 613 nsew power input
rlabel locali s 298660 163217 298799 163435 6 VPWR
port 613 nsew power input
rlabel locali s 298660 163435 298661 163543 6 VPWR
port 613 nsew power input
rlabel locali s 1259 162857 1340 162965 6 VPWR
port 613 nsew power input
rlabel locali s 1121 162965 1340 163183 6 VPWR
port 613 nsew power input
rlabel locali s 1104 163183 1340 163217 6 VPWR
port 613 nsew power input
rlabel locali s 1121 163217 1340 163435 6 VPWR
port 613 nsew power input
rlabel locali s 1259 163435 1340 163543 6 VPWR
port 613 nsew power input
rlabel locali s 298660 163945 298661 164053 6 VPWR
port 613 nsew power input
rlabel locali s 298660 164053 298799 164271 6 VPWR
port 613 nsew power input
rlabel locali s 298660 164271 298816 164305 6 VPWR
port 613 nsew power input
rlabel locali s 298660 164305 298799 164523 6 VPWR
port 613 nsew power input
rlabel locali s 298660 164523 298661 164631 6 VPWR
port 613 nsew power input
rlabel locali s 1259 163945 1340 164053 6 VPWR
port 613 nsew power input
rlabel locali s 1121 164053 1340 164271 6 VPWR
port 613 nsew power input
rlabel locali s 1104 164271 1340 164305 6 VPWR
port 613 nsew power input
rlabel locali s 1121 164305 1340 164523 6 VPWR
port 613 nsew power input
rlabel locali s 1259 164523 1340 164631 6 VPWR
port 613 nsew power input
rlabel locali s 298660 165033 298661 165141 6 VPWR
port 613 nsew power input
rlabel locali s 298660 165141 298799 165359 6 VPWR
port 613 nsew power input
rlabel locali s 298660 165359 298816 165393 6 VPWR
port 613 nsew power input
rlabel locali s 298660 165393 298799 165611 6 VPWR
port 613 nsew power input
rlabel locali s 298660 165611 298661 165719 6 VPWR
port 613 nsew power input
rlabel locali s 1259 165033 1340 165141 6 VPWR
port 613 nsew power input
rlabel locali s 1121 165141 1340 165359 6 VPWR
port 613 nsew power input
rlabel locali s 1104 165359 1340 165393 6 VPWR
port 613 nsew power input
rlabel locali s 1121 165393 1340 165611 6 VPWR
port 613 nsew power input
rlabel locali s 1259 165611 1340 165719 6 VPWR
port 613 nsew power input
rlabel locali s 298660 166121 298661 166229 6 VPWR
port 613 nsew power input
rlabel locali s 298660 166229 298799 166447 6 VPWR
port 613 nsew power input
rlabel locali s 298660 166447 298816 166481 6 VPWR
port 613 nsew power input
rlabel locali s 298660 166481 298799 166699 6 VPWR
port 613 nsew power input
rlabel locali s 298660 166699 298661 166807 6 VPWR
port 613 nsew power input
rlabel locali s 1259 166121 1340 166229 6 VPWR
port 613 nsew power input
rlabel locali s 1121 166229 1340 166447 6 VPWR
port 613 nsew power input
rlabel locali s 1104 166447 1340 166481 6 VPWR
port 613 nsew power input
rlabel locali s 1121 166481 1340 166699 6 VPWR
port 613 nsew power input
rlabel locali s 1259 166699 1340 166807 6 VPWR
port 613 nsew power input
rlabel locali s 298660 167209 298661 167317 6 VPWR
port 613 nsew power input
rlabel locali s 298660 167317 298799 167535 6 VPWR
port 613 nsew power input
rlabel locali s 298660 167535 298816 167569 6 VPWR
port 613 nsew power input
rlabel locali s 298660 167569 298799 167787 6 VPWR
port 613 nsew power input
rlabel locali s 298660 167787 298661 167895 6 VPWR
port 613 nsew power input
rlabel locali s 1259 167209 1340 167317 6 VPWR
port 613 nsew power input
rlabel locali s 1121 167317 1340 167535 6 VPWR
port 613 nsew power input
rlabel locali s 1104 167535 1340 167569 6 VPWR
port 613 nsew power input
rlabel locali s 1121 167569 1340 167787 6 VPWR
port 613 nsew power input
rlabel locali s 1259 167787 1340 167895 6 VPWR
port 613 nsew power input
rlabel locali s 298660 168297 298661 168405 6 VPWR
port 613 nsew power input
rlabel locali s 298660 168405 298799 168623 6 VPWR
port 613 nsew power input
rlabel locali s 298660 168623 298816 168657 6 VPWR
port 613 nsew power input
rlabel locali s 298660 168657 298799 168875 6 VPWR
port 613 nsew power input
rlabel locali s 298660 168875 298661 168983 6 VPWR
port 613 nsew power input
rlabel locali s 1259 168297 1340 168405 6 VPWR
port 613 nsew power input
rlabel locali s 1121 168405 1340 168623 6 VPWR
port 613 nsew power input
rlabel locali s 1104 168623 1340 168657 6 VPWR
port 613 nsew power input
rlabel locali s 1121 168657 1340 168875 6 VPWR
port 613 nsew power input
rlabel locali s 1259 168875 1340 168983 6 VPWR
port 613 nsew power input
rlabel locali s 298660 169385 298661 169493 6 VPWR
port 613 nsew power input
rlabel locali s 298660 169493 298799 169711 6 VPWR
port 613 nsew power input
rlabel locali s 298660 169711 298816 169745 6 VPWR
port 613 nsew power input
rlabel locali s 298660 169745 298799 169963 6 VPWR
port 613 nsew power input
rlabel locali s 298660 169963 298661 170071 6 VPWR
port 613 nsew power input
rlabel locali s 1259 169385 1340 169493 6 VPWR
port 613 nsew power input
rlabel locali s 1121 169493 1340 169711 6 VPWR
port 613 nsew power input
rlabel locali s 1104 169711 1340 169745 6 VPWR
port 613 nsew power input
rlabel locali s 1121 169745 1340 169963 6 VPWR
port 613 nsew power input
rlabel locali s 1259 169963 1340 170071 6 VPWR
port 613 nsew power input
rlabel locali s 298660 170473 298661 170581 6 VPWR
port 613 nsew power input
rlabel locali s 298660 170581 298799 170799 6 VPWR
port 613 nsew power input
rlabel locali s 298660 170799 298816 170833 6 VPWR
port 613 nsew power input
rlabel locali s 298660 170833 298799 171051 6 VPWR
port 613 nsew power input
rlabel locali s 298660 171051 298661 171159 6 VPWR
port 613 nsew power input
rlabel locali s 1259 170473 1340 170581 6 VPWR
port 613 nsew power input
rlabel locali s 1121 170581 1340 170799 6 VPWR
port 613 nsew power input
rlabel locali s 1104 170799 1340 170833 6 VPWR
port 613 nsew power input
rlabel locali s 1121 170833 1340 171051 6 VPWR
port 613 nsew power input
rlabel locali s 1259 171051 1340 171159 6 VPWR
port 613 nsew power input
rlabel locali s 298660 171561 298661 171669 6 VPWR
port 613 nsew power input
rlabel locali s 298660 171669 298799 171887 6 VPWR
port 613 nsew power input
rlabel locali s 298660 171887 298816 171921 6 VPWR
port 613 nsew power input
rlabel locali s 298660 171921 298799 172139 6 VPWR
port 613 nsew power input
rlabel locali s 298660 172139 298661 172247 6 VPWR
port 613 nsew power input
rlabel locali s 1259 171561 1340 171669 6 VPWR
port 613 nsew power input
rlabel locali s 1121 171669 1340 171887 6 VPWR
port 613 nsew power input
rlabel locali s 1104 171887 1340 171921 6 VPWR
port 613 nsew power input
rlabel locali s 1121 171921 1340 172139 6 VPWR
port 613 nsew power input
rlabel locali s 1259 172139 1340 172247 6 VPWR
port 613 nsew power input
rlabel locali s 298660 172649 298661 172757 6 VPWR
port 613 nsew power input
rlabel locali s 298660 172757 298799 172975 6 VPWR
port 613 nsew power input
rlabel locali s 298660 172975 298816 173009 6 VPWR
port 613 nsew power input
rlabel locali s 298660 173009 298799 173227 6 VPWR
port 613 nsew power input
rlabel locali s 298660 173227 298661 173335 6 VPWR
port 613 nsew power input
rlabel locali s 1259 172649 1340 172757 6 VPWR
port 613 nsew power input
rlabel locali s 1121 172757 1340 172975 6 VPWR
port 613 nsew power input
rlabel locali s 1104 172975 1340 173009 6 VPWR
port 613 nsew power input
rlabel locali s 1121 173009 1340 173227 6 VPWR
port 613 nsew power input
rlabel locali s 1259 173227 1340 173335 6 VPWR
port 613 nsew power input
rlabel locali s 298660 173737 298661 173845 6 VPWR
port 613 nsew power input
rlabel locali s 298660 173845 298799 174063 6 VPWR
port 613 nsew power input
rlabel locali s 298660 174063 298816 174097 6 VPWR
port 613 nsew power input
rlabel locali s 298660 174097 298799 174315 6 VPWR
port 613 nsew power input
rlabel locali s 298660 174315 298661 174423 6 VPWR
port 613 nsew power input
rlabel locali s 1259 173737 1340 173845 6 VPWR
port 613 nsew power input
rlabel locali s 1121 173845 1340 174063 6 VPWR
port 613 nsew power input
rlabel locali s 1104 174063 1340 174097 6 VPWR
port 613 nsew power input
rlabel locali s 1121 174097 1340 174315 6 VPWR
port 613 nsew power input
rlabel locali s 1259 174315 1340 174423 6 VPWR
port 613 nsew power input
rlabel locali s 298660 174825 298661 174933 6 VPWR
port 613 nsew power input
rlabel locali s 298660 174933 298799 175151 6 VPWR
port 613 nsew power input
rlabel locali s 298660 175151 298816 175185 6 VPWR
port 613 nsew power input
rlabel locali s 298660 175185 298799 175403 6 VPWR
port 613 nsew power input
rlabel locali s 298660 175403 298661 175511 6 VPWR
port 613 nsew power input
rlabel locali s 1259 174825 1340 174933 6 VPWR
port 613 nsew power input
rlabel locali s 1121 174933 1340 175151 6 VPWR
port 613 nsew power input
rlabel locali s 1104 175151 1340 175185 6 VPWR
port 613 nsew power input
rlabel locali s 1121 175185 1340 175403 6 VPWR
port 613 nsew power input
rlabel locali s 1259 175403 1340 175511 6 VPWR
port 613 nsew power input
rlabel locali s 298660 175913 298661 176021 6 VPWR
port 613 nsew power input
rlabel locali s 298660 176021 298799 176239 6 VPWR
port 613 nsew power input
rlabel locali s 298660 176239 298816 176273 6 VPWR
port 613 nsew power input
rlabel locali s 298660 176273 298799 176491 6 VPWR
port 613 nsew power input
rlabel locali s 298660 176491 298661 176599 6 VPWR
port 613 nsew power input
rlabel locali s 1259 175913 1340 176021 6 VPWR
port 613 nsew power input
rlabel locali s 1121 176021 1340 176239 6 VPWR
port 613 nsew power input
rlabel locali s 1104 176239 1340 176273 6 VPWR
port 613 nsew power input
rlabel locali s 1121 176273 1340 176491 6 VPWR
port 613 nsew power input
rlabel locali s 1259 176491 1340 176599 6 VPWR
port 613 nsew power input
rlabel locali s 298660 177001 298661 177109 6 VPWR
port 613 nsew power input
rlabel locali s 298660 177109 298799 177327 6 VPWR
port 613 nsew power input
rlabel locali s 298660 177327 298816 177361 6 VPWR
port 613 nsew power input
rlabel locali s 298660 177361 298799 177579 6 VPWR
port 613 nsew power input
rlabel locali s 298660 177579 298661 177687 6 VPWR
port 613 nsew power input
rlabel locali s 1259 177001 1340 177109 6 VPWR
port 613 nsew power input
rlabel locali s 1121 177109 1340 177327 6 VPWR
port 613 nsew power input
rlabel locali s 1104 177327 1340 177361 6 VPWR
port 613 nsew power input
rlabel locali s 1121 177361 1340 177579 6 VPWR
port 613 nsew power input
rlabel locali s 1259 177579 1340 177687 6 VPWR
port 613 nsew power input
rlabel locali s 298660 178089 298661 178197 6 VPWR
port 613 nsew power input
rlabel locali s 298660 178197 298799 178415 6 VPWR
port 613 nsew power input
rlabel locali s 298660 178415 298816 178449 6 VPWR
port 613 nsew power input
rlabel locali s 298660 178449 298799 178667 6 VPWR
port 613 nsew power input
rlabel locali s 298660 178667 298661 178775 6 VPWR
port 613 nsew power input
rlabel locali s 1259 178089 1340 178197 6 VPWR
port 613 nsew power input
rlabel locali s 1121 178197 1340 178415 6 VPWR
port 613 nsew power input
rlabel locali s 1104 178415 1340 178449 6 VPWR
port 613 nsew power input
rlabel locali s 1121 178449 1340 178667 6 VPWR
port 613 nsew power input
rlabel locali s 1259 178667 1340 178775 6 VPWR
port 613 nsew power input
rlabel locali s 298660 179177 298661 179285 6 VPWR
port 613 nsew power input
rlabel locali s 298660 179285 298799 179503 6 VPWR
port 613 nsew power input
rlabel locali s 298660 179503 298816 179537 6 VPWR
port 613 nsew power input
rlabel locali s 298660 179537 298799 179755 6 VPWR
port 613 nsew power input
rlabel locali s 298660 179755 298661 179863 6 VPWR
port 613 nsew power input
rlabel locali s 1259 179177 1340 179285 6 VPWR
port 613 nsew power input
rlabel locali s 1121 179285 1340 179503 6 VPWR
port 613 nsew power input
rlabel locali s 1104 179503 1340 179537 6 VPWR
port 613 nsew power input
rlabel locali s 1121 179537 1340 179755 6 VPWR
port 613 nsew power input
rlabel locali s 1259 179755 1340 179863 6 VPWR
port 613 nsew power input
rlabel locali s 298660 180265 298661 180373 6 VPWR
port 613 nsew power input
rlabel locali s 298660 180373 298799 180591 6 VPWR
port 613 nsew power input
rlabel locali s 298660 180591 298816 180625 6 VPWR
port 613 nsew power input
rlabel locali s 298660 180625 298799 180843 6 VPWR
port 613 nsew power input
rlabel locali s 298660 180843 298661 180951 6 VPWR
port 613 nsew power input
rlabel locali s 1259 180265 1340 180373 6 VPWR
port 613 nsew power input
rlabel locali s 1121 180373 1340 180591 6 VPWR
port 613 nsew power input
rlabel locali s 1104 180591 1340 180625 6 VPWR
port 613 nsew power input
rlabel locali s 1121 180625 1340 180843 6 VPWR
port 613 nsew power input
rlabel locali s 1259 180843 1340 180951 6 VPWR
port 613 nsew power input
rlabel locali s 298660 181353 298661 181461 6 VPWR
port 613 nsew power input
rlabel locali s 298660 181461 298799 181679 6 VPWR
port 613 nsew power input
rlabel locali s 298660 181679 298816 181713 6 VPWR
port 613 nsew power input
rlabel locali s 298660 181713 298799 181931 6 VPWR
port 613 nsew power input
rlabel locali s 298660 181931 298661 182039 6 VPWR
port 613 nsew power input
rlabel locali s 1259 181353 1340 181461 6 VPWR
port 613 nsew power input
rlabel locali s 1121 181461 1340 181679 6 VPWR
port 613 nsew power input
rlabel locali s 1104 181679 1340 181713 6 VPWR
port 613 nsew power input
rlabel locali s 1121 181713 1340 181931 6 VPWR
port 613 nsew power input
rlabel locali s 1259 181931 1340 182039 6 VPWR
port 613 nsew power input
rlabel locali s 298660 182441 298661 182549 6 VPWR
port 613 nsew power input
rlabel locali s 298660 182549 298799 182767 6 VPWR
port 613 nsew power input
rlabel locali s 298660 182767 298816 182801 6 VPWR
port 613 nsew power input
rlabel locali s 298660 182801 298799 183019 6 VPWR
port 613 nsew power input
rlabel locali s 298660 183019 298661 183127 6 VPWR
port 613 nsew power input
rlabel locali s 1259 182441 1340 182549 6 VPWR
port 613 nsew power input
rlabel locali s 1121 182549 1340 182767 6 VPWR
port 613 nsew power input
rlabel locali s 1104 182767 1340 182801 6 VPWR
port 613 nsew power input
rlabel locali s 1121 182801 1340 183019 6 VPWR
port 613 nsew power input
rlabel locali s 1259 183019 1340 183127 6 VPWR
port 613 nsew power input
rlabel locali s 298660 183529 298661 183637 6 VPWR
port 613 nsew power input
rlabel locali s 298660 183637 298799 183855 6 VPWR
port 613 nsew power input
rlabel locali s 298660 183855 298816 183889 6 VPWR
port 613 nsew power input
rlabel locali s 298660 183889 298799 184107 6 VPWR
port 613 nsew power input
rlabel locali s 298660 184107 298661 184215 6 VPWR
port 613 nsew power input
rlabel locali s 1259 183529 1340 183637 6 VPWR
port 613 nsew power input
rlabel locali s 1121 183637 1340 183855 6 VPWR
port 613 nsew power input
rlabel locali s 1104 183855 1340 183889 6 VPWR
port 613 nsew power input
rlabel locali s 1121 183889 1340 184107 6 VPWR
port 613 nsew power input
rlabel locali s 1259 184107 1340 184215 6 VPWR
port 613 nsew power input
rlabel locali s 298660 184617 298661 184725 6 VPWR
port 613 nsew power input
rlabel locali s 298660 184725 298799 184943 6 VPWR
port 613 nsew power input
rlabel locali s 298660 184943 298816 184977 6 VPWR
port 613 nsew power input
rlabel locali s 298660 184977 298799 185195 6 VPWR
port 613 nsew power input
rlabel locali s 298660 185195 298661 185303 6 VPWR
port 613 nsew power input
rlabel locali s 1259 184617 1340 184725 6 VPWR
port 613 nsew power input
rlabel locali s 1121 184725 1340 184943 6 VPWR
port 613 nsew power input
rlabel locali s 1104 184943 1340 184977 6 VPWR
port 613 nsew power input
rlabel locali s 1121 184977 1340 185195 6 VPWR
port 613 nsew power input
rlabel locali s 1259 185195 1340 185303 6 VPWR
port 613 nsew power input
rlabel locali s 298660 185705 298661 185813 6 VPWR
port 613 nsew power input
rlabel locali s 298660 185813 298799 186031 6 VPWR
port 613 nsew power input
rlabel locali s 298660 186031 298816 186065 6 VPWR
port 613 nsew power input
rlabel locali s 298660 186065 298799 186283 6 VPWR
port 613 nsew power input
rlabel locali s 298660 186283 298661 186391 6 VPWR
port 613 nsew power input
rlabel locali s 1259 185705 1340 185813 6 VPWR
port 613 nsew power input
rlabel locali s 1121 185813 1340 186031 6 VPWR
port 613 nsew power input
rlabel locali s 1104 186031 1340 186065 6 VPWR
port 613 nsew power input
rlabel locali s 1121 186065 1340 186283 6 VPWR
port 613 nsew power input
rlabel locali s 1259 186283 1340 186391 6 VPWR
port 613 nsew power input
rlabel locali s 298660 186793 298661 186901 6 VPWR
port 613 nsew power input
rlabel locali s 298660 186901 298799 187119 6 VPWR
port 613 nsew power input
rlabel locali s 298660 187119 298816 187153 6 VPWR
port 613 nsew power input
rlabel locali s 298660 187153 298799 187371 6 VPWR
port 613 nsew power input
rlabel locali s 298660 187371 298661 187479 6 VPWR
port 613 nsew power input
rlabel locali s 1259 186793 1340 186901 6 VPWR
port 613 nsew power input
rlabel locali s 1121 186901 1340 187119 6 VPWR
port 613 nsew power input
rlabel locali s 1104 187119 1340 187153 6 VPWR
port 613 nsew power input
rlabel locali s 1121 187153 1340 187371 6 VPWR
port 613 nsew power input
rlabel locali s 1259 187371 1340 187479 6 VPWR
port 613 nsew power input
rlabel locali s 298660 187881 298661 187989 6 VPWR
port 613 nsew power input
rlabel locali s 298660 187989 298799 188207 6 VPWR
port 613 nsew power input
rlabel locali s 298660 188207 298816 188241 6 VPWR
port 613 nsew power input
rlabel locali s 298660 188241 298799 188459 6 VPWR
port 613 nsew power input
rlabel locali s 298660 188459 298661 188567 6 VPWR
port 613 nsew power input
rlabel locali s 1259 187881 1340 187989 6 VPWR
port 613 nsew power input
rlabel locali s 1121 187989 1340 188207 6 VPWR
port 613 nsew power input
rlabel locali s 1104 188207 1340 188241 6 VPWR
port 613 nsew power input
rlabel locali s 1121 188241 1340 188459 6 VPWR
port 613 nsew power input
rlabel locali s 1259 188459 1340 188567 6 VPWR
port 613 nsew power input
rlabel locali s 298660 188969 298661 189077 6 VPWR
port 613 nsew power input
rlabel locali s 298660 189077 298799 189295 6 VPWR
port 613 nsew power input
rlabel locali s 298660 189295 298816 189329 6 VPWR
port 613 nsew power input
rlabel locali s 298660 189329 298799 189547 6 VPWR
port 613 nsew power input
rlabel locali s 298660 189547 298661 189655 6 VPWR
port 613 nsew power input
rlabel locali s 1259 188969 1340 189077 6 VPWR
port 613 nsew power input
rlabel locali s 1121 189077 1340 189295 6 VPWR
port 613 nsew power input
rlabel locali s 1104 189295 1340 189329 6 VPWR
port 613 nsew power input
rlabel locali s 1121 189329 1340 189547 6 VPWR
port 613 nsew power input
rlabel locali s 1259 189547 1340 189655 6 VPWR
port 613 nsew power input
rlabel locali s 298660 190057 298661 190165 6 VPWR
port 613 nsew power input
rlabel locali s 298660 190165 298799 190383 6 VPWR
port 613 nsew power input
rlabel locali s 298660 190383 298816 190417 6 VPWR
port 613 nsew power input
rlabel locali s 298660 190417 298799 190635 6 VPWR
port 613 nsew power input
rlabel locali s 298660 190635 298661 190743 6 VPWR
port 613 nsew power input
rlabel locali s 1259 190057 1340 190165 6 VPWR
port 613 nsew power input
rlabel locali s 1121 190165 1340 190383 6 VPWR
port 613 nsew power input
rlabel locali s 1104 190383 1340 190417 6 VPWR
port 613 nsew power input
rlabel locali s 1121 190417 1340 190635 6 VPWR
port 613 nsew power input
rlabel locali s 1259 190635 1340 190743 6 VPWR
port 613 nsew power input
rlabel locali s 298660 191145 298661 191253 6 VPWR
port 613 nsew power input
rlabel locali s 298660 191253 298799 191471 6 VPWR
port 613 nsew power input
rlabel locali s 298660 191471 298816 191505 6 VPWR
port 613 nsew power input
rlabel locali s 298660 191505 298799 191723 6 VPWR
port 613 nsew power input
rlabel locali s 298660 191723 298661 191831 6 VPWR
port 613 nsew power input
rlabel locali s 1259 191145 1340 191253 6 VPWR
port 613 nsew power input
rlabel locali s 1121 191253 1340 191471 6 VPWR
port 613 nsew power input
rlabel locali s 1104 191471 1340 191505 6 VPWR
port 613 nsew power input
rlabel locali s 1121 191505 1340 191723 6 VPWR
port 613 nsew power input
rlabel locali s 1259 191723 1340 191831 6 VPWR
port 613 nsew power input
rlabel locali s 298660 192233 298661 192341 6 VPWR
port 613 nsew power input
rlabel locali s 298660 192341 298799 192559 6 VPWR
port 613 nsew power input
rlabel locali s 298660 192559 298816 192593 6 VPWR
port 613 nsew power input
rlabel locali s 298660 192593 298799 192811 6 VPWR
port 613 nsew power input
rlabel locali s 298660 192811 298661 192919 6 VPWR
port 613 nsew power input
rlabel locali s 1259 192233 1340 192341 6 VPWR
port 613 nsew power input
rlabel locali s 1121 192341 1340 192559 6 VPWR
port 613 nsew power input
rlabel locali s 1104 192559 1340 192593 6 VPWR
port 613 nsew power input
rlabel locali s 1121 192593 1340 192811 6 VPWR
port 613 nsew power input
rlabel locali s 1259 192811 1340 192919 6 VPWR
port 613 nsew power input
rlabel locali s 298660 193321 298661 193429 6 VPWR
port 613 nsew power input
rlabel locali s 298660 193429 298799 193647 6 VPWR
port 613 nsew power input
rlabel locali s 298660 193647 298816 193681 6 VPWR
port 613 nsew power input
rlabel locali s 298660 193681 298799 193899 6 VPWR
port 613 nsew power input
rlabel locali s 298660 193899 298661 194007 6 VPWR
port 613 nsew power input
rlabel locali s 1259 193321 1340 193429 6 VPWR
port 613 nsew power input
rlabel locali s 1121 193429 1340 193647 6 VPWR
port 613 nsew power input
rlabel locali s 1104 193647 1340 193681 6 VPWR
port 613 nsew power input
rlabel locali s 1121 193681 1340 193899 6 VPWR
port 613 nsew power input
rlabel locali s 1259 193899 1340 194007 6 VPWR
port 613 nsew power input
rlabel locali s 298660 194409 298661 194517 6 VPWR
port 613 nsew power input
rlabel locali s 298660 194517 298799 194735 6 VPWR
port 613 nsew power input
rlabel locali s 298660 194735 298816 194769 6 VPWR
port 613 nsew power input
rlabel locali s 298660 194769 298799 194987 6 VPWR
port 613 nsew power input
rlabel locali s 298660 194987 298661 195095 6 VPWR
port 613 nsew power input
rlabel locali s 1259 194409 1340 194517 6 VPWR
port 613 nsew power input
rlabel locali s 1121 194517 1340 194735 6 VPWR
port 613 nsew power input
rlabel locali s 1104 194735 1340 194769 6 VPWR
port 613 nsew power input
rlabel locali s 1121 194769 1340 194987 6 VPWR
port 613 nsew power input
rlabel locali s 1259 194987 1340 195095 6 VPWR
port 613 nsew power input
rlabel locali s 298660 195497 298661 195605 6 VPWR
port 613 nsew power input
rlabel locali s 298660 195605 298799 195823 6 VPWR
port 613 nsew power input
rlabel locali s 298660 195823 298816 195857 6 VPWR
port 613 nsew power input
rlabel locali s 298660 195857 298799 196075 6 VPWR
port 613 nsew power input
rlabel locali s 298660 196075 298661 196183 6 VPWR
port 613 nsew power input
rlabel locali s 1259 195497 1340 195605 6 VPWR
port 613 nsew power input
rlabel locali s 1121 195605 1340 195823 6 VPWR
port 613 nsew power input
rlabel locali s 1104 195823 1340 195857 6 VPWR
port 613 nsew power input
rlabel locali s 1121 195857 1340 196075 6 VPWR
port 613 nsew power input
rlabel locali s 1259 196075 1340 196183 6 VPWR
port 613 nsew power input
rlabel locali s 298660 196585 298661 196693 6 VPWR
port 613 nsew power input
rlabel locali s 298660 196693 298799 196911 6 VPWR
port 613 nsew power input
rlabel locali s 298660 196911 298816 196945 6 VPWR
port 613 nsew power input
rlabel locali s 298660 196945 298799 197163 6 VPWR
port 613 nsew power input
rlabel locali s 298660 197163 298661 197271 6 VPWR
port 613 nsew power input
rlabel locali s 1259 196585 1340 196693 6 VPWR
port 613 nsew power input
rlabel locali s 1121 196693 1340 196911 6 VPWR
port 613 nsew power input
rlabel locali s 1104 196911 1340 196945 6 VPWR
port 613 nsew power input
rlabel locali s 1121 196945 1340 197163 6 VPWR
port 613 nsew power input
rlabel locali s 1259 197163 1340 197271 6 VPWR
port 613 nsew power input
rlabel locali s 298660 197673 298661 197781 6 VPWR
port 613 nsew power input
rlabel locali s 298660 197781 298799 197999 6 VPWR
port 613 nsew power input
rlabel locali s 298660 197999 298816 198033 6 VPWR
port 613 nsew power input
rlabel locali s 298660 198033 298799 198251 6 VPWR
port 613 nsew power input
rlabel locali s 298660 198251 298661 198359 6 VPWR
port 613 nsew power input
rlabel locali s 1259 197673 1340 197781 6 VPWR
port 613 nsew power input
rlabel locali s 1121 197781 1340 197999 6 VPWR
port 613 nsew power input
rlabel locali s 1104 197999 1340 198033 6 VPWR
port 613 nsew power input
rlabel locali s 1121 198033 1340 198251 6 VPWR
port 613 nsew power input
rlabel locali s 1259 198251 1340 198359 6 VPWR
port 613 nsew power input
rlabel locali s 298660 198761 298661 198869 6 VPWR
port 613 nsew power input
rlabel locali s 298660 198869 298799 199087 6 VPWR
port 613 nsew power input
rlabel locali s 298660 199087 298816 199121 6 VPWR
port 613 nsew power input
rlabel locali s 298660 199121 298799 199339 6 VPWR
port 613 nsew power input
rlabel locali s 298660 199339 298661 199447 6 VPWR
port 613 nsew power input
rlabel locali s 1259 198761 1340 198869 6 VPWR
port 613 nsew power input
rlabel locali s 1121 198869 1340 199087 6 VPWR
port 613 nsew power input
rlabel locali s 1104 199087 1340 199121 6 VPWR
port 613 nsew power input
rlabel locali s 1121 199121 1340 199339 6 VPWR
port 613 nsew power input
rlabel locali s 1259 199339 1340 199447 6 VPWR
port 613 nsew power input
rlabel locali s 298660 199849 298661 199957 6 VPWR
port 613 nsew power input
rlabel locali s 298660 199957 298799 200175 6 VPWR
port 613 nsew power input
rlabel locali s 298660 200175 298816 200209 6 VPWR
port 613 nsew power input
rlabel locali s 298660 200209 298799 200427 6 VPWR
port 613 nsew power input
rlabel locali s 298660 200427 298661 200535 6 VPWR
port 613 nsew power input
rlabel locali s 1259 199849 1340 199957 6 VPWR
port 613 nsew power input
rlabel locali s 1121 199957 1340 200175 6 VPWR
port 613 nsew power input
rlabel locali s 1104 200175 1340 200209 6 VPWR
port 613 nsew power input
rlabel locali s 1121 200209 1340 200427 6 VPWR
port 613 nsew power input
rlabel locali s 1259 200427 1340 200535 6 VPWR
port 613 nsew power input
rlabel locali s 298660 200937 298661 201045 6 VPWR
port 613 nsew power input
rlabel locali s 298660 201045 298799 201263 6 VPWR
port 613 nsew power input
rlabel locali s 298660 201263 298816 201297 6 VPWR
port 613 nsew power input
rlabel locali s 298660 201297 298799 201515 6 VPWR
port 613 nsew power input
rlabel locali s 298660 201515 298661 201623 6 VPWR
port 613 nsew power input
rlabel locali s 1259 200937 1340 201045 6 VPWR
port 613 nsew power input
rlabel locali s 1121 201045 1340 201263 6 VPWR
port 613 nsew power input
rlabel locali s 1104 201263 1340 201297 6 VPWR
port 613 nsew power input
rlabel locali s 1121 201297 1340 201515 6 VPWR
port 613 nsew power input
rlabel locali s 1259 201515 1340 201623 6 VPWR
port 613 nsew power input
rlabel locali s 298660 202025 298661 202133 6 VPWR
port 613 nsew power input
rlabel locali s 298660 202133 298799 202351 6 VPWR
port 613 nsew power input
rlabel locali s 298660 202351 298816 202385 6 VPWR
port 613 nsew power input
rlabel locali s 298660 202385 298799 202603 6 VPWR
port 613 nsew power input
rlabel locali s 298660 202603 298661 202711 6 VPWR
port 613 nsew power input
rlabel locali s 1259 202025 1340 202133 6 VPWR
port 613 nsew power input
rlabel locali s 1121 202133 1340 202351 6 VPWR
port 613 nsew power input
rlabel locali s 1104 202351 1340 202385 6 VPWR
port 613 nsew power input
rlabel locali s 1121 202385 1340 202603 6 VPWR
port 613 nsew power input
rlabel locali s 1259 202603 1340 202711 6 VPWR
port 613 nsew power input
rlabel locali s 298660 203113 298661 203221 6 VPWR
port 613 nsew power input
rlabel locali s 298660 203221 298799 203439 6 VPWR
port 613 nsew power input
rlabel locali s 298660 203439 298816 203473 6 VPWR
port 613 nsew power input
rlabel locali s 298660 203473 298799 203691 6 VPWR
port 613 nsew power input
rlabel locali s 298660 203691 298661 203799 6 VPWR
port 613 nsew power input
rlabel locali s 1259 203113 1340 203221 6 VPWR
port 613 nsew power input
rlabel locali s 1121 203221 1340 203439 6 VPWR
port 613 nsew power input
rlabel locali s 1104 203439 1340 203473 6 VPWR
port 613 nsew power input
rlabel locali s 1121 203473 1340 203691 6 VPWR
port 613 nsew power input
rlabel locali s 1259 203691 1340 203799 6 VPWR
port 613 nsew power input
rlabel locali s 298660 204201 298661 204309 6 VPWR
port 613 nsew power input
rlabel locali s 298660 204309 298799 204527 6 VPWR
port 613 nsew power input
rlabel locali s 298660 204527 298816 204561 6 VPWR
port 613 nsew power input
rlabel locali s 298660 204561 298799 204779 6 VPWR
port 613 nsew power input
rlabel locali s 298660 204779 298661 204887 6 VPWR
port 613 nsew power input
rlabel locali s 1259 204201 1340 204309 6 VPWR
port 613 nsew power input
rlabel locali s 1121 204309 1340 204527 6 VPWR
port 613 nsew power input
rlabel locali s 1104 204527 1340 204561 6 VPWR
port 613 nsew power input
rlabel locali s 1121 204561 1340 204779 6 VPWR
port 613 nsew power input
rlabel locali s 1259 204779 1340 204887 6 VPWR
port 613 nsew power input
rlabel locali s 298660 205289 298661 205397 6 VPWR
port 613 nsew power input
rlabel locali s 298660 205397 298799 205615 6 VPWR
port 613 nsew power input
rlabel locali s 298660 205615 298816 205649 6 VPWR
port 613 nsew power input
rlabel locali s 298660 205649 298799 205867 6 VPWR
port 613 nsew power input
rlabel locali s 298660 205867 298661 205975 6 VPWR
port 613 nsew power input
rlabel locali s 1259 205289 1340 205397 6 VPWR
port 613 nsew power input
rlabel locali s 1121 205397 1340 205615 6 VPWR
port 613 nsew power input
rlabel locali s 1104 205615 1340 205649 6 VPWR
port 613 nsew power input
rlabel locali s 1121 205649 1340 205867 6 VPWR
port 613 nsew power input
rlabel locali s 1259 205867 1340 205975 6 VPWR
port 613 nsew power input
rlabel locali s 298660 206377 298661 206485 6 VPWR
port 613 nsew power input
rlabel locali s 298660 206485 298799 206703 6 VPWR
port 613 nsew power input
rlabel locali s 298660 206703 298816 206737 6 VPWR
port 613 nsew power input
rlabel locali s 298660 206737 298799 206955 6 VPWR
port 613 nsew power input
rlabel locali s 298660 206955 298661 207063 6 VPWR
port 613 nsew power input
rlabel locali s 1259 206377 1340 206485 6 VPWR
port 613 nsew power input
rlabel locali s 1121 206485 1340 206703 6 VPWR
port 613 nsew power input
rlabel locali s 1104 206703 1340 206737 6 VPWR
port 613 nsew power input
rlabel locali s 1121 206737 1340 206955 6 VPWR
port 613 nsew power input
rlabel locali s 1259 206955 1340 207063 6 VPWR
port 613 nsew power input
rlabel locali s 298660 207465 298661 207573 6 VPWR
port 613 nsew power input
rlabel locali s 298660 207573 298799 207791 6 VPWR
port 613 nsew power input
rlabel locali s 298660 207791 298816 207825 6 VPWR
port 613 nsew power input
rlabel locali s 298660 207825 298799 208043 6 VPWR
port 613 nsew power input
rlabel locali s 298660 208043 298661 208151 6 VPWR
port 613 nsew power input
rlabel locali s 1259 207465 1340 207573 6 VPWR
port 613 nsew power input
rlabel locali s 1121 207573 1340 207791 6 VPWR
port 613 nsew power input
rlabel locali s 1104 207791 1340 207825 6 VPWR
port 613 nsew power input
rlabel locali s 1121 207825 1340 208043 6 VPWR
port 613 nsew power input
rlabel locali s 1259 208043 1340 208151 6 VPWR
port 613 nsew power input
rlabel locali s 298660 208553 298661 208661 6 VPWR
port 613 nsew power input
rlabel locali s 298660 208661 298799 208879 6 VPWR
port 613 nsew power input
rlabel locali s 298660 208879 298816 208913 6 VPWR
port 613 nsew power input
rlabel locali s 298660 208913 298799 209131 6 VPWR
port 613 nsew power input
rlabel locali s 298660 209131 298661 209239 6 VPWR
port 613 nsew power input
rlabel locali s 1259 208553 1340 208661 6 VPWR
port 613 nsew power input
rlabel locali s 1121 208661 1340 208879 6 VPWR
port 613 nsew power input
rlabel locali s 1104 208879 1340 208913 6 VPWR
port 613 nsew power input
rlabel locali s 1121 208913 1340 209131 6 VPWR
port 613 nsew power input
rlabel locali s 1259 209131 1340 209239 6 VPWR
port 613 nsew power input
rlabel locali s 298660 209641 298661 209749 6 VPWR
port 613 nsew power input
rlabel locali s 298660 209749 298799 209967 6 VPWR
port 613 nsew power input
rlabel locali s 298660 209967 298816 210001 6 VPWR
port 613 nsew power input
rlabel locali s 298660 210001 298799 210219 6 VPWR
port 613 nsew power input
rlabel locali s 298660 210219 298661 210327 6 VPWR
port 613 nsew power input
rlabel locali s 1259 209641 1340 209749 6 VPWR
port 613 nsew power input
rlabel locali s 1121 209749 1340 209967 6 VPWR
port 613 nsew power input
rlabel locali s 1104 209967 1340 210001 6 VPWR
port 613 nsew power input
rlabel locali s 1121 210001 1340 210219 6 VPWR
port 613 nsew power input
rlabel locali s 1259 210219 1340 210327 6 VPWR
port 613 nsew power input
rlabel locali s 298660 210729 298661 210837 6 VPWR
port 613 nsew power input
rlabel locali s 298660 210837 298799 211055 6 VPWR
port 613 nsew power input
rlabel locali s 298660 211055 298816 211089 6 VPWR
port 613 nsew power input
rlabel locali s 298660 211089 298799 211307 6 VPWR
port 613 nsew power input
rlabel locali s 298660 211307 298661 211415 6 VPWR
port 613 nsew power input
rlabel locali s 1259 210729 1340 210837 6 VPWR
port 613 nsew power input
rlabel locali s 1121 210837 1340 211055 6 VPWR
port 613 nsew power input
rlabel locali s 1104 211055 1340 211089 6 VPWR
port 613 nsew power input
rlabel locali s 1121 211089 1340 211307 6 VPWR
port 613 nsew power input
rlabel locali s 1259 211307 1340 211415 6 VPWR
port 613 nsew power input
rlabel locali s 298660 211817 298661 211925 6 VPWR
port 613 nsew power input
rlabel locali s 298660 211925 298799 212143 6 VPWR
port 613 nsew power input
rlabel locali s 298660 212143 298816 212177 6 VPWR
port 613 nsew power input
rlabel locali s 298660 212177 298799 212395 6 VPWR
port 613 nsew power input
rlabel locali s 298660 212395 298661 212503 6 VPWR
port 613 nsew power input
rlabel locali s 1259 211817 1340 211925 6 VPWR
port 613 nsew power input
rlabel locali s 1121 211925 1340 212143 6 VPWR
port 613 nsew power input
rlabel locali s 1104 212143 1340 212177 6 VPWR
port 613 nsew power input
rlabel locali s 1121 212177 1340 212395 6 VPWR
port 613 nsew power input
rlabel locali s 1259 212395 1340 212503 6 VPWR
port 613 nsew power input
rlabel locali s 298660 212905 298661 213013 6 VPWR
port 613 nsew power input
rlabel locali s 298660 213013 298799 213231 6 VPWR
port 613 nsew power input
rlabel locali s 298660 213231 298816 213265 6 VPWR
port 613 nsew power input
rlabel locali s 298660 213265 298799 213483 6 VPWR
port 613 nsew power input
rlabel locali s 298660 213483 298661 213591 6 VPWR
port 613 nsew power input
rlabel locali s 1259 212905 1340 213013 6 VPWR
port 613 nsew power input
rlabel locali s 1121 213013 1340 213231 6 VPWR
port 613 nsew power input
rlabel locali s 1104 213231 1340 213265 6 VPWR
port 613 nsew power input
rlabel locali s 1121 213265 1340 213483 6 VPWR
port 613 nsew power input
rlabel locali s 1259 213483 1340 213591 6 VPWR
port 613 nsew power input
rlabel locali s 298660 213993 298661 214101 6 VPWR
port 613 nsew power input
rlabel locali s 298660 214101 298799 214319 6 VPWR
port 613 nsew power input
rlabel locali s 298660 214319 298816 214353 6 VPWR
port 613 nsew power input
rlabel locali s 298660 214353 298799 214571 6 VPWR
port 613 nsew power input
rlabel locali s 298660 214571 298661 214679 6 VPWR
port 613 nsew power input
rlabel locali s 1259 213993 1340 214101 6 VPWR
port 613 nsew power input
rlabel locali s 1121 214101 1340 214319 6 VPWR
port 613 nsew power input
rlabel locali s 1104 214319 1340 214353 6 VPWR
port 613 nsew power input
rlabel locali s 1121 214353 1340 214571 6 VPWR
port 613 nsew power input
rlabel locali s 1259 214571 1340 214679 6 VPWR
port 613 nsew power input
rlabel locali s 298660 215081 298661 215189 6 VPWR
port 613 nsew power input
rlabel locali s 298660 215189 298799 215407 6 VPWR
port 613 nsew power input
rlabel locali s 298660 215407 298816 215441 6 VPWR
port 613 nsew power input
rlabel locali s 298660 215441 298799 215659 6 VPWR
port 613 nsew power input
rlabel locali s 298660 215659 298661 215767 6 VPWR
port 613 nsew power input
rlabel locali s 1259 215081 1340 215189 6 VPWR
port 613 nsew power input
rlabel locali s 1121 215189 1340 215407 6 VPWR
port 613 nsew power input
rlabel locali s 1104 215407 1340 215441 6 VPWR
port 613 nsew power input
rlabel locali s 1121 215441 1340 215659 6 VPWR
port 613 nsew power input
rlabel locali s 1259 215659 1340 215767 6 VPWR
port 613 nsew power input
rlabel locali s 298660 216169 298661 216277 6 VPWR
port 613 nsew power input
rlabel locali s 298660 216277 298799 216495 6 VPWR
port 613 nsew power input
rlabel locali s 298660 216495 298816 216529 6 VPWR
port 613 nsew power input
rlabel locali s 298660 216529 298799 216747 6 VPWR
port 613 nsew power input
rlabel locali s 298660 216747 298661 216855 6 VPWR
port 613 nsew power input
rlabel locali s 1259 216169 1340 216277 6 VPWR
port 613 nsew power input
rlabel locali s 1121 216277 1340 216495 6 VPWR
port 613 nsew power input
rlabel locali s 1104 216495 1340 216529 6 VPWR
port 613 nsew power input
rlabel locali s 1121 216529 1340 216747 6 VPWR
port 613 nsew power input
rlabel locali s 1259 216747 1340 216855 6 VPWR
port 613 nsew power input
rlabel locali s 298660 217257 298661 217365 6 VPWR
port 613 nsew power input
rlabel locali s 298660 217365 298799 217583 6 VPWR
port 613 nsew power input
rlabel locali s 298660 217583 298816 217617 6 VPWR
port 613 nsew power input
rlabel locali s 298660 217617 298799 217835 6 VPWR
port 613 nsew power input
rlabel locali s 298660 217835 298661 217943 6 VPWR
port 613 nsew power input
rlabel locali s 1259 217257 1340 217365 6 VPWR
port 613 nsew power input
rlabel locali s 1121 217365 1340 217583 6 VPWR
port 613 nsew power input
rlabel locali s 1104 217583 1340 217617 6 VPWR
port 613 nsew power input
rlabel locali s 1121 217617 1340 217835 6 VPWR
port 613 nsew power input
rlabel locali s 1259 217835 1340 217943 6 VPWR
port 613 nsew power input
rlabel locali s 298660 218345 298661 218453 6 VPWR
port 613 nsew power input
rlabel locali s 298660 218453 298799 218671 6 VPWR
port 613 nsew power input
rlabel locali s 298660 218671 298816 218705 6 VPWR
port 613 nsew power input
rlabel locali s 298660 218705 298799 218923 6 VPWR
port 613 nsew power input
rlabel locali s 298660 218923 298661 219031 6 VPWR
port 613 nsew power input
rlabel locali s 1259 218345 1340 218453 6 VPWR
port 613 nsew power input
rlabel locali s 1121 218453 1340 218671 6 VPWR
port 613 nsew power input
rlabel locali s 1104 218671 1340 218705 6 VPWR
port 613 nsew power input
rlabel locali s 1121 218705 1340 218923 6 VPWR
port 613 nsew power input
rlabel locali s 1259 218923 1340 219031 6 VPWR
port 613 nsew power input
rlabel locali s 298660 219433 298661 219541 6 VPWR
port 613 nsew power input
rlabel locali s 298660 219541 298799 219759 6 VPWR
port 613 nsew power input
rlabel locali s 298660 219759 298816 219793 6 VPWR
port 613 nsew power input
rlabel locali s 298660 219793 298799 220011 6 VPWR
port 613 nsew power input
rlabel locali s 298660 220011 298661 220119 6 VPWR
port 613 nsew power input
rlabel locali s 1259 219433 1340 219541 6 VPWR
port 613 nsew power input
rlabel locali s 1121 219541 1340 219759 6 VPWR
port 613 nsew power input
rlabel locali s 1104 219759 1340 219793 6 VPWR
port 613 nsew power input
rlabel locali s 1121 219793 1340 220011 6 VPWR
port 613 nsew power input
rlabel locali s 1259 220011 1340 220119 6 VPWR
port 613 nsew power input
rlabel locali s 298660 220521 298661 220629 6 VPWR
port 613 nsew power input
rlabel locali s 298660 220629 298799 220847 6 VPWR
port 613 nsew power input
rlabel locali s 298660 220847 298816 220881 6 VPWR
port 613 nsew power input
rlabel locali s 298660 220881 298799 221099 6 VPWR
port 613 nsew power input
rlabel locali s 298660 221099 298661 221207 6 VPWR
port 613 nsew power input
rlabel locali s 1259 220521 1340 220629 6 VPWR
port 613 nsew power input
rlabel locali s 1121 220629 1340 220847 6 VPWR
port 613 nsew power input
rlabel locali s 1104 220847 1340 220881 6 VPWR
port 613 nsew power input
rlabel locali s 1121 220881 1340 221099 6 VPWR
port 613 nsew power input
rlabel locali s 1259 221099 1340 221207 6 VPWR
port 613 nsew power input
rlabel locali s 298660 221609 298661 221717 6 VPWR
port 613 nsew power input
rlabel locali s 298660 221717 298799 221935 6 VPWR
port 613 nsew power input
rlabel locali s 298660 221935 298816 221969 6 VPWR
port 613 nsew power input
rlabel locali s 298660 221969 298799 222187 6 VPWR
port 613 nsew power input
rlabel locali s 298660 222187 298661 222295 6 VPWR
port 613 nsew power input
rlabel locali s 1259 221609 1340 221717 6 VPWR
port 613 nsew power input
rlabel locali s 1121 221717 1340 221935 6 VPWR
port 613 nsew power input
rlabel locali s 1104 221935 1340 221969 6 VPWR
port 613 nsew power input
rlabel locali s 1121 221969 1340 222187 6 VPWR
port 613 nsew power input
rlabel locali s 1259 222187 1340 222295 6 VPWR
port 613 nsew power input
rlabel locali s 298660 222697 298661 222805 6 VPWR
port 613 nsew power input
rlabel locali s 298660 222805 298799 223023 6 VPWR
port 613 nsew power input
rlabel locali s 298660 223023 298816 223057 6 VPWR
port 613 nsew power input
rlabel locali s 298660 223057 298799 223275 6 VPWR
port 613 nsew power input
rlabel locali s 298660 223275 298661 223383 6 VPWR
port 613 nsew power input
rlabel locali s 1259 222697 1340 222805 6 VPWR
port 613 nsew power input
rlabel locali s 1121 222805 1340 223023 6 VPWR
port 613 nsew power input
rlabel locali s 1104 223023 1340 223057 6 VPWR
port 613 nsew power input
rlabel locali s 1121 223057 1340 223275 6 VPWR
port 613 nsew power input
rlabel locali s 1259 223275 1340 223383 6 VPWR
port 613 nsew power input
rlabel locali s 298660 223785 298661 223893 6 VPWR
port 613 nsew power input
rlabel locali s 298660 223893 298799 224111 6 VPWR
port 613 nsew power input
rlabel locali s 298660 224111 298816 224145 6 VPWR
port 613 nsew power input
rlabel locali s 298660 224145 298799 224363 6 VPWR
port 613 nsew power input
rlabel locali s 298660 224363 298661 224471 6 VPWR
port 613 nsew power input
rlabel locali s 1259 223785 1340 223893 6 VPWR
port 613 nsew power input
rlabel locali s 1121 223893 1340 224111 6 VPWR
port 613 nsew power input
rlabel locali s 1104 224111 1340 224145 6 VPWR
port 613 nsew power input
rlabel locali s 1121 224145 1340 224363 6 VPWR
port 613 nsew power input
rlabel locali s 1259 224363 1340 224471 6 VPWR
port 613 nsew power input
rlabel locali s 298660 224873 298661 224981 6 VPWR
port 613 nsew power input
rlabel locali s 298660 224981 298799 225199 6 VPWR
port 613 nsew power input
rlabel locali s 298660 225199 298816 225233 6 VPWR
port 613 nsew power input
rlabel locali s 298660 225233 298799 225451 6 VPWR
port 613 nsew power input
rlabel locali s 298660 225451 298661 225559 6 VPWR
port 613 nsew power input
rlabel locali s 1259 224873 1340 224981 6 VPWR
port 613 nsew power input
rlabel locali s 1121 224981 1340 225199 6 VPWR
port 613 nsew power input
rlabel locali s 1104 225199 1340 225233 6 VPWR
port 613 nsew power input
rlabel locali s 1121 225233 1340 225451 6 VPWR
port 613 nsew power input
rlabel locali s 1259 225451 1340 225559 6 VPWR
port 613 nsew power input
rlabel locali s 298660 225961 298661 226069 6 VPWR
port 613 nsew power input
rlabel locali s 298660 226069 298799 226287 6 VPWR
port 613 nsew power input
rlabel locali s 298660 226287 298816 226321 6 VPWR
port 613 nsew power input
rlabel locali s 298660 226321 298799 226539 6 VPWR
port 613 nsew power input
rlabel locali s 298660 226539 298661 226647 6 VPWR
port 613 nsew power input
rlabel locali s 1259 225961 1340 226069 6 VPWR
port 613 nsew power input
rlabel locali s 1121 226069 1340 226287 6 VPWR
port 613 nsew power input
rlabel locali s 1104 226287 1340 226321 6 VPWR
port 613 nsew power input
rlabel locali s 1121 226321 1340 226539 6 VPWR
port 613 nsew power input
rlabel locali s 1259 226539 1340 226647 6 VPWR
port 613 nsew power input
rlabel locali s 298660 227049 298661 227157 6 VPWR
port 613 nsew power input
rlabel locali s 298660 227157 298799 227375 6 VPWR
port 613 nsew power input
rlabel locali s 298660 227375 298816 227409 6 VPWR
port 613 nsew power input
rlabel locali s 298660 227409 298799 227627 6 VPWR
port 613 nsew power input
rlabel locali s 298660 227627 298661 227735 6 VPWR
port 613 nsew power input
rlabel locali s 1259 227049 1340 227157 6 VPWR
port 613 nsew power input
rlabel locali s 1121 227157 1340 227375 6 VPWR
port 613 nsew power input
rlabel locali s 1104 227375 1340 227409 6 VPWR
port 613 nsew power input
rlabel locali s 1121 227409 1340 227627 6 VPWR
port 613 nsew power input
rlabel locali s 1259 227627 1340 227735 6 VPWR
port 613 nsew power input
rlabel locali s 298660 228137 298661 228245 6 VPWR
port 613 nsew power input
rlabel locali s 298660 228245 298799 228463 6 VPWR
port 613 nsew power input
rlabel locali s 298660 228463 298816 228497 6 VPWR
port 613 nsew power input
rlabel locali s 298660 228497 298799 228715 6 VPWR
port 613 nsew power input
rlabel locali s 298660 228715 298661 228823 6 VPWR
port 613 nsew power input
rlabel locali s 1259 228137 1340 228245 6 VPWR
port 613 nsew power input
rlabel locali s 1121 228245 1340 228463 6 VPWR
port 613 nsew power input
rlabel locali s 1104 228463 1340 228497 6 VPWR
port 613 nsew power input
rlabel locali s 1121 228497 1340 228715 6 VPWR
port 613 nsew power input
rlabel locali s 1259 228715 1340 228823 6 VPWR
port 613 nsew power input
rlabel locali s 298660 229225 298661 229333 6 VPWR
port 613 nsew power input
rlabel locali s 298660 229333 298799 229551 6 VPWR
port 613 nsew power input
rlabel locali s 298660 229551 298816 229585 6 VPWR
port 613 nsew power input
rlabel locali s 298660 229585 298799 229803 6 VPWR
port 613 nsew power input
rlabel locali s 298660 229803 298661 229911 6 VPWR
port 613 nsew power input
rlabel locali s 1259 229225 1340 229333 6 VPWR
port 613 nsew power input
rlabel locali s 1121 229333 1340 229551 6 VPWR
port 613 nsew power input
rlabel locali s 1104 229551 1340 229585 6 VPWR
port 613 nsew power input
rlabel locali s 1121 229585 1340 229803 6 VPWR
port 613 nsew power input
rlabel locali s 1259 229803 1340 229911 6 VPWR
port 613 nsew power input
rlabel locali s 298660 230313 298661 230421 6 VPWR
port 613 nsew power input
rlabel locali s 298660 230421 298799 230639 6 VPWR
port 613 nsew power input
rlabel locali s 298660 230639 298816 230673 6 VPWR
port 613 nsew power input
rlabel locali s 298660 230673 298799 230891 6 VPWR
port 613 nsew power input
rlabel locali s 298660 230891 298661 230999 6 VPWR
port 613 nsew power input
rlabel locali s 1259 230313 1340 230421 6 VPWR
port 613 nsew power input
rlabel locali s 1121 230421 1340 230639 6 VPWR
port 613 nsew power input
rlabel locali s 1104 230639 1340 230673 6 VPWR
port 613 nsew power input
rlabel locali s 1121 230673 1340 230891 6 VPWR
port 613 nsew power input
rlabel locali s 1259 230891 1340 230999 6 VPWR
port 613 nsew power input
rlabel locali s 298660 231401 298661 231509 6 VPWR
port 613 nsew power input
rlabel locali s 298660 231509 298799 231727 6 VPWR
port 613 nsew power input
rlabel locali s 298660 231727 298816 231761 6 VPWR
port 613 nsew power input
rlabel locali s 298660 231761 298799 231979 6 VPWR
port 613 nsew power input
rlabel locali s 298660 231979 298661 232087 6 VPWR
port 613 nsew power input
rlabel locali s 1259 231401 1340 231509 6 VPWR
port 613 nsew power input
rlabel locali s 1121 231509 1340 231727 6 VPWR
port 613 nsew power input
rlabel locali s 1104 231727 1340 231761 6 VPWR
port 613 nsew power input
rlabel locali s 1121 231761 1340 231979 6 VPWR
port 613 nsew power input
rlabel locali s 1259 231979 1340 232087 6 VPWR
port 613 nsew power input
rlabel locali s 298660 232489 298661 232597 6 VPWR
port 613 nsew power input
rlabel locali s 298660 232597 298799 232815 6 VPWR
port 613 nsew power input
rlabel locali s 298660 232815 298816 232849 6 VPWR
port 613 nsew power input
rlabel locali s 298660 232849 298799 233067 6 VPWR
port 613 nsew power input
rlabel locali s 298660 233067 298661 233175 6 VPWR
port 613 nsew power input
rlabel locali s 1259 232489 1340 232597 6 VPWR
port 613 nsew power input
rlabel locali s 1121 232597 1340 232815 6 VPWR
port 613 nsew power input
rlabel locali s 1104 232815 1340 232849 6 VPWR
port 613 nsew power input
rlabel locali s 1121 232849 1340 233067 6 VPWR
port 613 nsew power input
rlabel locali s 1259 233067 1340 233175 6 VPWR
port 613 nsew power input
rlabel locali s 298660 233577 298661 233685 6 VPWR
port 613 nsew power input
rlabel locali s 298660 233685 298799 233903 6 VPWR
port 613 nsew power input
rlabel locali s 298660 233903 298816 233937 6 VPWR
port 613 nsew power input
rlabel locali s 298660 233937 298799 234155 6 VPWR
port 613 nsew power input
rlabel locali s 298660 234155 298661 234263 6 VPWR
port 613 nsew power input
rlabel locali s 1259 233577 1340 233685 6 VPWR
port 613 nsew power input
rlabel locali s 1121 233685 1340 233903 6 VPWR
port 613 nsew power input
rlabel locali s 1104 233903 1340 233937 6 VPWR
port 613 nsew power input
rlabel locali s 1121 233937 1340 234155 6 VPWR
port 613 nsew power input
rlabel locali s 1259 234155 1340 234263 6 VPWR
port 613 nsew power input
rlabel locali s 298660 234665 298661 234773 6 VPWR
port 613 nsew power input
rlabel locali s 298660 234773 298799 234991 6 VPWR
port 613 nsew power input
rlabel locali s 298660 234991 298816 235025 6 VPWR
port 613 nsew power input
rlabel locali s 298660 235025 298799 235243 6 VPWR
port 613 nsew power input
rlabel locali s 298660 235243 298661 235351 6 VPWR
port 613 nsew power input
rlabel locali s 1259 234665 1340 234773 6 VPWR
port 613 nsew power input
rlabel locali s 1121 234773 1340 234991 6 VPWR
port 613 nsew power input
rlabel locali s 1104 234991 1340 235025 6 VPWR
port 613 nsew power input
rlabel locali s 1121 235025 1340 235243 6 VPWR
port 613 nsew power input
rlabel locali s 1259 235243 1340 235351 6 VPWR
port 613 nsew power input
rlabel locali s 298660 235753 298661 235861 6 VPWR
port 613 nsew power input
rlabel locali s 298660 235861 298799 236079 6 VPWR
port 613 nsew power input
rlabel locali s 298660 236079 298816 236113 6 VPWR
port 613 nsew power input
rlabel locali s 298660 236113 298799 236331 6 VPWR
port 613 nsew power input
rlabel locali s 298660 236331 298661 236439 6 VPWR
port 613 nsew power input
rlabel locali s 1259 235753 1340 235861 6 VPWR
port 613 nsew power input
rlabel locali s 1121 235861 1340 236079 6 VPWR
port 613 nsew power input
rlabel locali s 1104 236079 1340 236113 6 VPWR
port 613 nsew power input
rlabel locali s 1121 236113 1340 236331 6 VPWR
port 613 nsew power input
rlabel locali s 1259 236331 1340 236439 6 VPWR
port 613 nsew power input
rlabel locali s 298660 236841 298661 236949 6 VPWR
port 613 nsew power input
rlabel locali s 298660 236949 298799 237167 6 VPWR
port 613 nsew power input
rlabel locali s 298660 237167 298816 237201 6 VPWR
port 613 nsew power input
rlabel locali s 298660 237201 298799 237419 6 VPWR
port 613 nsew power input
rlabel locali s 298660 237419 298661 237527 6 VPWR
port 613 nsew power input
rlabel locali s 1259 236841 1340 236949 6 VPWR
port 613 nsew power input
rlabel locali s 1121 236949 1340 237167 6 VPWR
port 613 nsew power input
rlabel locali s 1104 237167 1340 237201 6 VPWR
port 613 nsew power input
rlabel locali s 1121 237201 1340 237419 6 VPWR
port 613 nsew power input
rlabel locali s 1259 237419 1340 237527 6 VPWR
port 613 nsew power input
rlabel locali s 298660 237929 298661 238037 6 VPWR
port 613 nsew power input
rlabel locali s 298660 238037 298799 238255 6 VPWR
port 613 nsew power input
rlabel locali s 298660 238255 298816 238289 6 VPWR
port 613 nsew power input
rlabel locali s 298660 238289 298799 238507 6 VPWR
port 613 nsew power input
rlabel locali s 298660 238507 298661 238615 6 VPWR
port 613 nsew power input
rlabel locali s 1259 237929 1340 238037 6 VPWR
port 613 nsew power input
rlabel locali s 1121 238037 1340 238255 6 VPWR
port 613 nsew power input
rlabel locali s 1104 238255 1340 238289 6 VPWR
port 613 nsew power input
rlabel locali s 1121 238289 1340 238507 6 VPWR
port 613 nsew power input
rlabel locali s 1259 238507 1340 238615 6 VPWR
port 613 nsew power input
rlabel locali s 298660 239017 298661 239125 6 VPWR
port 613 nsew power input
rlabel locali s 298660 239125 298799 239343 6 VPWR
port 613 nsew power input
rlabel locali s 298660 239343 298816 239377 6 VPWR
port 613 nsew power input
rlabel locali s 298660 239377 298799 239595 6 VPWR
port 613 nsew power input
rlabel locali s 298660 239595 298661 239703 6 VPWR
port 613 nsew power input
rlabel locali s 1259 239017 1340 239125 6 VPWR
port 613 nsew power input
rlabel locali s 1121 239125 1340 239343 6 VPWR
port 613 nsew power input
rlabel locali s 1104 239343 1340 239377 6 VPWR
port 613 nsew power input
rlabel locali s 1121 239377 1340 239595 6 VPWR
port 613 nsew power input
rlabel locali s 1259 239595 1340 239703 6 VPWR
port 613 nsew power input
rlabel locali s 298660 240105 298661 240213 6 VPWR
port 613 nsew power input
rlabel locali s 298660 240213 298799 240431 6 VPWR
port 613 nsew power input
rlabel locali s 298660 240431 298816 240465 6 VPWR
port 613 nsew power input
rlabel locali s 298660 240465 298799 240683 6 VPWR
port 613 nsew power input
rlabel locali s 298660 240683 298661 240791 6 VPWR
port 613 nsew power input
rlabel locali s 1259 240105 1340 240213 6 VPWR
port 613 nsew power input
rlabel locali s 1121 240213 1340 240431 6 VPWR
port 613 nsew power input
rlabel locali s 1104 240431 1340 240465 6 VPWR
port 613 nsew power input
rlabel locali s 1121 240465 1340 240683 6 VPWR
port 613 nsew power input
rlabel locali s 1259 240683 1340 240791 6 VPWR
port 613 nsew power input
rlabel locali s 298660 241193 298661 241301 6 VPWR
port 613 nsew power input
rlabel locali s 298660 241301 298799 241519 6 VPWR
port 613 nsew power input
rlabel locali s 298660 241519 298816 241553 6 VPWR
port 613 nsew power input
rlabel locali s 298660 241553 298799 241771 6 VPWR
port 613 nsew power input
rlabel locali s 298660 241771 298661 241879 6 VPWR
port 613 nsew power input
rlabel locali s 1259 241193 1340 241301 6 VPWR
port 613 nsew power input
rlabel locali s 1121 241301 1340 241519 6 VPWR
port 613 nsew power input
rlabel locali s 1104 241519 1340 241553 6 VPWR
port 613 nsew power input
rlabel locali s 1121 241553 1340 241771 6 VPWR
port 613 nsew power input
rlabel locali s 1259 241771 1340 241879 6 VPWR
port 613 nsew power input
rlabel locali s 298660 242281 298661 242389 6 VPWR
port 613 nsew power input
rlabel locali s 298660 242389 298799 242607 6 VPWR
port 613 nsew power input
rlabel locali s 298660 242607 298816 242641 6 VPWR
port 613 nsew power input
rlabel locali s 298660 242641 298799 242859 6 VPWR
port 613 nsew power input
rlabel locali s 298660 242859 298661 242967 6 VPWR
port 613 nsew power input
rlabel locali s 1259 242281 1340 242389 6 VPWR
port 613 nsew power input
rlabel locali s 1121 242389 1340 242607 6 VPWR
port 613 nsew power input
rlabel locali s 1104 242607 1340 242641 6 VPWR
port 613 nsew power input
rlabel locali s 1121 242641 1340 242859 6 VPWR
port 613 nsew power input
rlabel locali s 1259 242859 1340 242967 6 VPWR
port 613 nsew power input
rlabel locali s 298660 243369 298661 243477 6 VPWR
port 613 nsew power input
rlabel locali s 298660 243477 298799 243695 6 VPWR
port 613 nsew power input
rlabel locali s 298660 243695 298816 243729 6 VPWR
port 613 nsew power input
rlabel locali s 298660 243729 298799 243947 6 VPWR
port 613 nsew power input
rlabel locali s 298660 243947 298661 244055 6 VPWR
port 613 nsew power input
rlabel locali s 1259 243369 1340 243477 6 VPWR
port 613 nsew power input
rlabel locali s 1121 243477 1340 243695 6 VPWR
port 613 nsew power input
rlabel locali s 1104 243695 1340 243729 6 VPWR
port 613 nsew power input
rlabel locali s 1121 243729 1340 243947 6 VPWR
port 613 nsew power input
rlabel locali s 1259 243947 1340 244055 6 VPWR
port 613 nsew power input
rlabel locali s 298660 244457 298661 244565 6 VPWR
port 613 nsew power input
rlabel locali s 298660 244565 298799 244783 6 VPWR
port 613 nsew power input
rlabel locali s 298660 244783 298816 244817 6 VPWR
port 613 nsew power input
rlabel locali s 298660 244817 298799 245035 6 VPWR
port 613 nsew power input
rlabel locali s 298660 245035 298661 245143 6 VPWR
port 613 nsew power input
rlabel locali s 1259 244457 1340 244565 6 VPWR
port 613 nsew power input
rlabel locali s 1121 244565 1340 244783 6 VPWR
port 613 nsew power input
rlabel locali s 1104 244783 1340 244817 6 VPWR
port 613 nsew power input
rlabel locali s 1121 244817 1340 245035 6 VPWR
port 613 nsew power input
rlabel locali s 1259 245035 1340 245143 6 VPWR
port 613 nsew power input
rlabel locali s 298660 245545 298661 245653 6 VPWR
port 613 nsew power input
rlabel locali s 298660 245653 298799 245871 6 VPWR
port 613 nsew power input
rlabel locali s 298660 245871 298816 245905 6 VPWR
port 613 nsew power input
rlabel locali s 298660 245905 298799 246123 6 VPWR
port 613 nsew power input
rlabel locali s 298660 246123 298661 246231 6 VPWR
port 613 nsew power input
rlabel locali s 1259 245545 1340 245653 6 VPWR
port 613 nsew power input
rlabel locali s 1121 245653 1340 245871 6 VPWR
port 613 nsew power input
rlabel locali s 1104 245871 1340 245905 6 VPWR
port 613 nsew power input
rlabel locali s 1121 245905 1340 246123 6 VPWR
port 613 nsew power input
rlabel locali s 1259 246123 1340 246231 6 VPWR
port 613 nsew power input
rlabel locali s 298660 246633 298661 246741 6 VPWR
port 613 nsew power input
rlabel locali s 298660 246741 298799 246959 6 VPWR
port 613 nsew power input
rlabel locali s 298660 246959 298816 246993 6 VPWR
port 613 nsew power input
rlabel locali s 298660 246993 298799 247211 6 VPWR
port 613 nsew power input
rlabel locali s 298660 247211 298661 247319 6 VPWR
port 613 nsew power input
rlabel locali s 1259 246633 1340 246741 6 VPWR
port 613 nsew power input
rlabel locali s 1121 246741 1340 246959 6 VPWR
port 613 nsew power input
rlabel locali s 1104 246959 1340 246993 6 VPWR
port 613 nsew power input
rlabel locali s 1121 246993 1340 247211 6 VPWR
port 613 nsew power input
rlabel locali s 1259 247211 1340 247319 6 VPWR
port 613 nsew power input
rlabel locali s 298660 247721 298661 247829 6 VPWR
port 613 nsew power input
rlabel locali s 298660 247829 298799 248047 6 VPWR
port 613 nsew power input
rlabel locali s 298660 248047 298816 248081 6 VPWR
port 613 nsew power input
rlabel locali s 298660 248081 298799 248299 6 VPWR
port 613 nsew power input
rlabel locali s 298660 248299 298661 248407 6 VPWR
port 613 nsew power input
rlabel locali s 1259 247721 1340 247829 6 VPWR
port 613 nsew power input
rlabel locali s 1121 247829 1340 248047 6 VPWR
port 613 nsew power input
rlabel locali s 1104 248047 1340 248081 6 VPWR
port 613 nsew power input
rlabel locali s 1121 248081 1340 248299 6 VPWR
port 613 nsew power input
rlabel locali s 1259 248299 1340 248407 6 VPWR
port 613 nsew power input
rlabel locali s 298660 248809 298661 248917 6 VPWR
port 613 nsew power input
rlabel locali s 298660 248917 298799 249135 6 VPWR
port 613 nsew power input
rlabel locali s 298660 249135 298816 249169 6 VPWR
port 613 nsew power input
rlabel locali s 298660 249169 298799 249387 6 VPWR
port 613 nsew power input
rlabel locali s 298660 249387 298661 249495 6 VPWR
port 613 nsew power input
rlabel locali s 1259 248809 1340 248917 6 VPWR
port 613 nsew power input
rlabel locali s 1121 248917 1340 249135 6 VPWR
port 613 nsew power input
rlabel locali s 1104 249135 1340 249169 6 VPWR
port 613 nsew power input
rlabel locali s 1121 249169 1340 249387 6 VPWR
port 613 nsew power input
rlabel locali s 1259 249387 1340 249495 6 VPWR
port 613 nsew power input
rlabel locali s 298660 249897 298661 250005 6 VPWR
port 613 nsew power input
rlabel locali s 298660 250005 298799 250223 6 VPWR
port 613 nsew power input
rlabel locali s 298660 250223 298816 250257 6 VPWR
port 613 nsew power input
rlabel locali s 298660 250257 298799 250475 6 VPWR
port 613 nsew power input
rlabel locali s 298660 250475 298661 250583 6 VPWR
port 613 nsew power input
rlabel locali s 1259 249897 1340 250005 6 VPWR
port 613 nsew power input
rlabel locali s 1121 250005 1340 250223 6 VPWR
port 613 nsew power input
rlabel locali s 1104 250223 1340 250257 6 VPWR
port 613 nsew power input
rlabel locali s 1121 250257 1340 250475 6 VPWR
port 613 nsew power input
rlabel locali s 1259 250475 1340 250583 6 VPWR
port 613 nsew power input
rlabel locali s 298660 250985 298661 251093 6 VPWR
port 613 nsew power input
rlabel locali s 298660 251093 298799 251311 6 VPWR
port 613 nsew power input
rlabel locali s 298660 251311 298816 251345 6 VPWR
port 613 nsew power input
rlabel locali s 298660 251345 298799 251563 6 VPWR
port 613 nsew power input
rlabel locali s 298660 251563 298661 251671 6 VPWR
port 613 nsew power input
rlabel locali s 1259 250985 1340 251093 6 VPWR
port 613 nsew power input
rlabel locali s 1121 251093 1340 251311 6 VPWR
port 613 nsew power input
rlabel locali s 1104 251311 1340 251345 6 VPWR
port 613 nsew power input
rlabel locali s 1121 251345 1340 251563 6 VPWR
port 613 nsew power input
rlabel locali s 1259 251563 1340 251671 6 VPWR
port 613 nsew power input
rlabel locali s 298660 252073 298661 252181 6 VPWR
port 613 nsew power input
rlabel locali s 298660 252181 298799 252399 6 VPWR
port 613 nsew power input
rlabel locali s 298660 252399 298816 252433 6 VPWR
port 613 nsew power input
rlabel locali s 298660 252433 298799 252651 6 VPWR
port 613 nsew power input
rlabel locali s 298660 252651 298661 252759 6 VPWR
port 613 nsew power input
rlabel locali s 1259 252073 1340 252181 6 VPWR
port 613 nsew power input
rlabel locali s 1121 252181 1340 252399 6 VPWR
port 613 nsew power input
rlabel locali s 1104 252399 1340 252433 6 VPWR
port 613 nsew power input
rlabel locali s 1121 252433 1340 252651 6 VPWR
port 613 nsew power input
rlabel locali s 1259 252651 1340 252759 6 VPWR
port 613 nsew power input
rlabel locali s 298660 253161 298661 253269 6 VPWR
port 613 nsew power input
rlabel locali s 298660 253269 298799 253487 6 VPWR
port 613 nsew power input
rlabel locali s 298660 253487 298816 253521 6 VPWR
port 613 nsew power input
rlabel locali s 298660 253521 298799 253739 6 VPWR
port 613 nsew power input
rlabel locali s 298660 253739 298661 253847 6 VPWR
port 613 nsew power input
rlabel locali s 1259 253161 1340 253269 6 VPWR
port 613 nsew power input
rlabel locali s 1121 253269 1340 253487 6 VPWR
port 613 nsew power input
rlabel locali s 1104 253487 1340 253521 6 VPWR
port 613 nsew power input
rlabel locali s 1121 253521 1340 253739 6 VPWR
port 613 nsew power input
rlabel locali s 1259 253739 1340 253847 6 VPWR
port 613 nsew power input
rlabel locali s 298660 254249 298661 254357 6 VPWR
port 613 nsew power input
rlabel locali s 298660 254357 298799 254575 6 VPWR
port 613 nsew power input
rlabel locali s 298660 254575 298816 254609 6 VPWR
port 613 nsew power input
rlabel locali s 298660 254609 298799 254827 6 VPWR
port 613 nsew power input
rlabel locali s 298660 254827 298661 254935 6 VPWR
port 613 nsew power input
rlabel locali s 1259 254249 1340 254357 6 VPWR
port 613 nsew power input
rlabel locali s 1121 254357 1340 254575 6 VPWR
port 613 nsew power input
rlabel locali s 1104 254575 1340 254609 6 VPWR
port 613 nsew power input
rlabel locali s 1121 254609 1340 254827 6 VPWR
port 613 nsew power input
rlabel locali s 1259 254827 1340 254935 6 VPWR
port 613 nsew power input
rlabel locali s 298660 255337 298661 255445 6 VPWR
port 613 nsew power input
rlabel locali s 298660 255445 298799 255663 6 VPWR
port 613 nsew power input
rlabel locali s 298660 255663 298816 255697 6 VPWR
port 613 nsew power input
rlabel locali s 298660 255697 298799 255915 6 VPWR
port 613 nsew power input
rlabel locali s 298660 255915 298661 256023 6 VPWR
port 613 nsew power input
rlabel locali s 1259 255337 1340 255445 6 VPWR
port 613 nsew power input
rlabel locali s 1121 255445 1340 255663 6 VPWR
port 613 nsew power input
rlabel locali s 1104 255663 1340 255697 6 VPWR
port 613 nsew power input
rlabel locali s 1121 255697 1340 255915 6 VPWR
port 613 nsew power input
rlabel locali s 1259 255915 1340 256023 6 VPWR
port 613 nsew power input
rlabel locali s 298660 256425 298661 256533 6 VPWR
port 613 nsew power input
rlabel locali s 298660 256533 298799 256751 6 VPWR
port 613 nsew power input
rlabel locali s 298660 256751 298816 256785 6 VPWR
port 613 nsew power input
rlabel locali s 298660 256785 298799 257003 6 VPWR
port 613 nsew power input
rlabel locali s 298660 257003 298661 257111 6 VPWR
port 613 nsew power input
rlabel locali s 1259 256425 1340 256533 6 VPWR
port 613 nsew power input
rlabel locali s 1121 256533 1340 256751 6 VPWR
port 613 nsew power input
rlabel locali s 1104 256751 1340 256785 6 VPWR
port 613 nsew power input
rlabel locali s 1121 256785 1340 257003 6 VPWR
port 613 nsew power input
rlabel locali s 1259 257003 1340 257111 6 VPWR
port 613 nsew power input
rlabel locali s 298660 257513 298661 257621 6 VPWR
port 613 nsew power input
rlabel locali s 298660 257621 298799 257839 6 VPWR
port 613 nsew power input
rlabel locali s 298660 257839 298816 257873 6 VPWR
port 613 nsew power input
rlabel locali s 298660 257873 298799 258091 6 VPWR
port 613 nsew power input
rlabel locali s 298660 258091 298661 258199 6 VPWR
port 613 nsew power input
rlabel locali s 1259 257513 1340 257621 6 VPWR
port 613 nsew power input
rlabel locali s 1121 257621 1340 257839 6 VPWR
port 613 nsew power input
rlabel locali s 1104 257839 1340 257873 6 VPWR
port 613 nsew power input
rlabel locali s 1121 257873 1340 258091 6 VPWR
port 613 nsew power input
rlabel locali s 1259 258091 1340 258199 6 VPWR
port 613 nsew power input
rlabel locali s 298660 258601 298661 258709 6 VPWR
port 613 nsew power input
rlabel locali s 298660 258709 298799 258927 6 VPWR
port 613 nsew power input
rlabel locali s 298660 258927 298816 258961 6 VPWR
port 613 nsew power input
rlabel locali s 298660 258961 298799 259179 6 VPWR
port 613 nsew power input
rlabel locali s 298660 259179 298661 259287 6 VPWR
port 613 nsew power input
rlabel locali s 1259 258601 1340 258709 6 VPWR
port 613 nsew power input
rlabel locali s 1121 258709 1340 258927 6 VPWR
port 613 nsew power input
rlabel locali s 1104 258927 1340 258961 6 VPWR
port 613 nsew power input
rlabel locali s 1121 258961 1340 259179 6 VPWR
port 613 nsew power input
rlabel locali s 1259 259179 1340 259287 6 VPWR
port 613 nsew power input
rlabel locali s 298660 259689 298661 259797 6 VPWR
port 613 nsew power input
rlabel locali s 298660 259797 298799 260015 6 VPWR
port 613 nsew power input
rlabel locali s 298660 260015 298816 260049 6 VPWR
port 613 nsew power input
rlabel locali s 298660 260049 298799 260267 6 VPWR
port 613 nsew power input
rlabel locali s 298660 260267 298661 260375 6 VPWR
port 613 nsew power input
rlabel locali s 1259 259689 1340 259797 6 VPWR
port 613 nsew power input
rlabel locali s 1121 259797 1340 260015 6 VPWR
port 613 nsew power input
rlabel locali s 1104 260015 1340 260049 6 VPWR
port 613 nsew power input
rlabel locali s 1121 260049 1340 260267 6 VPWR
port 613 nsew power input
rlabel locali s 1259 260267 1340 260375 6 VPWR
port 613 nsew power input
rlabel locali s 298660 260777 298661 260885 6 VPWR
port 613 nsew power input
rlabel locali s 298660 260885 298799 261103 6 VPWR
port 613 nsew power input
rlabel locali s 298660 261103 298816 261137 6 VPWR
port 613 nsew power input
rlabel locali s 298660 261137 298799 261355 6 VPWR
port 613 nsew power input
rlabel locali s 298660 261355 298661 261463 6 VPWR
port 613 nsew power input
rlabel locali s 1259 260777 1340 260885 6 VPWR
port 613 nsew power input
rlabel locali s 1121 260885 1340 261103 6 VPWR
port 613 nsew power input
rlabel locali s 1104 261103 1340 261137 6 VPWR
port 613 nsew power input
rlabel locali s 1121 261137 1340 261355 6 VPWR
port 613 nsew power input
rlabel locali s 1259 261355 1340 261463 6 VPWR
port 613 nsew power input
rlabel locali s 298660 261865 298661 261973 6 VPWR
port 613 nsew power input
rlabel locali s 298660 261973 298799 262191 6 VPWR
port 613 nsew power input
rlabel locali s 298660 262191 298816 262225 6 VPWR
port 613 nsew power input
rlabel locali s 298660 262225 298799 262443 6 VPWR
port 613 nsew power input
rlabel locali s 298660 262443 298661 262551 6 VPWR
port 613 nsew power input
rlabel locali s 1259 261865 1340 261973 6 VPWR
port 613 nsew power input
rlabel locali s 1121 261973 1340 262191 6 VPWR
port 613 nsew power input
rlabel locali s 1104 262191 1340 262225 6 VPWR
port 613 nsew power input
rlabel locali s 1121 262225 1340 262443 6 VPWR
port 613 nsew power input
rlabel locali s 1259 262443 1340 262551 6 VPWR
port 613 nsew power input
rlabel locali s 298660 262953 298661 263061 6 VPWR
port 613 nsew power input
rlabel locali s 298660 263061 298799 263279 6 VPWR
port 613 nsew power input
rlabel locali s 298660 263279 298816 263313 6 VPWR
port 613 nsew power input
rlabel locali s 298660 263313 298799 263531 6 VPWR
port 613 nsew power input
rlabel locali s 298660 263531 298661 263639 6 VPWR
port 613 nsew power input
rlabel locali s 1259 262953 1340 263061 6 VPWR
port 613 nsew power input
rlabel locali s 1121 263061 1340 263279 6 VPWR
port 613 nsew power input
rlabel locali s 1104 263279 1340 263313 6 VPWR
port 613 nsew power input
rlabel locali s 1121 263313 1340 263531 6 VPWR
port 613 nsew power input
rlabel locali s 1259 263531 1340 263639 6 VPWR
port 613 nsew power input
rlabel locali s 298660 264041 298661 264149 6 VPWR
port 613 nsew power input
rlabel locali s 298660 264149 298799 264367 6 VPWR
port 613 nsew power input
rlabel locali s 298660 264367 298816 264401 6 VPWR
port 613 nsew power input
rlabel locali s 298660 264401 298799 264619 6 VPWR
port 613 nsew power input
rlabel locali s 298660 264619 298661 264727 6 VPWR
port 613 nsew power input
rlabel locali s 1259 264041 1340 264149 6 VPWR
port 613 nsew power input
rlabel locali s 1121 264149 1340 264367 6 VPWR
port 613 nsew power input
rlabel locali s 1104 264367 1340 264401 6 VPWR
port 613 nsew power input
rlabel locali s 1121 264401 1340 264619 6 VPWR
port 613 nsew power input
rlabel locali s 1259 264619 1340 264727 6 VPWR
port 613 nsew power input
rlabel locali s 298660 265129 298661 265237 6 VPWR
port 613 nsew power input
rlabel locali s 298660 265237 298799 265455 6 VPWR
port 613 nsew power input
rlabel locali s 298660 265455 298816 265489 6 VPWR
port 613 nsew power input
rlabel locali s 298660 265489 298799 265707 6 VPWR
port 613 nsew power input
rlabel locali s 298660 265707 298661 265815 6 VPWR
port 613 nsew power input
rlabel locali s 1259 265129 1340 265237 6 VPWR
port 613 nsew power input
rlabel locali s 1121 265237 1340 265455 6 VPWR
port 613 nsew power input
rlabel locali s 1104 265455 1340 265489 6 VPWR
port 613 nsew power input
rlabel locali s 1121 265489 1340 265707 6 VPWR
port 613 nsew power input
rlabel locali s 1259 265707 1340 265815 6 VPWR
port 613 nsew power input
rlabel locali s 298660 266217 298661 266325 6 VPWR
port 613 nsew power input
rlabel locali s 298660 266325 298799 266543 6 VPWR
port 613 nsew power input
rlabel locali s 298660 266543 298816 266577 6 VPWR
port 613 nsew power input
rlabel locali s 298660 266577 298799 266795 6 VPWR
port 613 nsew power input
rlabel locali s 298660 266795 298661 266903 6 VPWR
port 613 nsew power input
rlabel locali s 1259 266217 1340 266325 6 VPWR
port 613 nsew power input
rlabel locali s 1121 266325 1340 266543 6 VPWR
port 613 nsew power input
rlabel locali s 1104 266543 1340 266577 6 VPWR
port 613 nsew power input
rlabel locali s 1121 266577 1340 266795 6 VPWR
port 613 nsew power input
rlabel locali s 1259 266795 1340 266903 6 VPWR
port 613 nsew power input
rlabel locali s 298660 267305 298661 267413 6 VPWR
port 613 nsew power input
rlabel locali s 298660 267413 298799 267631 6 VPWR
port 613 nsew power input
rlabel locali s 298660 267631 298816 267665 6 VPWR
port 613 nsew power input
rlabel locali s 298660 267665 298799 267883 6 VPWR
port 613 nsew power input
rlabel locali s 298660 267883 298661 267991 6 VPWR
port 613 nsew power input
rlabel locali s 1259 267305 1340 267413 6 VPWR
port 613 nsew power input
rlabel locali s 1121 267413 1340 267631 6 VPWR
port 613 nsew power input
rlabel locali s 1104 267631 1340 267665 6 VPWR
port 613 nsew power input
rlabel locali s 1121 267665 1340 267883 6 VPWR
port 613 nsew power input
rlabel locali s 1259 267883 1340 267991 6 VPWR
port 613 nsew power input
rlabel locali s 298660 268393 298661 268501 6 VPWR
port 613 nsew power input
rlabel locali s 298660 268501 298799 268719 6 VPWR
port 613 nsew power input
rlabel locali s 298660 268719 298816 268753 6 VPWR
port 613 nsew power input
rlabel locali s 298660 268753 298799 268971 6 VPWR
port 613 nsew power input
rlabel locali s 298660 268971 298661 269079 6 VPWR
port 613 nsew power input
rlabel locali s 1259 268393 1340 268501 6 VPWR
port 613 nsew power input
rlabel locali s 1121 268501 1340 268719 6 VPWR
port 613 nsew power input
rlabel locali s 1104 268719 1340 268753 6 VPWR
port 613 nsew power input
rlabel locali s 1121 268753 1340 268971 6 VPWR
port 613 nsew power input
rlabel locali s 1259 268971 1340 269079 6 VPWR
port 613 nsew power input
rlabel locali s 298660 269481 298661 269589 6 VPWR
port 613 nsew power input
rlabel locali s 298660 269589 298799 269807 6 VPWR
port 613 nsew power input
rlabel locali s 298660 269807 298816 269841 6 VPWR
port 613 nsew power input
rlabel locali s 298660 269841 298799 270059 6 VPWR
port 613 nsew power input
rlabel locali s 298660 270059 298661 270167 6 VPWR
port 613 nsew power input
rlabel locali s 1259 269481 1340 269589 6 VPWR
port 613 nsew power input
rlabel locali s 1121 269589 1340 269807 6 VPWR
port 613 nsew power input
rlabel locali s 1104 269807 1340 269841 6 VPWR
port 613 nsew power input
rlabel locali s 1121 269841 1340 270059 6 VPWR
port 613 nsew power input
rlabel locali s 1259 270059 1340 270167 6 VPWR
port 613 nsew power input
rlabel locali s 298660 270569 298661 270677 6 VPWR
port 613 nsew power input
rlabel locali s 298660 270677 298799 270895 6 VPWR
port 613 nsew power input
rlabel locali s 298660 270895 298816 270929 6 VPWR
port 613 nsew power input
rlabel locali s 298660 270929 298799 271147 6 VPWR
port 613 nsew power input
rlabel locali s 298660 271147 298661 271255 6 VPWR
port 613 nsew power input
rlabel locali s 1259 270569 1340 270677 6 VPWR
port 613 nsew power input
rlabel locali s 1121 270677 1340 270895 6 VPWR
port 613 nsew power input
rlabel locali s 1104 270895 1340 270929 6 VPWR
port 613 nsew power input
rlabel locali s 1121 270929 1340 271147 6 VPWR
port 613 nsew power input
rlabel locali s 1259 271147 1340 271255 6 VPWR
port 613 nsew power input
rlabel locali s 298660 271657 298661 271765 6 VPWR
port 613 nsew power input
rlabel locali s 298660 271765 298799 271983 6 VPWR
port 613 nsew power input
rlabel locali s 298660 271983 298816 272017 6 VPWR
port 613 nsew power input
rlabel locali s 298660 272017 298799 272235 6 VPWR
port 613 nsew power input
rlabel locali s 298660 272235 298661 272343 6 VPWR
port 613 nsew power input
rlabel locali s 1259 271657 1340 271765 6 VPWR
port 613 nsew power input
rlabel locali s 1121 271765 1340 271983 6 VPWR
port 613 nsew power input
rlabel locali s 1104 271983 1340 272017 6 VPWR
port 613 nsew power input
rlabel locali s 1121 272017 1340 272235 6 VPWR
port 613 nsew power input
rlabel locali s 1259 272235 1340 272343 6 VPWR
port 613 nsew power input
rlabel locali s 298660 272745 298661 272853 6 VPWR
port 613 nsew power input
rlabel locali s 298660 272853 298799 273071 6 VPWR
port 613 nsew power input
rlabel locali s 298660 273071 298816 273105 6 VPWR
port 613 nsew power input
rlabel locali s 298660 273105 298799 273323 6 VPWR
port 613 nsew power input
rlabel locali s 298660 273323 298661 273431 6 VPWR
port 613 nsew power input
rlabel locali s 1259 272745 1340 272853 6 VPWR
port 613 nsew power input
rlabel locali s 1121 272853 1340 273071 6 VPWR
port 613 nsew power input
rlabel locali s 1104 273071 1340 273105 6 VPWR
port 613 nsew power input
rlabel locali s 1121 273105 1340 273323 6 VPWR
port 613 nsew power input
rlabel locali s 1259 273323 1340 273431 6 VPWR
port 613 nsew power input
rlabel locali s 298660 273833 298661 273941 6 VPWR
port 613 nsew power input
rlabel locali s 298660 273941 298799 274159 6 VPWR
port 613 nsew power input
rlabel locali s 298660 274159 298816 274193 6 VPWR
port 613 nsew power input
rlabel locali s 298660 274193 298799 274411 6 VPWR
port 613 nsew power input
rlabel locali s 298660 274411 298661 274519 6 VPWR
port 613 nsew power input
rlabel locali s 1259 273833 1340 273941 6 VPWR
port 613 nsew power input
rlabel locali s 1121 273941 1340 274159 6 VPWR
port 613 nsew power input
rlabel locali s 1104 274159 1340 274193 6 VPWR
port 613 nsew power input
rlabel locali s 1121 274193 1340 274411 6 VPWR
port 613 nsew power input
rlabel locali s 1259 274411 1340 274519 6 VPWR
port 613 nsew power input
rlabel locali s 298660 274921 298661 275029 6 VPWR
port 613 nsew power input
rlabel locali s 298660 275029 298799 275247 6 VPWR
port 613 nsew power input
rlabel locali s 298660 275247 298816 275281 6 VPWR
port 613 nsew power input
rlabel locali s 298660 275281 298799 275499 6 VPWR
port 613 nsew power input
rlabel locali s 298660 275499 298661 275607 6 VPWR
port 613 nsew power input
rlabel locali s 1259 274921 1340 275029 6 VPWR
port 613 nsew power input
rlabel locali s 1121 275029 1340 275247 6 VPWR
port 613 nsew power input
rlabel locali s 1104 275247 1340 275281 6 VPWR
port 613 nsew power input
rlabel locali s 1121 275281 1340 275499 6 VPWR
port 613 nsew power input
rlabel locali s 1259 275499 1340 275607 6 VPWR
port 613 nsew power input
rlabel locali s 298660 276009 298661 276117 6 VPWR
port 613 nsew power input
rlabel locali s 298660 276117 298799 276335 6 VPWR
port 613 nsew power input
rlabel locali s 298660 276335 298816 276369 6 VPWR
port 613 nsew power input
rlabel locali s 298660 276369 298799 276587 6 VPWR
port 613 nsew power input
rlabel locali s 298660 276587 298661 276695 6 VPWR
port 613 nsew power input
rlabel locali s 1259 276009 1340 276117 6 VPWR
port 613 nsew power input
rlabel locali s 1121 276117 1340 276335 6 VPWR
port 613 nsew power input
rlabel locali s 1104 276335 1340 276369 6 VPWR
port 613 nsew power input
rlabel locali s 1121 276369 1340 276587 6 VPWR
port 613 nsew power input
rlabel locali s 1259 276587 1340 276695 6 VPWR
port 613 nsew power input
rlabel locali s 298660 277097 298661 277205 6 VPWR
port 613 nsew power input
rlabel locali s 298660 277205 298799 277423 6 VPWR
port 613 nsew power input
rlabel locali s 298660 277423 298816 277457 6 VPWR
port 613 nsew power input
rlabel locali s 298660 277457 298799 277675 6 VPWR
port 613 nsew power input
rlabel locali s 298660 277675 298661 277783 6 VPWR
port 613 nsew power input
rlabel locali s 1259 277097 1340 277205 6 VPWR
port 613 nsew power input
rlabel locali s 1121 277205 1340 277423 6 VPWR
port 613 nsew power input
rlabel locali s 1104 277423 1340 277457 6 VPWR
port 613 nsew power input
rlabel locali s 1121 277457 1340 277675 6 VPWR
port 613 nsew power input
rlabel locali s 1259 277675 1340 277783 6 VPWR
port 613 nsew power input
rlabel locali s 298660 278185 298661 278293 6 VPWR
port 613 nsew power input
rlabel locali s 298660 278293 298799 278511 6 VPWR
port 613 nsew power input
rlabel locali s 298660 278511 298816 278545 6 VPWR
port 613 nsew power input
rlabel locali s 298660 278545 298799 278763 6 VPWR
port 613 nsew power input
rlabel locali s 298660 278763 298661 278871 6 VPWR
port 613 nsew power input
rlabel locali s 1259 278185 1340 278293 6 VPWR
port 613 nsew power input
rlabel locali s 1121 278293 1340 278511 6 VPWR
port 613 nsew power input
rlabel locali s 1104 278511 1340 278545 6 VPWR
port 613 nsew power input
rlabel locali s 1121 278545 1340 278763 6 VPWR
port 613 nsew power input
rlabel locali s 1259 278763 1340 278871 6 VPWR
port 613 nsew power input
rlabel locali s 298660 279273 298661 279381 6 VPWR
port 613 nsew power input
rlabel locali s 298660 279381 298799 279599 6 VPWR
port 613 nsew power input
rlabel locali s 298660 279599 298816 279633 6 VPWR
port 613 nsew power input
rlabel locali s 298660 279633 298799 279851 6 VPWR
port 613 nsew power input
rlabel locali s 298660 279851 298661 279959 6 VPWR
port 613 nsew power input
rlabel locali s 1259 279273 1340 279381 6 VPWR
port 613 nsew power input
rlabel locali s 1121 279381 1340 279599 6 VPWR
port 613 nsew power input
rlabel locali s 1104 279599 1340 279633 6 VPWR
port 613 nsew power input
rlabel locali s 1121 279633 1340 279851 6 VPWR
port 613 nsew power input
rlabel locali s 1259 279851 1340 279959 6 VPWR
port 613 nsew power input
rlabel locali s 298660 280361 298661 280469 6 VPWR
port 613 nsew power input
rlabel locali s 298660 280469 298799 280687 6 VPWR
port 613 nsew power input
rlabel locali s 298660 280687 298816 280721 6 VPWR
port 613 nsew power input
rlabel locali s 298660 280721 298799 280939 6 VPWR
port 613 nsew power input
rlabel locali s 298660 280939 298661 281047 6 VPWR
port 613 nsew power input
rlabel locali s 1259 280361 1340 280469 6 VPWR
port 613 nsew power input
rlabel locali s 1121 280469 1340 280687 6 VPWR
port 613 nsew power input
rlabel locali s 1104 280687 1340 280721 6 VPWR
port 613 nsew power input
rlabel locali s 1121 280721 1340 280939 6 VPWR
port 613 nsew power input
rlabel locali s 1259 280939 1340 281047 6 VPWR
port 613 nsew power input
rlabel locali s 298660 281449 298661 281557 6 VPWR
port 613 nsew power input
rlabel locali s 298660 281557 298799 281775 6 VPWR
port 613 nsew power input
rlabel locali s 298660 281775 298816 281809 6 VPWR
port 613 nsew power input
rlabel locali s 298660 281809 298799 282027 6 VPWR
port 613 nsew power input
rlabel locali s 298660 282027 298661 282135 6 VPWR
port 613 nsew power input
rlabel locali s 1259 281449 1340 281557 6 VPWR
port 613 nsew power input
rlabel locali s 1121 281557 1340 281775 6 VPWR
port 613 nsew power input
rlabel locali s 1104 281775 1340 281809 6 VPWR
port 613 nsew power input
rlabel locali s 1121 281809 1340 282027 6 VPWR
port 613 nsew power input
rlabel locali s 1259 282027 1340 282135 6 VPWR
port 613 nsew power input
rlabel locali s 298660 282537 298661 282645 6 VPWR
port 613 nsew power input
rlabel locali s 298660 282645 298799 282863 6 VPWR
port 613 nsew power input
rlabel locali s 298660 282863 298816 282897 6 VPWR
port 613 nsew power input
rlabel locali s 298660 282897 298799 283115 6 VPWR
port 613 nsew power input
rlabel locali s 298660 283115 298661 283223 6 VPWR
port 613 nsew power input
rlabel locali s 1259 282537 1340 282645 6 VPWR
port 613 nsew power input
rlabel locali s 1121 282645 1340 282863 6 VPWR
port 613 nsew power input
rlabel locali s 1104 282863 1340 282897 6 VPWR
port 613 nsew power input
rlabel locali s 1121 282897 1340 283115 6 VPWR
port 613 nsew power input
rlabel locali s 1259 283115 1340 283223 6 VPWR
port 613 nsew power input
rlabel locali s 298660 283625 298661 283733 6 VPWR
port 613 nsew power input
rlabel locali s 298660 283733 298799 283951 6 VPWR
port 613 nsew power input
rlabel locali s 298660 283951 298816 283985 6 VPWR
port 613 nsew power input
rlabel locali s 298660 283985 298799 284203 6 VPWR
port 613 nsew power input
rlabel locali s 298660 284203 298661 284311 6 VPWR
port 613 nsew power input
rlabel locali s 1259 283625 1340 283733 6 VPWR
port 613 nsew power input
rlabel locali s 1121 283733 1340 283951 6 VPWR
port 613 nsew power input
rlabel locali s 1104 283951 1340 283985 6 VPWR
port 613 nsew power input
rlabel locali s 1121 283985 1340 284203 6 VPWR
port 613 nsew power input
rlabel locali s 1259 284203 1340 284311 6 VPWR
port 613 nsew power input
rlabel locali s 298660 284713 298661 284821 6 VPWR
port 613 nsew power input
rlabel locali s 298660 284821 298799 285039 6 VPWR
port 613 nsew power input
rlabel locali s 298660 285039 298816 285073 6 VPWR
port 613 nsew power input
rlabel locali s 298660 285073 298799 285291 6 VPWR
port 613 nsew power input
rlabel locali s 298660 285291 298661 285399 6 VPWR
port 613 nsew power input
rlabel locali s 1259 284713 1340 284821 6 VPWR
port 613 nsew power input
rlabel locali s 1121 284821 1340 285039 6 VPWR
port 613 nsew power input
rlabel locali s 1104 285039 1340 285073 6 VPWR
port 613 nsew power input
rlabel locali s 1121 285073 1340 285291 6 VPWR
port 613 nsew power input
rlabel locali s 1259 285291 1340 285399 6 VPWR
port 613 nsew power input
rlabel locali s 298660 285801 298661 285909 6 VPWR
port 613 nsew power input
rlabel locali s 298660 285909 298799 286127 6 VPWR
port 613 nsew power input
rlabel locali s 298660 286127 298816 286161 6 VPWR
port 613 nsew power input
rlabel locali s 298660 286161 298799 286379 6 VPWR
port 613 nsew power input
rlabel locali s 298660 286379 298661 286487 6 VPWR
port 613 nsew power input
rlabel locali s 1259 285801 1340 285909 6 VPWR
port 613 nsew power input
rlabel locali s 1121 285909 1340 286127 6 VPWR
port 613 nsew power input
rlabel locali s 1104 286127 1340 286161 6 VPWR
port 613 nsew power input
rlabel locali s 1121 286161 1340 286379 6 VPWR
port 613 nsew power input
rlabel locali s 1259 286379 1340 286487 6 VPWR
port 613 nsew power input
rlabel locali s 298660 286889 298661 286997 6 VPWR
port 613 nsew power input
rlabel locali s 298660 286997 298799 287215 6 VPWR
port 613 nsew power input
rlabel locali s 298660 287215 298816 287249 6 VPWR
port 613 nsew power input
rlabel locali s 298660 287249 298799 287467 6 VPWR
port 613 nsew power input
rlabel locali s 298660 287467 298661 287575 6 VPWR
port 613 nsew power input
rlabel locali s 1259 286889 1340 286997 6 VPWR
port 613 nsew power input
rlabel locali s 1121 286997 1340 287215 6 VPWR
port 613 nsew power input
rlabel locali s 1104 287215 1340 287249 6 VPWR
port 613 nsew power input
rlabel locali s 1121 287249 1340 287467 6 VPWR
port 613 nsew power input
rlabel locali s 1259 287467 1340 287575 6 VPWR
port 613 nsew power input
rlabel locali s 298660 287977 298661 288085 6 VPWR
port 613 nsew power input
rlabel locali s 298660 288085 298799 288303 6 VPWR
port 613 nsew power input
rlabel locali s 298660 288303 298816 288337 6 VPWR
port 613 nsew power input
rlabel locali s 298660 288337 298799 288555 6 VPWR
port 613 nsew power input
rlabel locali s 298660 288555 298661 288663 6 VPWR
port 613 nsew power input
rlabel locali s 1259 287977 1340 288085 6 VPWR
port 613 nsew power input
rlabel locali s 1121 288085 1340 288303 6 VPWR
port 613 nsew power input
rlabel locali s 1104 288303 1340 288337 6 VPWR
port 613 nsew power input
rlabel locali s 1121 288337 1340 288555 6 VPWR
port 613 nsew power input
rlabel locali s 1259 288555 1340 288663 6 VPWR
port 613 nsew power input
rlabel locali s 298660 289065 298661 289173 6 VPWR
port 613 nsew power input
rlabel locali s 298660 289173 298799 289391 6 VPWR
port 613 nsew power input
rlabel locali s 298660 289391 298816 289425 6 VPWR
port 613 nsew power input
rlabel locali s 298660 289425 298799 289643 6 VPWR
port 613 nsew power input
rlabel locali s 298660 289643 298661 289751 6 VPWR
port 613 nsew power input
rlabel locali s 1259 289065 1340 289173 6 VPWR
port 613 nsew power input
rlabel locali s 1121 289173 1340 289391 6 VPWR
port 613 nsew power input
rlabel locali s 1104 289391 1340 289425 6 VPWR
port 613 nsew power input
rlabel locali s 1121 289425 1340 289643 6 VPWR
port 613 nsew power input
rlabel locali s 1259 289643 1340 289751 6 VPWR
port 613 nsew power input
rlabel locali s 298660 290153 298661 290261 6 VPWR
port 613 nsew power input
rlabel locali s 298660 290261 298799 290479 6 VPWR
port 613 nsew power input
rlabel locali s 298660 290479 298816 290513 6 VPWR
port 613 nsew power input
rlabel locali s 298660 290513 298799 290731 6 VPWR
port 613 nsew power input
rlabel locali s 298660 290731 298661 290839 6 VPWR
port 613 nsew power input
rlabel locali s 1259 290153 1340 290261 6 VPWR
port 613 nsew power input
rlabel locali s 1121 290261 1340 290479 6 VPWR
port 613 nsew power input
rlabel locali s 1104 290479 1340 290513 6 VPWR
port 613 nsew power input
rlabel locali s 1121 290513 1340 290731 6 VPWR
port 613 nsew power input
rlabel locali s 1259 290731 1340 290839 6 VPWR
port 613 nsew power input
rlabel locali s 298660 291241 298661 291349 6 VPWR
port 613 nsew power input
rlabel locali s 298660 291349 298799 291567 6 VPWR
port 613 nsew power input
rlabel locali s 298660 291567 298816 291601 6 VPWR
port 613 nsew power input
rlabel locali s 298660 291601 298799 291819 6 VPWR
port 613 nsew power input
rlabel locali s 298660 291819 298661 291927 6 VPWR
port 613 nsew power input
rlabel locali s 1259 291241 1340 291349 6 VPWR
port 613 nsew power input
rlabel locali s 1121 291349 1340 291567 6 VPWR
port 613 nsew power input
rlabel locali s 1104 291567 1340 291601 6 VPWR
port 613 nsew power input
rlabel locali s 1121 291601 1340 291819 6 VPWR
port 613 nsew power input
rlabel locali s 1259 291819 1340 291927 6 VPWR
port 613 nsew power input
rlabel locali s 298660 292329 298661 292437 6 VPWR
port 613 nsew power input
rlabel locali s 298660 292437 298799 292655 6 VPWR
port 613 nsew power input
rlabel locali s 298660 292655 298816 292689 6 VPWR
port 613 nsew power input
rlabel locali s 298660 292689 298799 292907 6 VPWR
port 613 nsew power input
rlabel locali s 298660 292907 298661 293015 6 VPWR
port 613 nsew power input
rlabel locali s 1259 292329 1340 292437 6 VPWR
port 613 nsew power input
rlabel locali s 1121 292437 1340 292655 6 VPWR
port 613 nsew power input
rlabel locali s 1104 292655 1340 292689 6 VPWR
port 613 nsew power input
rlabel locali s 1121 292689 1340 292907 6 VPWR
port 613 nsew power input
rlabel locali s 1259 292907 1340 293015 6 VPWR
port 613 nsew power input
rlabel locali s 298660 293417 298661 293525 6 VPWR
port 613 nsew power input
rlabel locali s 298660 293525 298799 293743 6 VPWR
port 613 nsew power input
rlabel locali s 298660 293743 298816 293777 6 VPWR
port 613 nsew power input
rlabel locali s 298660 293777 298799 293995 6 VPWR
port 613 nsew power input
rlabel locali s 298660 293995 298661 294103 6 VPWR
port 613 nsew power input
rlabel locali s 1259 293417 1340 293525 6 VPWR
port 613 nsew power input
rlabel locali s 1121 293525 1340 293743 6 VPWR
port 613 nsew power input
rlabel locali s 1104 293743 1340 293777 6 VPWR
port 613 nsew power input
rlabel locali s 1121 293777 1340 293995 6 VPWR
port 613 nsew power input
rlabel locali s 1259 293995 1340 294103 6 VPWR
port 613 nsew power input
rlabel locali s 298660 294505 298661 294613 6 VPWR
port 613 nsew power input
rlabel locali s 298660 294613 298799 294831 6 VPWR
port 613 nsew power input
rlabel locali s 298660 294831 298816 294865 6 VPWR
port 613 nsew power input
rlabel locali s 298660 294865 298799 295083 6 VPWR
port 613 nsew power input
rlabel locali s 298660 295083 298661 295191 6 VPWR
port 613 nsew power input
rlabel locali s 1259 294505 1340 294613 6 VPWR
port 613 nsew power input
rlabel locali s 1121 294613 1340 294831 6 VPWR
port 613 nsew power input
rlabel locali s 1104 294831 1340 294865 6 VPWR
port 613 nsew power input
rlabel locali s 1121 294865 1340 295083 6 VPWR
port 613 nsew power input
rlabel locali s 1259 295083 1340 295191 6 VPWR
port 613 nsew power input
rlabel locali s 298660 295593 298661 295701 6 VPWR
port 613 nsew power input
rlabel locali s 298660 295701 298799 295919 6 VPWR
port 613 nsew power input
rlabel locali s 298660 295919 298816 295953 6 VPWR
port 613 nsew power input
rlabel locali s 298660 295953 298799 296171 6 VPWR
port 613 nsew power input
rlabel locali s 298660 296171 298661 296279 6 VPWR
port 613 nsew power input
rlabel locali s 1259 295593 1340 295701 6 VPWR
port 613 nsew power input
rlabel locali s 1121 295701 1340 295919 6 VPWR
port 613 nsew power input
rlabel locali s 1104 295919 1340 295953 6 VPWR
port 613 nsew power input
rlabel locali s 1121 295953 1340 296171 6 VPWR
port 613 nsew power input
rlabel locali s 1259 296171 1340 296279 6 VPWR
port 613 nsew power input
rlabel locali s 298660 296681 298661 296789 6 VPWR
port 613 nsew power input
rlabel locali s 298660 296789 298799 297007 6 VPWR
port 613 nsew power input
rlabel locali s 298660 297007 298816 297041 6 VPWR
port 613 nsew power input
rlabel locali s 298660 297041 298799 297259 6 VPWR
port 613 nsew power input
rlabel locali s 298660 297259 298661 297367 6 VPWR
port 613 nsew power input
rlabel locali s 1259 296681 1340 296789 6 VPWR
port 613 nsew power input
rlabel locali s 1121 296789 1340 297007 6 VPWR
port 613 nsew power input
rlabel locali s 1104 297007 1340 297041 6 VPWR
port 613 nsew power input
rlabel locali s 1121 297041 1340 297259 6 VPWR
port 613 nsew power input
rlabel locali s 1259 297259 1340 297367 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 2138 298854 2459 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 2138 1340 2459 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 2981 298854 3547 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 2981 1340 3547 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 4069 298854 4635 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 4069 1340 4635 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 5157 298854 5723 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 5157 1340 5723 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 6245 298854 6811 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 6245 1340 6811 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 7333 298854 7899 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 7333 1340 7899 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 8421 298854 8987 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 8421 1340 8987 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 9509 298854 10075 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 9509 1340 10075 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 10597 298854 11163 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 10597 1340 11163 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 11685 298854 12251 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 11685 1340 12251 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 12773 298854 13339 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 12773 1340 13339 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 13861 298854 14427 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 13861 1340 14427 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 14949 298854 15515 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 14949 1340 15515 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 16037 298854 16603 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 16037 1340 16603 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 17125 298854 17691 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 17125 1340 17691 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 18213 298854 18779 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 18213 1340 18779 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 19301 298854 19867 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 19301 1340 19867 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 20389 298854 20955 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 20389 1340 20955 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 21477 298854 22043 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 21477 1340 22043 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 22565 298854 23131 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 22565 1340 23131 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 23653 298854 24219 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 23653 1340 24219 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 24741 298854 25307 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 24741 1340 25307 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 25829 298854 26395 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 25829 1340 26395 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 26917 298854 27483 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 26917 1340 27483 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 28005 298854 28571 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 28005 1340 28571 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 29093 298854 29659 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 29093 1340 29659 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 30181 298854 30747 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 30181 1340 30747 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 31269 298854 31835 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 31269 1340 31835 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 32357 298854 32923 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 32357 1340 32923 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 33445 298854 34011 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 33445 1340 34011 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 34533 298854 35099 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 34533 1340 35099 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 35621 298854 36187 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 35621 1340 36187 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 36709 298854 37275 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 36709 1340 37275 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 37797 298854 38363 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 37797 1340 38363 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 38885 298854 39451 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 38885 1340 39451 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 39973 298854 40539 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 39973 1340 40539 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 41061 298854 41627 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 41061 1340 41627 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 42149 298854 42715 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 42149 1340 42715 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 43237 298854 43803 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 43237 1340 43803 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 44325 298854 44891 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 44325 1340 44891 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 45413 298854 45979 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 45413 1340 45979 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 46501 298854 47067 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 46501 1340 47067 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 47589 298854 48155 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 47589 1340 48155 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 48677 298854 49243 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 48677 1340 49243 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 49765 298854 50331 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 49765 1340 50331 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 50853 298854 51419 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 50853 1340 51419 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 51941 298854 52507 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 51941 1340 52507 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 53029 298854 53595 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 53029 1340 53595 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 54117 298854 54683 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 54117 1340 54683 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 55205 298854 55771 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 55205 1340 55771 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 56293 298854 56859 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 56293 1340 56859 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 57381 298854 57947 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 57381 1340 57947 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 58469 298854 59035 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 58469 1340 59035 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 59557 298854 60123 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 59557 1340 60123 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 60645 298854 61211 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 60645 1340 61211 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 61733 298854 62299 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 61733 1340 62299 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 62821 298854 63387 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 62821 1340 63387 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 63909 298854 64475 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 63909 1340 64475 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 64997 298854 65563 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 64997 1340 65563 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 66085 298854 66651 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 66085 1340 66651 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 67173 298854 67739 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 67173 1340 67739 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 68261 298854 68827 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 68261 1340 68827 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 69349 298854 69915 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 69349 1340 69915 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 70437 298854 71003 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 70437 1340 71003 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 71525 298854 72091 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 71525 1340 72091 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 72613 298854 73179 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 72613 1340 73179 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 73701 298854 74267 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 73701 1340 74267 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 74789 298854 75355 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 74789 1340 75355 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 75877 298854 76443 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 75877 1340 76443 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 76965 298854 77531 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 76965 1340 77531 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 78053 298854 78619 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 78053 1340 78619 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 79141 298854 79707 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 79141 1340 79707 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 80229 298854 80795 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 80229 1340 80795 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 81317 298854 81883 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 81317 1340 81883 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 82405 298854 82971 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 82405 1340 82971 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 83493 298854 84059 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 83493 1340 84059 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 84581 298854 85147 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 84581 1340 85147 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 85669 298854 86235 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 85669 1340 86235 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 86757 298854 87323 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 86757 1340 87323 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 87845 298854 88411 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 87845 1340 88411 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 88933 298854 89499 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 88933 1340 89499 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 90021 298854 90587 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 90021 1340 90587 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 91109 298854 91675 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 91109 1340 91675 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 92197 298854 92763 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 92197 1340 92763 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 93285 298854 93851 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 93285 1340 93851 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 94373 298854 94939 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 94373 1340 94939 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 95461 298854 96027 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 95461 1340 96027 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 96549 298854 97115 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 96549 1340 97115 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 97637 298854 98203 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 97637 1340 98203 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 98725 298854 99291 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 98725 1340 99291 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 99813 298854 100379 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 99813 1340 100379 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 100901 298854 101467 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 100901 1340 101467 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 101989 298854 102555 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 101989 1340 102555 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 103077 298854 103643 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 103077 1340 103643 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 104165 298854 104731 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 104165 1340 104731 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 105253 298854 105819 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 105253 1340 105819 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 106341 298854 106907 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 106341 1340 106907 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 107429 298854 107995 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 107429 1340 107995 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 108517 298854 109083 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 108517 1340 109083 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 109605 298854 110171 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 109605 1340 110171 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 110693 298854 111259 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 110693 1340 111259 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 111781 298854 112347 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 111781 1340 112347 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 112869 298854 113435 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 112869 1340 113435 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 113957 298854 114523 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 113957 1340 114523 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 115045 298854 115611 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 115045 1340 115611 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 116133 298854 116699 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 116133 1340 116699 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 117221 298854 117787 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 117221 1340 117787 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 118309 298854 118875 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 118309 1340 118875 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 119397 298854 119963 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 119397 1340 119963 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 120485 298854 121051 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 120485 1340 121051 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 121573 298854 122139 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 121573 1340 122139 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 122661 298854 123227 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 122661 1340 123227 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 123749 298854 124315 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 123749 1340 124315 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 124837 298854 125403 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 124837 1340 125403 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 125925 298854 126491 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 125925 1340 126491 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 127013 298854 127579 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 127013 1340 127579 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 128101 298854 128667 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 128101 1340 128667 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 129189 298854 129755 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 129189 1340 129755 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 130277 298854 130843 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 130277 1340 130843 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 131365 298854 131931 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 131365 1340 131931 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 132453 298854 133019 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 132453 1340 133019 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 133541 298854 134107 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 133541 1340 134107 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 134629 298854 135195 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 134629 1340 135195 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 135717 298854 136283 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 135717 1340 136283 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 136805 298854 137371 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 136805 1340 137371 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 137893 298854 138459 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 137893 1340 138459 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 138981 298854 139547 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 138981 1340 139547 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 140069 298854 140635 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 140069 1340 140635 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 141157 298854 141723 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 141157 1340 141723 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 142245 298854 142811 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 142245 1340 142811 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 143333 298854 143899 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 143333 1340 143899 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 144421 298854 144987 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 144421 1340 144987 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 145509 298854 146075 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 145509 1340 146075 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 146597 298854 147163 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 146597 1340 147163 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 147685 298854 148251 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 147685 1340 148251 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 148773 298854 149339 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 148773 1340 149339 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 149861 298854 150427 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 149861 1340 150427 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 150949 298854 151515 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 150949 1340 151515 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 152037 298854 152603 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 152037 1340 152603 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 153125 298854 153691 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 153125 1340 153691 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 154213 298854 154779 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 154213 1340 154779 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 155301 298854 155867 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 155301 1340 155867 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 156389 298854 156955 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 156389 1340 156955 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 157477 298854 158043 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 157477 1340 158043 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 158565 298854 159131 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 158565 1340 159131 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 159653 298854 160219 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 159653 1340 160219 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 160741 298854 161307 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 160741 1340 161307 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 161829 298854 162395 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 161829 1340 162395 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 162917 298854 163483 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 162917 1340 163483 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 164005 298854 164571 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 164005 1340 164571 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 165093 298854 165659 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 165093 1340 165659 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 166181 298854 166747 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 166181 1340 166747 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 167269 298854 167835 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 167269 1340 167835 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 168357 298854 168923 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 168357 1340 168923 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 169445 298854 170011 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 169445 1340 170011 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 170533 298854 171099 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 170533 1340 171099 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 171621 298854 172187 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 171621 1340 172187 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 172709 298854 173275 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 172709 1340 173275 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 173797 298854 174363 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 173797 1340 174363 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 174885 298854 175451 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 174885 1340 175451 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 175973 298854 176539 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 175973 1340 176539 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 177061 298854 177627 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 177061 1340 177627 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 178149 298854 178715 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 178149 1340 178715 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 179237 298854 179803 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 179237 1340 179803 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 180325 298854 180891 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 180325 1340 180891 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 181413 298854 181979 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 181413 1340 181979 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 182501 298854 183067 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 182501 1340 183067 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 183589 298854 184155 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 183589 1340 184155 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 184677 298854 185243 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 184677 1340 185243 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 185765 298854 186331 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 185765 1340 186331 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 186853 298854 187419 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 186853 1340 187419 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 187941 298854 188507 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 187941 1340 188507 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 189029 298854 189595 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 189029 1340 189595 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 190117 298854 190683 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 190117 1340 190683 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 191205 298854 191771 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 191205 1340 191771 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 192293 298854 192859 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 192293 1340 192859 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 193381 298854 193947 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 193381 1340 193947 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 194469 298854 195035 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 194469 1340 195035 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 195557 298854 196123 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 195557 1340 196123 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 196645 298854 197211 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 196645 1340 197211 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 197733 298854 198299 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 197733 1340 198299 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 198821 298854 199387 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 198821 1340 199387 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 199909 298854 200475 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 199909 1340 200475 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 200997 298854 201563 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 200997 1340 201563 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 202085 298854 202651 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 202085 1340 202651 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 203173 298854 203739 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 203173 1340 203739 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 204261 298854 204827 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 204261 1340 204827 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 205349 298854 205915 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 205349 1340 205915 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 206437 298854 207003 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 206437 1340 207003 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 207525 298854 208091 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 207525 1340 208091 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 208613 298854 209179 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 208613 1340 209179 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 209701 298854 210267 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 209701 1340 210267 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 210789 298854 211355 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 210789 1340 211355 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 211877 298854 212443 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 211877 1340 212443 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 212965 298854 213531 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 212965 1340 213531 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 214053 298854 214619 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 214053 1340 214619 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 215141 298854 215707 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 215141 1340 215707 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 216229 298854 216795 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 216229 1340 216795 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 217317 298854 217883 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 217317 1340 217883 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 218405 298854 218971 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 218405 1340 218971 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 219493 298854 220059 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 219493 1340 220059 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 220581 298854 221147 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 220581 1340 221147 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 221669 298854 222235 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 221669 1340 222235 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 222757 298854 223323 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 222757 1340 223323 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 223845 298854 224411 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 223845 1340 224411 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 224933 298854 225499 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 224933 1340 225499 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 226021 298854 226587 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 226021 1340 226587 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 227109 298854 227675 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 227109 1340 227675 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 228197 298854 228763 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 228197 1340 228763 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 229285 298854 229851 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 229285 1340 229851 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 230373 298854 230939 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 230373 1340 230939 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 231461 298854 232027 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 231461 1340 232027 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 232549 298854 233115 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 232549 1340 233115 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 233637 298854 234203 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 233637 1340 234203 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 234725 298854 235291 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 234725 1340 235291 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 235813 298854 236379 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 235813 1340 236379 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 236901 298854 237467 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 236901 1340 237467 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 237989 298854 238555 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 237989 1340 238555 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 239077 298854 239643 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 239077 1340 239643 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 240165 298854 240731 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 240165 1340 240731 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 241253 298854 241819 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 241253 1340 241819 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 242341 298854 242907 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 242341 1340 242907 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 243429 298854 243995 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 243429 1340 243995 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 244517 298854 245083 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 244517 1340 245083 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 245605 298854 246171 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 245605 1340 246171 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 246693 298854 247259 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 246693 1340 247259 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 247781 298854 248347 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 247781 1340 248347 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 248869 298854 249435 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 248869 1340 249435 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 249957 298854 250523 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 249957 1340 250523 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 251045 298854 251611 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 251045 1340 251611 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 252133 298854 252699 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 252133 1340 252699 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 253221 298854 253787 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 253221 1340 253787 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 254309 298854 254875 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 254309 1340 254875 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 255397 298854 255963 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 255397 1340 255963 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 256485 298854 257051 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 256485 1340 257051 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 257573 298854 258139 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 257573 1340 258139 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 258661 298854 259227 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 258661 1340 259227 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 259749 298854 260315 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 259749 1340 260315 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 260837 298854 261403 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 260837 1340 261403 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 261925 298854 262491 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 261925 1340 262491 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 263013 298854 263579 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 263013 1340 263579 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 264101 298854 264667 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 264101 1340 264667 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 265189 298854 265755 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 265189 1340 265755 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 266277 298854 266843 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 266277 1340 266843 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 267365 298854 267931 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 267365 1340 267931 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 268453 298854 269019 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 268453 1340 269019 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 269541 298854 270107 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 269541 1340 270107 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 270629 298854 271195 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 270629 1340 271195 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 271717 298854 272283 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 271717 1340 272283 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 272805 298854 273371 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 272805 1340 273371 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 273893 298854 274459 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 273893 1340 274459 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 274981 298854 275547 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 274981 1340 275547 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 276069 298854 276635 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 276069 1340 276635 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 277157 298854 277723 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 277157 1340 277723 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 278245 298854 278811 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 278245 1340 278811 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 279333 298854 279899 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 279333 1340 279899 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 280421 298854 280987 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 280421 1340 280987 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 281509 298854 282075 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 281509 1340 282075 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 282597 298854 283163 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 282597 1340 283163 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 283685 298854 284251 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 283685 1340 284251 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 284773 298854 285339 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 284773 1340 285339 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 285861 298854 286427 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 285861 1340 286427 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 286949 298854 287515 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 286949 1340 287515 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 288037 298854 288603 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 288037 1340 288603 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 289125 298854 289691 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 289125 1340 289691 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 290213 298854 290779 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 290213 1340 290779 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 291301 298854 291867 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 291301 1340 291867 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 292389 298854 292955 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 292389 1340 292955 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 293477 298854 294043 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 293477 1340 294043 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 294565 298854 295131 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 294565 1340 295131 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 295653 298854 296219 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 295653 1340 296219 6 VPWR
port 613 nsew power input
rlabel nwell s 298660 296741 298854 297307 6 VPWR
port 613 nsew power input
rlabel nwell s 1066 296741 1340 297307 6 VPWR
port 613 nsew power input
rlabel metal5 s 299456 934 300056 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 296688 934 297008 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 265968 934 266288 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 235248 934 235568 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 204528 934 204848 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 173808 934 174128 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 143088 934 143408 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 112368 934 112688 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 81648 934 81968 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 50928 934 51248 936 6 VGND
port 614 nsew ground input
rlabel metal5 s 20208 934 20528 936 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 934 464 936 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 936 300056 1340 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 1340 300056 1536 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 1340 1340 1536 6 VGND
port 614 nsew ground input
rlabel metal5 s 299456 1536 300056 1538 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 1536 464 1538 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 13645 300056 13965 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 13645 1340 13965 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 28963 300056 29283 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 28963 1340 29283 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 44281 300056 44601 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 44281 1340 44601 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 59599 300056 59919 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 59599 1340 59919 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 74917 300056 75237 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 74917 1340 75237 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 90235 300056 90555 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 90235 1340 90555 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 105553 300056 105873 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 105553 1340 105873 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 120871 300056 121191 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 120871 1340 121191 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 136189 300056 136509 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 136189 1340 136509 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 151507 300056 151827 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 151507 1340 151827 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 166825 300056 167145 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 166825 1340 167145 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 182143 300056 182463 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 182143 1340 182463 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 197461 300056 197781 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 197461 1340 197781 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 212779 300056 213099 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 212779 1340 213099 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 228097 300056 228417 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 228097 1340 228417 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 243415 300056 243735 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 243415 1340 243735 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 258733 300056 259053 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 258733 1340 259053 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 274051 300056 274371 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 274051 1340 274371 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 289369 300056 289689 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 289369 1340 289689 6 VGND
port 614 nsew ground input
rlabel metal5 s 299456 298206 300056 298208 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 298206 464 298208 6 VGND
port 614 nsew ground input
rlabel metal5 s 298660 298208 300056 298660 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 298208 1340 298660 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 298660 300056 298808 6 VGND
port 614 nsew ground input
rlabel metal5 s 299456 298808 300056 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 296688 298808 297008 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 265968 298808 266288 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 235248 298808 235568 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 204528 298808 204848 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 173808 298808 174128 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 143088 298808 143408 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 112368 298808 112688 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 81648 298808 81968 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 50928 298808 51248 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s 20208 298808 20528 298810 6 VGND
port 614 nsew ground input
rlabel metal5 s -136 298808 464 298810 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 958 299874 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 1278 299874 1514 6 VGND
port 614 nsew ground input
rlabel via4 s 296730 958 296966 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 296730 1278 296966 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 266010 958 266246 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 266010 1278 266246 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 235290 958 235526 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 235290 1278 235526 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 204570 958 204806 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 204570 1278 204806 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 173850 958 174086 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 173850 1278 174086 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 143130 958 143366 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 143130 1278 143366 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 112410 958 112646 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 112410 1278 112646 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 81690 958 81926 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 81690 1278 81926 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 50970 958 51206 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 50970 1278 51206 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 20250 958 20486 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 20250 1278 20486 1340 6 VGND
port 614 nsew ground input
rlabel via4 s 46 958 282 1194 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 13687 299874 13923 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 29005 299874 29241 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 44323 299874 44559 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 59641 299874 59877 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 74959 299874 75195 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 90277 299874 90513 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 105595 299874 105831 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 120913 299874 121149 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 136231 299874 136467 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 151549 299874 151785 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 166867 299874 167103 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 182185 299874 182421 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 197503 299874 197739 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 212821 299874 213057 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 228139 299874 228375 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 243457 299874 243693 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 258775 299874 259011 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 274093 299874 274329 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 289411 299874 289647 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 298230 299874 298466 6 VGND
port 614 nsew ground input
rlabel via4 s 299638 298550 299874 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 46 1278 282 1514 6 VGND
port 614 nsew ground input
rlabel via4 s 46 13687 282 13923 6 VGND
port 614 nsew ground input
rlabel via4 s 46 29005 282 29241 6 VGND
port 614 nsew ground input
rlabel via4 s 46 44323 282 44559 6 VGND
port 614 nsew ground input
rlabel via4 s 46 59641 282 59877 6 VGND
port 614 nsew ground input
rlabel via4 s 46 74959 282 75195 6 VGND
port 614 nsew ground input
rlabel via4 s 46 90277 282 90513 6 VGND
port 614 nsew ground input
rlabel via4 s 46 105595 282 105831 6 VGND
port 614 nsew ground input
rlabel via4 s 46 120913 282 121149 6 VGND
port 614 nsew ground input
rlabel via4 s 46 136231 282 136467 6 VGND
port 614 nsew ground input
rlabel via4 s 46 151549 282 151785 6 VGND
port 614 nsew ground input
rlabel via4 s 46 166867 282 167103 6 VGND
port 614 nsew ground input
rlabel via4 s 46 182185 282 182421 6 VGND
port 614 nsew ground input
rlabel via4 s 46 197503 282 197739 6 VGND
port 614 nsew ground input
rlabel via4 s 46 212821 282 213057 6 VGND
port 614 nsew ground input
rlabel via4 s 46 228139 282 228375 6 VGND
port 614 nsew ground input
rlabel via4 s 46 243457 282 243693 6 VGND
port 614 nsew ground input
rlabel via4 s 46 258775 282 259011 6 VGND
port 614 nsew ground input
rlabel via4 s 46 274093 282 274329 6 VGND
port 614 nsew ground input
rlabel via4 s 46 289411 282 289647 6 VGND
port 614 nsew ground input
rlabel via4 s 46 298230 282 298466 6 VGND
port 614 nsew ground input
rlabel via4 s 296730 298660 296966 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 266010 298660 266246 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 235290 298660 235526 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 204570 298660 204806 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 173850 298660 174086 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 143130 298660 143366 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 112410 298660 112646 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 81690 298660 81926 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 50970 298660 51206 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 20250 298660 20486 298786 6 VGND
port 614 nsew ground input
rlabel via4 s 46 298550 282 298786 6 VGND
port 614 nsew ground input
rlabel metal4 s 299456 936 300056 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 296688 936 297008 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 265968 936 266288 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 235248 936 235568 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 204528 936 204848 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 173808 936 174128 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 143088 936 143408 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 112368 936 112688 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 81648 936 81968 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 50928 936 51248 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 20208 936 20528 1340 6 VGND
port 614 nsew ground input
rlabel metal4 s 296688 298660 297008 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 265968 298660 266288 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 235248 298660 235568 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 204528 298660 204848 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 173808 298660 174128 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 143088 298660 143408 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 112368 298660 112688 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 81648 298660 81968 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 50928 298660 51248 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s 20208 298660 20528 298808 6 VGND
port 614 nsew ground input
rlabel metal4 s -136 936 464 298808 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 2672 298816 2768 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 2672 1340 2768 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 3760 298816 3856 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 3760 1340 3856 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 4848 298816 4944 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 4848 1340 4944 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 5936 298816 6032 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 5936 1340 6032 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 7024 298816 7120 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 7024 1340 7120 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 8112 298816 8208 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 8112 1340 8208 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 9200 298816 9296 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 9200 1340 9296 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 10288 298816 10384 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 10288 1340 10384 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 11376 298816 11472 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 11376 1340 11472 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 12464 298816 12560 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 12464 1340 12560 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 13552 298816 13648 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 13552 1340 13648 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 14640 298816 14736 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 14640 1340 14736 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 15728 298816 15824 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 15728 1340 15824 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 16816 298816 16912 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 16816 1340 16912 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 17904 298816 18000 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 17904 1340 18000 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 18992 298816 19088 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 18992 1340 19088 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 20080 298816 20176 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 20080 1340 20176 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 21168 298816 21264 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 21168 1340 21264 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 22256 298816 22352 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 22256 1340 22352 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 23344 298816 23440 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 23344 1340 23440 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 24432 298816 24528 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 24432 1340 24528 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 25520 298816 25616 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 25520 1340 25616 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 26608 298816 26704 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 26608 1340 26704 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 27696 298816 27792 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 27696 1340 27792 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 28784 298816 28880 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 28784 1340 28880 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 29872 298816 29968 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 29872 1340 29968 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 30960 298816 31056 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 30960 1340 31056 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 32048 298816 32144 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 32048 1340 32144 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 33136 298816 33232 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 33136 1340 33232 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 34224 298816 34320 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 34224 1340 34320 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 35312 298816 35408 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 35312 1340 35408 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 36400 298816 36496 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 36400 1340 36496 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 37488 298816 37584 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 37488 1340 37584 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 38576 298816 38672 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 38576 1340 38672 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 39664 298816 39760 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 39664 1340 39760 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 40752 298816 40848 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 40752 1340 40848 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 41840 298816 41936 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 41840 1340 41936 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 42928 298816 43024 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 42928 1340 43024 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 44016 298816 44112 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 44016 1340 44112 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 45104 298816 45200 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 45104 1340 45200 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 46192 298816 46288 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 46192 1340 46288 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 47280 298816 47376 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 47280 1340 47376 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 48368 298816 48464 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 48368 1340 48464 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 49456 298816 49552 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 49456 1340 49552 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 50544 298816 50640 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 50544 1340 50640 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 51632 298816 51728 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 51632 1340 51728 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 52720 298816 52816 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 52720 1340 52816 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 53808 298816 53904 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 53808 1340 53904 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 54896 298816 54992 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 54896 1340 54992 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 55984 298816 56080 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 55984 1340 56080 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 57072 298816 57168 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 57072 1340 57168 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 58160 298816 58256 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 58160 1340 58256 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 59248 298816 59344 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 59248 1340 59344 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 60336 298816 60432 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 60336 1340 60432 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 61424 298816 61520 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 61424 1340 61520 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 62512 298816 62608 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 62512 1340 62608 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 63600 298816 63696 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 63600 1340 63696 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 64688 298816 64784 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 64688 1340 64784 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 65776 298816 65872 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 65776 1340 65872 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 66864 298816 66960 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 66864 1340 66960 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 67952 298816 68048 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 67952 1340 68048 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 69040 298816 69136 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 69040 1340 69136 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 70128 298816 70224 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 70128 1340 70224 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 71216 298816 71312 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 71216 1340 71312 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 72304 298816 72400 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 72304 1340 72400 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 73392 298816 73488 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 73392 1340 73488 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 74480 298816 74576 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 74480 1340 74576 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 75568 298816 75664 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 75568 1340 75664 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 76656 298816 76752 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 76656 1340 76752 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 77744 298816 77840 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 77744 1340 77840 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 78832 298816 78928 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 78832 1340 78928 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 79920 298816 80016 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 79920 1340 80016 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 81008 298816 81104 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 81008 1340 81104 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 82096 298816 82192 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 82096 1340 82192 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 83184 298816 83280 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 83184 1340 83280 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 84272 298816 84368 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 84272 1340 84368 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 85360 298816 85456 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 85360 1340 85456 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 86448 298816 86544 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 86448 1340 86544 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 87536 298816 87632 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 87536 1340 87632 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 88624 298816 88720 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 88624 1340 88720 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 89712 298816 89808 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 89712 1340 89808 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 90800 298816 90896 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 90800 1340 90896 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 91888 298816 91984 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 91888 1340 91984 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 92976 298816 93072 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 92976 1340 93072 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 94064 298816 94160 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 94064 1340 94160 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 95152 298816 95248 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 95152 1340 95248 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 96240 298816 96336 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 96240 1340 96336 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 97328 298816 97424 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 97328 1340 97424 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 98416 298816 98512 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 98416 1340 98512 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 99504 298816 99600 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 99504 1340 99600 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 100592 298816 100688 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 100592 1340 100688 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 101680 298816 101776 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 101680 1340 101776 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 102768 298816 102864 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 102768 1340 102864 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 103856 298816 103952 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 103856 1340 103952 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 104944 298816 105040 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 104944 1340 105040 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 106032 298816 106128 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 106032 1340 106128 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 107120 298816 107216 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 107120 1340 107216 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 108208 298816 108304 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 108208 1340 108304 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 109296 298816 109392 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 109296 1340 109392 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 110384 298816 110480 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 110384 1340 110480 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 111472 298816 111568 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 111472 1340 111568 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 112560 298816 112656 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 112560 1340 112656 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 113648 298816 113744 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 113648 1340 113744 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 114736 298816 114832 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 114736 1340 114832 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 115824 298816 115920 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 115824 1340 115920 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 116912 298816 117008 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 116912 1340 117008 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 118000 298816 118096 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 118000 1340 118096 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 119088 298816 119184 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 119088 1340 119184 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 120176 298816 120272 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 120176 1340 120272 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 121264 298816 121360 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 121264 1340 121360 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 122352 298816 122448 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 122352 1340 122448 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 123440 298816 123536 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 123440 1340 123536 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 124528 298816 124624 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 124528 1340 124624 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 125616 298816 125712 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 125616 1340 125712 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 126704 298816 126800 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 126704 1340 126800 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 127792 298816 127888 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 127792 1340 127888 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 128880 298816 128976 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 128880 1340 128976 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 129968 298816 130064 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 129968 1340 130064 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 131056 298816 131152 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 131056 1340 131152 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 132144 298816 132240 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 132144 1340 132240 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 133232 298816 133328 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 133232 1340 133328 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 134320 298816 134416 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 134320 1340 134416 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 135408 298816 135504 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 135408 1340 135504 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 136496 298816 136592 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 136496 1340 136592 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 137584 298816 137680 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 137584 1340 137680 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 138672 298816 138768 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 138672 1340 138768 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 139760 298816 139856 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 139760 1340 139856 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 140848 298816 140944 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 140848 1340 140944 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 141936 298816 142032 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 141936 1340 142032 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 143024 298816 143120 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 143024 1340 143120 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 144112 298816 144208 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 144112 1340 144208 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 145200 298816 145296 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 145200 1340 145296 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 146288 298816 146384 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 146288 1340 146384 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 147376 298816 147472 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 147376 1340 147472 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 148464 298816 148560 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 148464 1340 148560 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 149552 298816 149648 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 149552 1340 149648 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 150640 298816 150736 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 150640 1340 150736 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 151728 298816 151824 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 151728 1340 151824 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 152816 298816 152912 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 152816 1340 152912 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 153904 298816 154000 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 153904 1340 154000 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 154992 298816 155088 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 154992 1340 155088 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 156080 298816 156176 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 156080 1340 156176 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 157168 298816 157264 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 157168 1340 157264 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 158256 298816 158352 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 158256 1340 158352 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 159344 298816 159440 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 159344 1340 159440 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 160432 298816 160528 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 160432 1340 160528 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 161520 298816 161616 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 161520 1340 161616 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 162608 298816 162704 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 162608 1340 162704 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 163696 298816 163792 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 163696 1340 163792 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 164784 298816 164880 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 164784 1340 164880 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 165872 298816 165968 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 165872 1340 165968 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 166960 298816 167056 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 166960 1340 167056 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 168048 298816 168144 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 168048 1340 168144 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 169136 298816 169232 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 169136 1340 169232 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 170224 298816 170320 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 170224 1340 170320 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 171312 298816 171408 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 171312 1340 171408 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 172400 298816 172496 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 172400 1340 172496 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 173488 298816 173584 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 173488 1340 173584 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 174576 298816 174672 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 174576 1340 174672 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 175664 298816 175760 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 175664 1340 175760 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 176752 298816 176848 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 176752 1340 176848 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 177840 298816 177936 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 177840 1340 177936 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 178928 298816 179024 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 178928 1340 179024 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 180016 298816 180112 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 180016 1340 180112 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 181104 298816 181200 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 181104 1340 181200 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 182192 298816 182288 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 182192 1340 182288 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 183280 298816 183376 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 183280 1340 183376 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 184368 298816 184464 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 184368 1340 184464 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 185456 298816 185552 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 185456 1340 185552 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 186544 298816 186640 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 186544 1340 186640 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 187632 298816 187728 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 187632 1340 187728 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 188720 298816 188816 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 188720 1340 188816 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 189808 298816 189904 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 189808 1340 189904 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 190896 298816 190992 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 190896 1340 190992 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 191984 298816 192080 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 191984 1340 192080 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 193072 298816 193168 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 193072 1340 193168 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 194160 298816 194256 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 194160 1340 194256 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 195248 298816 195344 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 195248 1340 195344 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 196336 298816 196432 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 196336 1340 196432 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 197424 298816 197520 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 197424 1340 197520 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 198512 298816 198608 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 198512 1340 198608 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 199600 298816 199696 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 199600 1340 199696 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 200688 298816 200784 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 200688 1340 200784 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 201776 298816 201872 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 201776 1340 201872 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 202864 298816 202960 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 202864 1340 202960 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 203952 298816 204048 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 203952 1340 204048 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 205040 298816 205136 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 205040 1340 205136 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 206128 298816 206224 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 206128 1340 206224 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 207216 298816 207312 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 207216 1340 207312 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 208304 298816 208400 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 208304 1340 208400 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 209392 298816 209488 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 209392 1340 209488 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 210480 298816 210576 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 210480 1340 210576 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 211568 298816 211664 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 211568 1340 211664 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 212656 298816 212752 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 212656 1340 212752 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 213744 298816 213840 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 213744 1340 213840 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 214832 298816 214928 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 214832 1340 214928 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 215920 298816 216016 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 215920 1340 216016 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 217008 298816 217104 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 217008 1340 217104 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 218096 298816 218192 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 218096 1340 218192 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 219184 298816 219280 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 219184 1340 219280 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 220272 298816 220368 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 220272 1340 220368 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 221360 298816 221456 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 221360 1340 221456 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 222448 298816 222544 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 222448 1340 222544 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 223536 298816 223632 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 223536 1340 223632 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 224624 298816 224720 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 224624 1340 224720 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 225712 298816 225808 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 225712 1340 225808 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 226800 298816 226896 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 226800 1340 226896 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 227888 298816 227984 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 227888 1340 227984 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 228976 298816 229072 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 228976 1340 229072 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 230064 298816 230160 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 230064 1340 230160 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 231152 298816 231248 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 231152 1340 231248 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 232240 298816 232336 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 232240 1340 232336 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 233328 298816 233424 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 233328 1340 233424 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 234416 298816 234512 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 234416 1340 234512 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 235504 298816 235600 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 235504 1340 235600 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 236592 298816 236688 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 236592 1340 236688 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 237680 298816 237776 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 237680 1340 237776 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 238768 298816 238864 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 238768 1340 238864 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 239856 298816 239952 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 239856 1340 239952 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 240944 298816 241040 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 240944 1340 241040 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 242032 298816 242128 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 242032 1340 242128 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 243120 298816 243216 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 243120 1340 243216 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 244208 298816 244304 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 244208 1340 244304 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 245296 298816 245392 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 245296 1340 245392 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 246384 298816 246480 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 246384 1340 246480 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 247472 298816 247568 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 247472 1340 247568 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 248560 298816 248656 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 248560 1340 248656 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 249648 298816 249744 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 249648 1340 249744 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 250736 298816 250832 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 250736 1340 250832 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 251824 298816 251920 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 251824 1340 251920 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 252912 298816 253008 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 252912 1340 253008 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 254000 298816 254096 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 254000 1340 254096 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 255088 298816 255184 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 255088 1340 255184 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 256176 298816 256272 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 256176 1340 256272 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 257264 298816 257360 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 257264 1340 257360 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 258352 298816 258448 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 258352 1340 258448 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 259440 298816 259536 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 259440 1340 259536 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 260528 298816 260624 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 260528 1340 260624 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 261616 298816 261712 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 261616 1340 261712 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 262704 298816 262800 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 262704 1340 262800 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 263792 298816 263888 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 263792 1340 263888 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 264880 298816 264976 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 264880 1340 264976 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 265968 298816 266064 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 265968 1340 266064 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 267056 298816 267152 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 267056 1340 267152 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 268144 298816 268240 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 268144 1340 268240 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 269232 298816 269328 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 269232 1340 269328 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 270320 298816 270416 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 270320 1340 270416 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 271408 298816 271504 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 271408 1340 271504 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 272496 298816 272592 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 272496 1340 272592 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 273584 298816 273680 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 273584 1340 273680 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 274672 298816 274768 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 274672 1340 274768 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 275760 298816 275856 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 275760 1340 275856 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 276848 298816 276944 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 276848 1340 276944 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 277936 298816 278032 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 277936 1340 278032 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 279024 298816 279120 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 279024 1340 279120 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 280112 298816 280208 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 280112 1340 280208 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 281200 298816 281296 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 281200 1340 281296 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 282288 298816 282384 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 282288 1340 282384 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 283376 298816 283472 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 283376 1340 283472 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 284464 298816 284560 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 284464 1340 284560 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 285552 298816 285648 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 285552 1340 285648 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 286640 298816 286736 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 286640 1340 286736 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 287728 298816 287824 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 287728 1340 287824 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 288816 298816 288912 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 288816 1340 288912 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 289904 298816 290000 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 289904 1340 290000 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 290992 298816 291088 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 290992 1340 291088 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 292080 298816 292176 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 292080 1340 292176 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 293168 298816 293264 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 293168 1340 293264 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 294256 298816 294352 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 294256 1340 294352 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 295344 298816 295440 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 295344 1340 295440 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 296432 298816 296528 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 296432 1340 296528 6 VGND
port 614 nsew ground input
rlabel metal1 s 298660 297520 298816 297616 6 VGND
port 614 nsew ground input
rlabel metal1 s 1104 297520 1340 297616 6 VGND
port 614 nsew ground input
rlabel viali s 298753 2703 298787 2737 6 VGND
port 614 nsew ground input
rlabel viali s 298661 2703 298695 2737 6 VGND
port 614 nsew ground input
rlabel viali s 1317 2703 1340 2737 6 VGND
port 614 nsew ground input
rlabel viali s 1225 2703 1259 2737 6 VGND
port 614 nsew ground input
rlabel viali s 1133 2703 1167 2737 6 VGND
port 614 nsew ground input
rlabel viali s 298753 3791 298787 3825 6 VGND
port 614 nsew ground input
rlabel viali s 298661 3791 298695 3825 6 VGND
port 614 nsew ground input
rlabel viali s 1317 3791 1340 3825 6 VGND
port 614 nsew ground input
rlabel viali s 1225 3791 1259 3825 6 VGND
port 614 nsew ground input
rlabel viali s 1133 3791 1167 3825 6 VGND
port 614 nsew ground input
rlabel viali s 298753 4879 298787 4913 6 VGND
port 614 nsew ground input
rlabel viali s 298661 4879 298695 4913 6 VGND
port 614 nsew ground input
rlabel viali s 1317 4879 1340 4913 6 VGND
port 614 nsew ground input
rlabel viali s 1225 4879 1259 4913 6 VGND
port 614 nsew ground input
rlabel viali s 1133 4879 1167 4913 6 VGND
port 614 nsew ground input
rlabel viali s 298753 5967 298787 6001 6 VGND
port 614 nsew ground input
rlabel viali s 298661 5967 298695 6001 6 VGND
port 614 nsew ground input
rlabel viali s 1317 5967 1340 6001 6 VGND
port 614 nsew ground input
rlabel viali s 1225 5967 1259 6001 6 VGND
port 614 nsew ground input
rlabel viali s 1133 5967 1167 6001 6 VGND
port 614 nsew ground input
rlabel viali s 298753 7055 298787 7089 6 VGND
port 614 nsew ground input
rlabel viali s 298661 7055 298695 7089 6 VGND
port 614 nsew ground input
rlabel viali s 1317 7055 1340 7089 6 VGND
port 614 nsew ground input
rlabel viali s 1225 7055 1259 7089 6 VGND
port 614 nsew ground input
rlabel viali s 1133 7055 1167 7089 6 VGND
port 614 nsew ground input
rlabel viali s 298753 8143 298787 8177 6 VGND
port 614 nsew ground input
rlabel viali s 298661 8143 298695 8177 6 VGND
port 614 nsew ground input
rlabel viali s 1317 8143 1340 8177 6 VGND
port 614 nsew ground input
rlabel viali s 1225 8143 1259 8177 6 VGND
port 614 nsew ground input
rlabel viali s 1133 8143 1167 8177 6 VGND
port 614 nsew ground input
rlabel viali s 298753 9231 298787 9265 6 VGND
port 614 nsew ground input
rlabel viali s 298661 9231 298695 9265 6 VGND
port 614 nsew ground input
rlabel viali s 1317 9231 1340 9265 6 VGND
port 614 nsew ground input
rlabel viali s 1225 9231 1259 9265 6 VGND
port 614 nsew ground input
rlabel viali s 1133 9231 1167 9265 6 VGND
port 614 nsew ground input
rlabel viali s 298753 10319 298787 10353 6 VGND
port 614 nsew ground input
rlabel viali s 298661 10319 298695 10353 6 VGND
port 614 nsew ground input
rlabel viali s 1317 10319 1340 10353 6 VGND
port 614 nsew ground input
rlabel viali s 1225 10319 1259 10353 6 VGND
port 614 nsew ground input
rlabel viali s 1133 10319 1167 10353 6 VGND
port 614 nsew ground input
rlabel viali s 298753 11407 298787 11441 6 VGND
port 614 nsew ground input
rlabel viali s 298661 11407 298695 11441 6 VGND
port 614 nsew ground input
rlabel viali s 1317 11407 1340 11441 6 VGND
port 614 nsew ground input
rlabel viali s 1225 11407 1259 11441 6 VGND
port 614 nsew ground input
rlabel viali s 1133 11407 1167 11441 6 VGND
port 614 nsew ground input
rlabel viali s 298753 12495 298787 12529 6 VGND
port 614 nsew ground input
rlabel viali s 298661 12495 298695 12529 6 VGND
port 614 nsew ground input
rlabel viali s 1317 12495 1340 12529 6 VGND
port 614 nsew ground input
rlabel viali s 1225 12495 1259 12529 6 VGND
port 614 nsew ground input
rlabel viali s 1133 12495 1167 12529 6 VGND
port 614 nsew ground input
rlabel viali s 298753 13583 298787 13617 6 VGND
port 614 nsew ground input
rlabel viali s 298661 13583 298695 13617 6 VGND
port 614 nsew ground input
rlabel viali s 1317 13583 1340 13617 6 VGND
port 614 nsew ground input
rlabel viali s 1225 13583 1259 13617 6 VGND
port 614 nsew ground input
rlabel viali s 1133 13583 1167 13617 6 VGND
port 614 nsew ground input
rlabel viali s 298753 14671 298787 14705 6 VGND
port 614 nsew ground input
rlabel viali s 298661 14671 298695 14705 6 VGND
port 614 nsew ground input
rlabel viali s 1317 14671 1340 14705 6 VGND
port 614 nsew ground input
rlabel viali s 1225 14671 1259 14705 6 VGND
port 614 nsew ground input
rlabel viali s 1133 14671 1167 14705 6 VGND
port 614 nsew ground input
rlabel viali s 298753 15759 298787 15793 6 VGND
port 614 nsew ground input
rlabel viali s 298661 15759 298695 15793 6 VGND
port 614 nsew ground input
rlabel viali s 1317 15759 1340 15793 6 VGND
port 614 nsew ground input
rlabel viali s 1225 15759 1259 15793 6 VGND
port 614 nsew ground input
rlabel viali s 1133 15759 1167 15793 6 VGND
port 614 nsew ground input
rlabel viali s 298753 16847 298787 16881 6 VGND
port 614 nsew ground input
rlabel viali s 298661 16847 298695 16881 6 VGND
port 614 nsew ground input
rlabel viali s 1317 16847 1340 16881 6 VGND
port 614 nsew ground input
rlabel viali s 1225 16847 1259 16881 6 VGND
port 614 nsew ground input
rlabel viali s 1133 16847 1167 16881 6 VGND
port 614 nsew ground input
rlabel viali s 298753 17935 298787 17969 6 VGND
port 614 nsew ground input
rlabel viali s 298661 17935 298695 17969 6 VGND
port 614 nsew ground input
rlabel viali s 1317 17935 1340 17969 6 VGND
port 614 nsew ground input
rlabel viali s 1225 17935 1259 17969 6 VGND
port 614 nsew ground input
rlabel viali s 1133 17935 1167 17969 6 VGND
port 614 nsew ground input
rlabel viali s 298753 19023 298787 19057 6 VGND
port 614 nsew ground input
rlabel viali s 298661 19023 298695 19057 6 VGND
port 614 nsew ground input
rlabel viali s 1317 19023 1340 19057 6 VGND
port 614 nsew ground input
rlabel viali s 1225 19023 1259 19057 6 VGND
port 614 nsew ground input
rlabel viali s 1133 19023 1167 19057 6 VGND
port 614 nsew ground input
rlabel viali s 298753 20111 298787 20145 6 VGND
port 614 nsew ground input
rlabel viali s 298661 20111 298695 20145 6 VGND
port 614 nsew ground input
rlabel viali s 1317 20111 1340 20145 6 VGND
port 614 nsew ground input
rlabel viali s 1225 20111 1259 20145 6 VGND
port 614 nsew ground input
rlabel viali s 1133 20111 1167 20145 6 VGND
port 614 nsew ground input
rlabel viali s 298753 21199 298787 21233 6 VGND
port 614 nsew ground input
rlabel viali s 298661 21199 298695 21233 6 VGND
port 614 nsew ground input
rlabel viali s 1317 21199 1340 21233 6 VGND
port 614 nsew ground input
rlabel viali s 1225 21199 1259 21233 6 VGND
port 614 nsew ground input
rlabel viali s 1133 21199 1167 21233 6 VGND
port 614 nsew ground input
rlabel viali s 298753 22287 298787 22321 6 VGND
port 614 nsew ground input
rlabel viali s 298661 22287 298695 22321 6 VGND
port 614 nsew ground input
rlabel viali s 1317 22287 1340 22321 6 VGND
port 614 nsew ground input
rlabel viali s 1225 22287 1259 22321 6 VGND
port 614 nsew ground input
rlabel viali s 1133 22287 1167 22321 6 VGND
port 614 nsew ground input
rlabel viali s 298753 23375 298787 23409 6 VGND
port 614 nsew ground input
rlabel viali s 298661 23375 298695 23409 6 VGND
port 614 nsew ground input
rlabel viali s 1317 23375 1340 23409 6 VGND
port 614 nsew ground input
rlabel viali s 1225 23375 1259 23409 6 VGND
port 614 nsew ground input
rlabel viali s 1133 23375 1167 23409 6 VGND
port 614 nsew ground input
rlabel viali s 298753 24463 298787 24497 6 VGND
port 614 nsew ground input
rlabel viali s 298661 24463 298695 24497 6 VGND
port 614 nsew ground input
rlabel viali s 1317 24463 1340 24497 6 VGND
port 614 nsew ground input
rlabel viali s 1225 24463 1259 24497 6 VGND
port 614 nsew ground input
rlabel viali s 1133 24463 1167 24497 6 VGND
port 614 nsew ground input
rlabel viali s 298753 25551 298787 25585 6 VGND
port 614 nsew ground input
rlabel viali s 298661 25551 298695 25585 6 VGND
port 614 nsew ground input
rlabel viali s 1317 25551 1340 25585 6 VGND
port 614 nsew ground input
rlabel viali s 1225 25551 1259 25585 6 VGND
port 614 nsew ground input
rlabel viali s 1133 25551 1167 25585 6 VGND
port 614 nsew ground input
rlabel viali s 298753 26639 298787 26673 6 VGND
port 614 nsew ground input
rlabel viali s 298661 26639 298695 26673 6 VGND
port 614 nsew ground input
rlabel viali s 1317 26639 1340 26673 6 VGND
port 614 nsew ground input
rlabel viali s 1225 26639 1259 26673 6 VGND
port 614 nsew ground input
rlabel viali s 1133 26639 1167 26673 6 VGND
port 614 nsew ground input
rlabel viali s 298753 27727 298787 27761 6 VGND
port 614 nsew ground input
rlabel viali s 298661 27727 298695 27761 6 VGND
port 614 nsew ground input
rlabel viali s 1317 27727 1340 27761 6 VGND
port 614 nsew ground input
rlabel viali s 1225 27727 1259 27761 6 VGND
port 614 nsew ground input
rlabel viali s 1133 27727 1167 27761 6 VGND
port 614 nsew ground input
rlabel viali s 298753 28815 298787 28849 6 VGND
port 614 nsew ground input
rlabel viali s 298661 28815 298695 28849 6 VGND
port 614 nsew ground input
rlabel viali s 1317 28815 1340 28849 6 VGND
port 614 nsew ground input
rlabel viali s 1225 28815 1259 28849 6 VGND
port 614 nsew ground input
rlabel viali s 1133 28815 1167 28849 6 VGND
port 614 nsew ground input
rlabel viali s 298753 29903 298787 29937 6 VGND
port 614 nsew ground input
rlabel viali s 298661 29903 298695 29937 6 VGND
port 614 nsew ground input
rlabel viali s 1317 29903 1340 29937 6 VGND
port 614 nsew ground input
rlabel viali s 1225 29903 1259 29937 6 VGND
port 614 nsew ground input
rlabel viali s 1133 29903 1167 29937 6 VGND
port 614 nsew ground input
rlabel viali s 298753 30991 298787 31025 6 VGND
port 614 nsew ground input
rlabel viali s 298661 30991 298695 31025 6 VGND
port 614 nsew ground input
rlabel viali s 1317 30991 1340 31025 6 VGND
port 614 nsew ground input
rlabel viali s 1225 30991 1259 31025 6 VGND
port 614 nsew ground input
rlabel viali s 1133 30991 1167 31025 6 VGND
port 614 nsew ground input
rlabel viali s 298753 32079 298787 32113 6 VGND
port 614 nsew ground input
rlabel viali s 298661 32079 298695 32113 6 VGND
port 614 nsew ground input
rlabel viali s 1317 32079 1340 32113 6 VGND
port 614 nsew ground input
rlabel viali s 1225 32079 1259 32113 6 VGND
port 614 nsew ground input
rlabel viali s 1133 32079 1167 32113 6 VGND
port 614 nsew ground input
rlabel viali s 298753 33167 298787 33201 6 VGND
port 614 nsew ground input
rlabel viali s 298661 33167 298695 33201 6 VGND
port 614 nsew ground input
rlabel viali s 1317 33167 1340 33201 6 VGND
port 614 nsew ground input
rlabel viali s 1225 33167 1259 33201 6 VGND
port 614 nsew ground input
rlabel viali s 1133 33167 1167 33201 6 VGND
port 614 nsew ground input
rlabel viali s 298753 34255 298787 34289 6 VGND
port 614 nsew ground input
rlabel viali s 298661 34255 298695 34289 6 VGND
port 614 nsew ground input
rlabel viali s 1317 34255 1340 34289 6 VGND
port 614 nsew ground input
rlabel viali s 1225 34255 1259 34289 6 VGND
port 614 nsew ground input
rlabel viali s 1133 34255 1167 34289 6 VGND
port 614 nsew ground input
rlabel viali s 298753 35343 298787 35377 6 VGND
port 614 nsew ground input
rlabel viali s 298661 35343 298695 35377 6 VGND
port 614 nsew ground input
rlabel viali s 1317 35343 1340 35377 6 VGND
port 614 nsew ground input
rlabel viali s 1225 35343 1259 35377 6 VGND
port 614 nsew ground input
rlabel viali s 1133 35343 1167 35377 6 VGND
port 614 nsew ground input
rlabel viali s 298753 36431 298787 36465 6 VGND
port 614 nsew ground input
rlabel viali s 298661 36431 298695 36465 6 VGND
port 614 nsew ground input
rlabel viali s 1317 36431 1340 36465 6 VGND
port 614 nsew ground input
rlabel viali s 1225 36431 1259 36465 6 VGND
port 614 nsew ground input
rlabel viali s 1133 36431 1167 36465 6 VGND
port 614 nsew ground input
rlabel viali s 298753 37519 298787 37553 6 VGND
port 614 nsew ground input
rlabel viali s 298661 37519 298695 37553 6 VGND
port 614 nsew ground input
rlabel viali s 1317 37519 1340 37553 6 VGND
port 614 nsew ground input
rlabel viali s 1225 37519 1259 37553 6 VGND
port 614 nsew ground input
rlabel viali s 1133 37519 1167 37553 6 VGND
port 614 nsew ground input
rlabel viali s 298753 38607 298787 38641 6 VGND
port 614 nsew ground input
rlabel viali s 298661 38607 298695 38641 6 VGND
port 614 nsew ground input
rlabel viali s 1317 38607 1340 38641 6 VGND
port 614 nsew ground input
rlabel viali s 1225 38607 1259 38641 6 VGND
port 614 nsew ground input
rlabel viali s 1133 38607 1167 38641 6 VGND
port 614 nsew ground input
rlabel viali s 298753 39695 298787 39729 6 VGND
port 614 nsew ground input
rlabel viali s 298661 39695 298695 39729 6 VGND
port 614 nsew ground input
rlabel viali s 1317 39695 1340 39729 6 VGND
port 614 nsew ground input
rlabel viali s 1225 39695 1259 39729 6 VGND
port 614 nsew ground input
rlabel viali s 1133 39695 1167 39729 6 VGND
port 614 nsew ground input
rlabel viali s 298753 40783 298787 40817 6 VGND
port 614 nsew ground input
rlabel viali s 298661 40783 298695 40817 6 VGND
port 614 nsew ground input
rlabel viali s 1317 40783 1340 40817 6 VGND
port 614 nsew ground input
rlabel viali s 1225 40783 1259 40817 6 VGND
port 614 nsew ground input
rlabel viali s 1133 40783 1167 40817 6 VGND
port 614 nsew ground input
rlabel viali s 298753 41871 298787 41905 6 VGND
port 614 nsew ground input
rlabel viali s 298661 41871 298695 41905 6 VGND
port 614 nsew ground input
rlabel viali s 1317 41871 1340 41905 6 VGND
port 614 nsew ground input
rlabel viali s 1225 41871 1259 41905 6 VGND
port 614 nsew ground input
rlabel viali s 1133 41871 1167 41905 6 VGND
port 614 nsew ground input
rlabel viali s 298753 42959 298787 42993 6 VGND
port 614 nsew ground input
rlabel viali s 298661 42959 298695 42993 6 VGND
port 614 nsew ground input
rlabel viali s 1317 42959 1340 42993 6 VGND
port 614 nsew ground input
rlabel viali s 1225 42959 1259 42993 6 VGND
port 614 nsew ground input
rlabel viali s 1133 42959 1167 42993 6 VGND
port 614 nsew ground input
rlabel viali s 298753 44047 298787 44081 6 VGND
port 614 nsew ground input
rlabel viali s 298661 44047 298695 44081 6 VGND
port 614 nsew ground input
rlabel viali s 1317 44047 1340 44081 6 VGND
port 614 nsew ground input
rlabel viali s 1225 44047 1259 44081 6 VGND
port 614 nsew ground input
rlabel viali s 1133 44047 1167 44081 6 VGND
port 614 nsew ground input
rlabel viali s 298753 45135 298787 45169 6 VGND
port 614 nsew ground input
rlabel viali s 298661 45135 298695 45169 6 VGND
port 614 nsew ground input
rlabel viali s 1317 45135 1340 45169 6 VGND
port 614 nsew ground input
rlabel viali s 1225 45135 1259 45169 6 VGND
port 614 nsew ground input
rlabel viali s 1133 45135 1167 45169 6 VGND
port 614 nsew ground input
rlabel viali s 298753 46223 298787 46257 6 VGND
port 614 nsew ground input
rlabel viali s 298661 46223 298695 46257 6 VGND
port 614 nsew ground input
rlabel viali s 1317 46223 1340 46257 6 VGND
port 614 nsew ground input
rlabel viali s 1225 46223 1259 46257 6 VGND
port 614 nsew ground input
rlabel viali s 1133 46223 1167 46257 6 VGND
port 614 nsew ground input
rlabel viali s 298753 47311 298787 47345 6 VGND
port 614 nsew ground input
rlabel viali s 298661 47311 298695 47345 6 VGND
port 614 nsew ground input
rlabel viali s 1317 47311 1340 47345 6 VGND
port 614 nsew ground input
rlabel viali s 1225 47311 1259 47345 6 VGND
port 614 nsew ground input
rlabel viali s 1133 47311 1167 47345 6 VGND
port 614 nsew ground input
rlabel viali s 298753 48399 298787 48433 6 VGND
port 614 nsew ground input
rlabel viali s 298661 48399 298695 48433 6 VGND
port 614 nsew ground input
rlabel viali s 1317 48399 1340 48433 6 VGND
port 614 nsew ground input
rlabel viali s 1225 48399 1259 48433 6 VGND
port 614 nsew ground input
rlabel viali s 1133 48399 1167 48433 6 VGND
port 614 nsew ground input
rlabel viali s 298753 49487 298787 49521 6 VGND
port 614 nsew ground input
rlabel viali s 298661 49487 298695 49521 6 VGND
port 614 nsew ground input
rlabel viali s 1317 49487 1340 49521 6 VGND
port 614 nsew ground input
rlabel viali s 1225 49487 1259 49521 6 VGND
port 614 nsew ground input
rlabel viali s 1133 49487 1167 49521 6 VGND
port 614 nsew ground input
rlabel viali s 298753 50575 298787 50609 6 VGND
port 614 nsew ground input
rlabel viali s 298661 50575 298695 50609 6 VGND
port 614 nsew ground input
rlabel viali s 1317 50575 1340 50609 6 VGND
port 614 nsew ground input
rlabel viali s 1225 50575 1259 50609 6 VGND
port 614 nsew ground input
rlabel viali s 1133 50575 1167 50609 6 VGND
port 614 nsew ground input
rlabel viali s 298753 51663 298787 51697 6 VGND
port 614 nsew ground input
rlabel viali s 298661 51663 298695 51697 6 VGND
port 614 nsew ground input
rlabel viali s 1317 51663 1340 51697 6 VGND
port 614 nsew ground input
rlabel viali s 1225 51663 1259 51697 6 VGND
port 614 nsew ground input
rlabel viali s 1133 51663 1167 51697 6 VGND
port 614 nsew ground input
rlabel viali s 298753 52751 298787 52785 6 VGND
port 614 nsew ground input
rlabel viali s 298661 52751 298695 52785 6 VGND
port 614 nsew ground input
rlabel viali s 1317 52751 1340 52785 6 VGND
port 614 nsew ground input
rlabel viali s 1225 52751 1259 52785 6 VGND
port 614 nsew ground input
rlabel viali s 1133 52751 1167 52785 6 VGND
port 614 nsew ground input
rlabel viali s 298753 53839 298787 53873 6 VGND
port 614 nsew ground input
rlabel viali s 298661 53839 298695 53873 6 VGND
port 614 nsew ground input
rlabel viali s 1317 53839 1340 53873 6 VGND
port 614 nsew ground input
rlabel viali s 1225 53839 1259 53873 6 VGND
port 614 nsew ground input
rlabel viali s 1133 53839 1167 53873 6 VGND
port 614 nsew ground input
rlabel viali s 298753 54927 298787 54961 6 VGND
port 614 nsew ground input
rlabel viali s 298661 54927 298695 54961 6 VGND
port 614 nsew ground input
rlabel viali s 1317 54927 1340 54961 6 VGND
port 614 nsew ground input
rlabel viali s 1225 54927 1259 54961 6 VGND
port 614 nsew ground input
rlabel viali s 1133 54927 1167 54961 6 VGND
port 614 nsew ground input
rlabel viali s 298753 56015 298787 56049 6 VGND
port 614 nsew ground input
rlabel viali s 298661 56015 298695 56049 6 VGND
port 614 nsew ground input
rlabel viali s 1317 56015 1340 56049 6 VGND
port 614 nsew ground input
rlabel viali s 1225 56015 1259 56049 6 VGND
port 614 nsew ground input
rlabel viali s 1133 56015 1167 56049 6 VGND
port 614 nsew ground input
rlabel viali s 298753 57103 298787 57137 6 VGND
port 614 nsew ground input
rlabel viali s 298661 57103 298695 57137 6 VGND
port 614 nsew ground input
rlabel viali s 1317 57103 1340 57137 6 VGND
port 614 nsew ground input
rlabel viali s 1225 57103 1259 57137 6 VGND
port 614 nsew ground input
rlabel viali s 1133 57103 1167 57137 6 VGND
port 614 nsew ground input
rlabel viali s 298753 58191 298787 58225 6 VGND
port 614 nsew ground input
rlabel viali s 298661 58191 298695 58225 6 VGND
port 614 nsew ground input
rlabel viali s 1317 58191 1340 58225 6 VGND
port 614 nsew ground input
rlabel viali s 1225 58191 1259 58225 6 VGND
port 614 nsew ground input
rlabel viali s 1133 58191 1167 58225 6 VGND
port 614 nsew ground input
rlabel viali s 298753 59279 298787 59313 6 VGND
port 614 nsew ground input
rlabel viali s 298661 59279 298695 59313 6 VGND
port 614 nsew ground input
rlabel viali s 1317 59279 1340 59313 6 VGND
port 614 nsew ground input
rlabel viali s 1225 59279 1259 59313 6 VGND
port 614 nsew ground input
rlabel viali s 1133 59279 1167 59313 6 VGND
port 614 nsew ground input
rlabel viali s 298753 60367 298787 60401 6 VGND
port 614 nsew ground input
rlabel viali s 298661 60367 298695 60401 6 VGND
port 614 nsew ground input
rlabel viali s 1317 60367 1340 60401 6 VGND
port 614 nsew ground input
rlabel viali s 1225 60367 1259 60401 6 VGND
port 614 nsew ground input
rlabel viali s 1133 60367 1167 60401 6 VGND
port 614 nsew ground input
rlabel viali s 298753 61455 298787 61489 6 VGND
port 614 nsew ground input
rlabel viali s 298661 61455 298695 61489 6 VGND
port 614 nsew ground input
rlabel viali s 1317 61455 1340 61489 6 VGND
port 614 nsew ground input
rlabel viali s 1225 61455 1259 61489 6 VGND
port 614 nsew ground input
rlabel viali s 1133 61455 1167 61489 6 VGND
port 614 nsew ground input
rlabel viali s 298753 62543 298787 62577 6 VGND
port 614 nsew ground input
rlabel viali s 298661 62543 298695 62577 6 VGND
port 614 nsew ground input
rlabel viali s 1317 62543 1340 62577 6 VGND
port 614 nsew ground input
rlabel viali s 1225 62543 1259 62577 6 VGND
port 614 nsew ground input
rlabel viali s 1133 62543 1167 62577 6 VGND
port 614 nsew ground input
rlabel viali s 298753 63631 298787 63665 6 VGND
port 614 nsew ground input
rlabel viali s 298661 63631 298695 63665 6 VGND
port 614 nsew ground input
rlabel viali s 1317 63631 1340 63665 6 VGND
port 614 nsew ground input
rlabel viali s 1225 63631 1259 63665 6 VGND
port 614 nsew ground input
rlabel viali s 1133 63631 1167 63665 6 VGND
port 614 nsew ground input
rlabel viali s 298753 64719 298787 64753 6 VGND
port 614 nsew ground input
rlabel viali s 298661 64719 298695 64753 6 VGND
port 614 nsew ground input
rlabel viali s 1317 64719 1340 64753 6 VGND
port 614 nsew ground input
rlabel viali s 1225 64719 1259 64753 6 VGND
port 614 nsew ground input
rlabel viali s 1133 64719 1167 64753 6 VGND
port 614 nsew ground input
rlabel viali s 298753 65807 298787 65841 6 VGND
port 614 nsew ground input
rlabel viali s 298661 65807 298695 65841 6 VGND
port 614 nsew ground input
rlabel viali s 1317 65807 1340 65841 6 VGND
port 614 nsew ground input
rlabel viali s 1225 65807 1259 65841 6 VGND
port 614 nsew ground input
rlabel viali s 1133 65807 1167 65841 6 VGND
port 614 nsew ground input
rlabel viali s 298753 66895 298787 66929 6 VGND
port 614 nsew ground input
rlabel viali s 298661 66895 298695 66929 6 VGND
port 614 nsew ground input
rlabel viali s 1317 66895 1340 66929 6 VGND
port 614 nsew ground input
rlabel viali s 1225 66895 1259 66929 6 VGND
port 614 nsew ground input
rlabel viali s 1133 66895 1167 66929 6 VGND
port 614 nsew ground input
rlabel viali s 298753 67983 298787 68017 6 VGND
port 614 nsew ground input
rlabel viali s 298661 67983 298695 68017 6 VGND
port 614 nsew ground input
rlabel viali s 1317 67983 1340 68017 6 VGND
port 614 nsew ground input
rlabel viali s 1225 67983 1259 68017 6 VGND
port 614 nsew ground input
rlabel viali s 1133 67983 1167 68017 6 VGND
port 614 nsew ground input
rlabel viali s 298753 69071 298787 69105 6 VGND
port 614 nsew ground input
rlabel viali s 298661 69071 298695 69105 6 VGND
port 614 nsew ground input
rlabel viali s 1317 69071 1340 69105 6 VGND
port 614 nsew ground input
rlabel viali s 1225 69071 1259 69105 6 VGND
port 614 nsew ground input
rlabel viali s 1133 69071 1167 69105 6 VGND
port 614 nsew ground input
rlabel viali s 298753 70159 298787 70193 6 VGND
port 614 nsew ground input
rlabel viali s 298661 70159 298695 70193 6 VGND
port 614 nsew ground input
rlabel viali s 1317 70159 1340 70193 6 VGND
port 614 nsew ground input
rlabel viali s 1225 70159 1259 70193 6 VGND
port 614 nsew ground input
rlabel viali s 1133 70159 1167 70193 6 VGND
port 614 nsew ground input
rlabel viali s 298753 71247 298787 71281 6 VGND
port 614 nsew ground input
rlabel viali s 298661 71247 298695 71281 6 VGND
port 614 nsew ground input
rlabel viali s 1317 71247 1340 71281 6 VGND
port 614 nsew ground input
rlabel viali s 1225 71247 1259 71281 6 VGND
port 614 nsew ground input
rlabel viali s 1133 71247 1167 71281 6 VGND
port 614 nsew ground input
rlabel viali s 298753 72335 298787 72369 6 VGND
port 614 nsew ground input
rlabel viali s 298661 72335 298695 72369 6 VGND
port 614 nsew ground input
rlabel viali s 1317 72335 1340 72369 6 VGND
port 614 nsew ground input
rlabel viali s 1225 72335 1259 72369 6 VGND
port 614 nsew ground input
rlabel viali s 1133 72335 1167 72369 6 VGND
port 614 nsew ground input
rlabel viali s 298753 73423 298787 73457 6 VGND
port 614 nsew ground input
rlabel viali s 298661 73423 298695 73457 6 VGND
port 614 nsew ground input
rlabel viali s 1317 73423 1340 73457 6 VGND
port 614 nsew ground input
rlabel viali s 1225 73423 1259 73457 6 VGND
port 614 nsew ground input
rlabel viali s 1133 73423 1167 73457 6 VGND
port 614 nsew ground input
rlabel viali s 298753 74511 298787 74545 6 VGND
port 614 nsew ground input
rlabel viali s 298661 74511 298695 74545 6 VGND
port 614 nsew ground input
rlabel viali s 1317 74511 1340 74545 6 VGND
port 614 nsew ground input
rlabel viali s 1225 74511 1259 74545 6 VGND
port 614 nsew ground input
rlabel viali s 1133 74511 1167 74545 6 VGND
port 614 nsew ground input
rlabel viali s 298753 75599 298787 75633 6 VGND
port 614 nsew ground input
rlabel viali s 298661 75599 298695 75633 6 VGND
port 614 nsew ground input
rlabel viali s 1317 75599 1340 75633 6 VGND
port 614 nsew ground input
rlabel viali s 1225 75599 1259 75633 6 VGND
port 614 nsew ground input
rlabel viali s 1133 75599 1167 75633 6 VGND
port 614 nsew ground input
rlabel viali s 298753 76687 298787 76721 6 VGND
port 614 nsew ground input
rlabel viali s 298661 76687 298695 76721 6 VGND
port 614 nsew ground input
rlabel viali s 1317 76687 1340 76721 6 VGND
port 614 nsew ground input
rlabel viali s 1225 76687 1259 76721 6 VGND
port 614 nsew ground input
rlabel viali s 1133 76687 1167 76721 6 VGND
port 614 nsew ground input
rlabel viali s 298753 77775 298787 77809 6 VGND
port 614 nsew ground input
rlabel viali s 298661 77775 298695 77809 6 VGND
port 614 nsew ground input
rlabel viali s 1317 77775 1340 77809 6 VGND
port 614 nsew ground input
rlabel viali s 1225 77775 1259 77809 6 VGND
port 614 nsew ground input
rlabel viali s 1133 77775 1167 77809 6 VGND
port 614 nsew ground input
rlabel viali s 298753 78863 298787 78897 6 VGND
port 614 nsew ground input
rlabel viali s 298661 78863 298695 78897 6 VGND
port 614 nsew ground input
rlabel viali s 1317 78863 1340 78897 6 VGND
port 614 nsew ground input
rlabel viali s 1225 78863 1259 78897 6 VGND
port 614 nsew ground input
rlabel viali s 1133 78863 1167 78897 6 VGND
port 614 nsew ground input
rlabel viali s 298753 79951 298787 79985 6 VGND
port 614 nsew ground input
rlabel viali s 298661 79951 298695 79985 6 VGND
port 614 nsew ground input
rlabel viali s 1317 79951 1340 79985 6 VGND
port 614 nsew ground input
rlabel viali s 1225 79951 1259 79985 6 VGND
port 614 nsew ground input
rlabel viali s 1133 79951 1167 79985 6 VGND
port 614 nsew ground input
rlabel viali s 298753 81039 298787 81073 6 VGND
port 614 nsew ground input
rlabel viali s 298661 81039 298695 81073 6 VGND
port 614 nsew ground input
rlabel viali s 1317 81039 1340 81073 6 VGND
port 614 nsew ground input
rlabel viali s 1225 81039 1259 81073 6 VGND
port 614 nsew ground input
rlabel viali s 1133 81039 1167 81073 6 VGND
port 614 nsew ground input
rlabel viali s 298753 82127 298787 82161 6 VGND
port 614 nsew ground input
rlabel viali s 298661 82127 298695 82161 6 VGND
port 614 nsew ground input
rlabel viali s 1317 82127 1340 82161 6 VGND
port 614 nsew ground input
rlabel viali s 1225 82127 1259 82161 6 VGND
port 614 nsew ground input
rlabel viali s 1133 82127 1167 82161 6 VGND
port 614 nsew ground input
rlabel viali s 298753 83215 298787 83249 6 VGND
port 614 nsew ground input
rlabel viali s 298661 83215 298695 83249 6 VGND
port 614 nsew ground input
rlabel viali s 1317 83215 1340 83249 6 VGND
port 614 nsew ground input
rlabel viali s 1225 83215 1259 83249 6 VGND
port 614 nsew ground input
rlabel viali s 1133 83215 1167 83249 6 VGND
port 614 nsew ground input
rlabel viali s 298753 84303 298787 84337 6 VGND
port 614 nsew ground input
rlabel viali s 298661 84303 298695 84337 6 VGND
port 614 nsew ground input
rlabel viali s 1317 84303 1340 84337 6 VGND
port 614 nsew ground input
rlabel viali s 1225 84303 1259 84337 6 VGND
port 614 nsew ground input
rlabel viali s 1133 84303 1167 84337 6 VGND
port 614 nsew ground input
rlabel viali s 298753 85391 298787 85425 6 VGND
port 614 nsew ground input
rlabel viali s 298661 85391 298695 85425 6 VGND
port 614 nsew ground input
rlabel viali s 1317 85391 1340 85425 6 VGND
port 614 nsew ground input
rlabel viali s 1225 85391 1259 85425 6 VGND
port 614 nsew ground input
rlabel viali s 1133 85391 1167 85425 6 VGND
port 614 nsew ground input
rlabel viali s 298753 86479 298787 86513 6 VGND
port 614 nsew ground input
rlabel viali s 298661 86479 298695 86513 6 VGND
port 614 nsew ground input
rlabel viali s 1317 86479 1340 86513 6 VGND
port 614 nsew ground input
rlabel viali s 1225 86479 1259 86513 6 VGND
port 614 nsew ground input
rlabel viali s 1133 86479 1167 86513 6 VGND
port 614 nsew ground input
rlabel viali s 298753 87567 298787 87601 6 VGND
port 614 nsew ground input
rlabel viali s 298661 87567 298695 87601 6 VGND
port 614 nsew ground input
rlabel viali s 1317 87567 1340 87601 6 VGND
port 614 nsew ground input
rlabel viali s 1225 87567 1259 87601 6 VGND
port 614 nsew ground input
rlabel viali s 1133 87567 1167 87601 6 VGND
port 614 nsew ground input
rlabel viali s 298753 88655 298787 88689 6 VGND
port 614 nsew ground input
rlabel viali s 298661 88655 298695 88689 6 VGND
port 614 nsew ground input
rlabel viali s 1317 88655 1340 88689 6 VGND
port 614 nsew ground input
rlabel viali s 1225 88655 1259 88689 6 VGND
port 614 nsew ground input
rlabel viali s 1133 88655 1167 88689 6 VGND
port 614 nsew ground input
rlabel viali s 298753 89743 298787 89777 6 VGND
port 614 nsew ground input
rlabel viali s 298661 89743 298695 89777 6 VGND
port 614 nsew ground input
rlabel viali s 1317 89743 1340 89777 6 VGND
port 614 nsew ground input
rlabel viali s 1225 89743 1259 89777 6 VGND
port 614 nsew ground input
rlabel viali s 1133 89743 1167 89777 6 VGND
port 614 nsew ground input
rlabel viali s 298753 90831 298787 90865 6 VGND
port 614 nsew ground input
rlabel viali s 298661 90831 298695 90865 6 VGND
port 614 nsew ground input
rlabel viali s 1317 90831 1340 90865 6 VGND
port 614 nsew ground input
rlabel viali s 1225 90831 1259 90865 6 VGND
port 614 nsew ground input
rlabel viali s 1133 90831 1167 90865 6 VGND
port 614 nsew ground input
rlabel viali s 298753 91919 298787 91953 6 VGND
port 614 nsew ground input
rlabel viali s 298661 91919 298695 91953 6 VGND
port 614 nsew ground input
rlabel viali s 1317 91919 1340 91953 6 VGND
port 614 nsew ground input
rlabel viali s 1225 91919 1259 91953 6 VGND
port 614 nsew ground input
rlabel viali s 1133 91919 1167 91953 6 VGND
port 614 nsew ground input
rlabel viali s 298753 93007 298787 93041 6 VGND
port 614 nsew ground input
rlabel viali s 298661 93007 298695 93041 6 VGND
port 614 nsew ground input
rlabel viali s 1317 93007 1340 93041 6 VGND
port 614 nsew ground input
rlabel viali s 1225 93007 1259 93041 6 VGND
port 614 nsew ground input
rlabel viali s 1133 93007 1167 93041 6 VGND
port 614 nsew ground input
rlabel viali s 298753 94095 298787 94129 6 VGND
port 614 nsew ground input
rlabel viali s 298661 94095 298695 94129 6 VGND
port 614 nsew ground input
rlabel viali s 1317 94095 1340 94129 6 VGND
port 614 nsew ground input
rlabel viali s 1225 94095 1259 94129 6 VGND
port 614 nsew ground input
rlabel viali s 1133 94095 1167 94129 6 VGND
port 614 nsew ground input
rlabel viali s 298753 95183 298787 95217 6 VGND
port 614 nsew ground input
rlabel viali s 298661 95183 298695 95217 6 VGND
port 614 nsew ground input
rlabel viali s 1317 95183 1340 95217 6 VGND
port 614 nsew ground input
rlabel viali s 1225 95183 1259 95217 6 VGND
port 614 nsew ground input
rlabel viali s 1133 95183 1167 95217 6 VGND
port 614 nsew ground input
rlabel viali s 298753 96271 298787 96305 6 VGND
port 614 nsew ground input
rlabel viali s 298661 96271 298695 96305 6 VGND
port 614 nsew ground input
rlabel viali s 1317 96271 1340 96305 6 VGND
port 614 nsew ground input
rlabel viali s 1225 96271 1259 96305 6 VGND
port 614 nsew ground input
rlabel viali s 1133 96271 1167 96305 6 VGND
port 614 nsew ground input
rlabel viali s 298753 97359 298787 97393 6 VGND
port 614 nsew ground input
rlabel viali s 298661 97359 298695 97393 6 VGND
port 614 nsew ground input
rlabel viali s 1317 97359 1340 97393 6 VGND
port 614 nsew ground input
rlabel viali s 1225 97359 1259 97393 6 VGND
port 614 nsew ground input
rlabel viali s 1133 97359 1167 97393 6 VGND
port 614 nsew ground input
rlabel viali s 298753 98447 298787 98481 6 VGND
port 614 nsew ground input
rlabel viali s 298661 98447 298695 98481 6 VGND
port 614 nsew ground input
rlabel viali s 1317 98447 1340 98481 6 VGND
port 614 nsew ground input
rlabel viali s 1225 98447 1259 98481 6 VGND
port 614 nsew ground input
rlabel viali s 1133 98447 1167 98481 6 VGND
port 614 nsew ground input
rlabel viali s 298753 99535 298787 99569 6 VGND
port 614 nsew ground input
rlabel viali s 298661 99535 298695 99569 6 VGND
port 614 nsew ground input
rlabel viali s 1317 99535 1340 99569 6 VGND
port 614 nsew ground input
rlabel viali s 1225 99535 1259 99569 6 VGND
port 614 nsew ground input
rlabel viali s 1133 99535 1167 99569 6 VGND
port 614 nsew ground input
rlabel viali s 298753 100623 298787 100657 6 VGND
port 614 nsew ground input
rlabel viali s 298661 100623 298695 100657 6 VGND
port 614 nsew ground input
rlabel viali s 1317 100623 1340 100657 6 VGND
port 614 nsew ground input
rlabel viali s 1225 100623 1259 100657 6 VGND
port 614 nsew ground input
rlabel viali s 1133 100623 1167 100657 6 VGND
port 614 nsew ground input
rlabel viali s 298753 101711 298787 101745 6 VGND
port 614 nsew ground input
rlabel viali s 298661 101711 298695 101745 6 VGND
port 614 nsew ground input
rlabel viali s 1317 101711 1340 101745 6 VGND
port 614 nsew ground input
rlabel viali s 1225 101711 1259 101745 6 VGND
port 614 nsew ground input
rlabel viali s 1133 101711 1167 101745 6 VGND
port 614 nsew ground input
rlabel viali s 298753 102799 298787 102833 6 VGND
port 614 nsew ground input
rlabel viali s 298661 102799 298695 102833 6 VGND
port 614 nsew ground input
rlabel viali s 1317 102799 1340 102833 6 VGND
port 614 nsew ground input
rlabel viali s 1225 102799 1259 102833 6 VGND
port 614 nsew ground input
rlabel viali s 1133 102799 1167 102833 6 VGND
port 614 nsew ground input
rlabel viali s 298753 103887 298787 103921 6 VGND
port 614 nsew ground input
rlabel viali s 298661 103887 298695 103921 6 VGND
port 614 nsew ground input
rlabel viali s 1317 103887 1340 103921 6 VGND
port 614 nsew ground input
rlabel viali s 1225 103887 1259 103921 6 VGND
port 614 nsew ground input
rlabel viali s 1133 103887 1167 103921 6 VGND
port 614 nsew ground input
rlabel viali s 298753 104975 298787 105009 6 VGND
port 614 nsew ground input
rlabel viali s 298661 104975 298695 105009 6 VGND
port 614 nsew ground input
rlabel viali s 1317 104975 1340 105009 6 VGND
port 614 nsew ground input
rlabel viali s 1225 104975 1259 105009 6 VGND
port 614 nsew ground input
rlabel viali s 1133 104975 1167 105009 6 VGND
port 614 nsew ground input
rlabel viali s 298753 106063 298787 106097 6 VGND
port 614 nsew ground input
rlabel viali s 298661 106063 298695 106097 6 VGND
port 614 nsew ground input
rlabel viali s 1317 106063 1340 106097 6 VGND
port 614 nsew ground input
rlabel viali s 1225 106063 1259 106097 6 VGND
port 614 nsew ground input
rlabel viali s 1133 106063 1167 106097 6 VGND
port 614 nsew ground input
rlabel viali s 298753 107151 298787 107185 6 VGND
port 614 nsew ground input
rlabel viali s 298661 107151 298695 107185 6 VGND
port 614 nsew ground input
rlabel viali s 1317 107151 1340 107185 6 VGND
port 614 nsew ground input
rlabel viali s 1225 107151 1259 107185 6 VGND
port 614 nsew ground input
rlabel viali s 1133 107151 1167 107185 6 VGND
port 614 nsew ground input
rlabel viali s 298753 108239 298787 108273 6 VGND
port 614 nsew ground input
rlabel viali s 298661 108239 298695 108273 6 VGND
port 614 nsew ground input
rlabel viali s 1317 108239 1340 108273 6 VGND
port 614 nsew ground input
rlabel viali s 1225 108239 1259 108273 6 VGND
port 614 nsew ground input
rlabel viali s 1133 108239 1167 108273 6 VGND
port 614 nsew ground input
rlabel viali s 298753 109327 298787 109361 6 VGND
port 614 nsew ground input
rlabel viali s 298661 109327 298695 109361 6 VGND
port 614 nsew ground input
rlabel viali s 1317 109327 1340 109361 6 VGND
port 614 nsew ground input
rlabel viali s 1225 109327 1259 109361 6 VGND
port 614 nsew ground input
rlabel viali s 1133 109327 1167 109361 6 VGND
port 614 nsew ground input
rlabel viali s 298753 110415 298787 110449 6 VGND
port 614 nsew ground input
rlabel viali s 298661 110415 298695 110449 6 VGND
port 614 nsew ground input
rlabel viali s 1317 110415 1340 110449 6 VGND
port 614 nsew ground input
rlabel viali s 1225 110415 1259 110449 6 VGND
port 614 nsew ground input
rlabel viali s 1133 110415 1167 110449 6 VGND
port 614 nsew ground input
rlabel viali s 298753 111503 298787 111537 6 VGND
port 614 nsew ground input
rlabel viali s 298661 111503 298695 111537 6 VGND
port 614 nsew ground input
rlabel viali s 1317 111503 1340 111537 6 VGND
port 614 nsew ground input
rlabel viali s 1225 111503 1259 111537 6 VGND
port 614 nsew ground input
rlabel viali s 1133 111503 1167 111537 6 VGND
port 614 nsew ground input
rlabel viali s 298753 112591 298787 112625 6 VGND
port 614 nsew ground input
rlabel viali s 298661 112591 298695 112625 6 VGND
port 614 nsew ground input
rlabel viali s 1317 112591 1340 112625 6 VGND
port 614 nsew ground input
rlabel viali s 1225 112591 1259 112625 6 VGND
port 614 nsew ground input
rlabel viali s 1133 112591 1167 112625 6 VGND
port 614 nsew ground input
rlabel viali s 298753 113679 298787 113713 6 VGND
port 614 nsew ground input
rlabel viali s 298661 113679 298695 113713 6 VGND
port 614 nsew ground input
rlabel viali s 1317 113679 1340 113713 6 VGND
port 614 nsew ground input
rlabel viali s 1225 113679 1259 113713 6 VGND
port 614 nsew ground input
rlabel viali s 1133 113679 1167 113713 6 VGND
port 614 nsew ground input
rlabel viali s 298753 114767 298787 114801 6 VGND
port 614 nsew ground input
rlabel viali s 298661 114767 298695 114801 6 VGND
port 614 nsew ground input
rlabel viali s 1317 114767 1340 114801 6 VGND
port 614 nsew ground input
rlabel viali s 1225 114767 1259 114801 6 VGND
port 614 nsew ground input
rlabel viali s 1133 114767 1167 114801 6 VGND
port 614 nsew ground input
rlabel viali s 298753 115855 298787 115889 6 VGND
port 614 nsew ground input
rlabel viali s 298661 115855 298695 115889 6 VGND
port 614 nsew ground input
rlabel viali s 1317 115855 1340 115889 6 VGND
port 614 nsew ground input
rlabel viali s 1225 115855 1259 115889 6 VGND
port 614 nsew ground input
rlabel viali s 1133 115855 1167 115889 6 VGND
port 614 nsew ground input
rlabel viali s 298753 116943 298787 116977 6 VGND
port 614 nsew ground input
rlabel viali s 298661 116943 298695 116977 6 VGND
port 614 nsew ground input
rlabel viali s 1317 116943 1340 116977 6 VGND
port 614 nsew ground input
rlabel viali s 1225 116943 1259 116977 6 VGND
port 614 nsew ground input
rlabel viali s 1133 116943 1167 116977 6 VGND
port 614 nsew ground input
rlabel viali s 298753 118031 298787 118065 6 VGND
port 614 nsew ground input
rlabel viali s 298661 118031 298695 118065 6 VGND
port 614 nsew ground input
rlabel viali s 1317 118031 1340 118065 6 VGND
port 614 nsew ground input
rlabel viali s 1225 118031 1259 118065 6 VGND
port 614 nsew ground input
rlabel viali s 1133 118031 1167 118065 6 VGND
port 614 nsew ground input
rlabel viali s 298753 119119 298787 119153 6 VGND
port 614 nsew ground input
rlabel viali s 298661 119119 298695 119153 6 VGND
port 614 nsew ground input
rlabel viali s 1317 119119 1340 119153 6 VGND
port 614 nsew ground input
rlabel viali s 1225 119119 1259 119153 6 VGND
port 614 nsew ground input
rlabel viali s 1133 119119 1167 119153 6 VGND
port 614 nsew ground input
rlabel viali s 298753 120207 298787 120241 6 VGND
port 614 nsew ground input
rlabel viali s 298661 120207 298695 120241 6 VGND
port 614 nsew ground input
rlabel viali s 1317 120207 1340 120241 6 VGND
port 614 nsew ground input
rlabel viali s 1225 120207 1259 120241 6 VGND
port 614 nsew ground input
rlabel viali s 1133 120207 1167 120241 6 VGND
port 614 nsew ground input
rlabel viali s 298753 121295 298787 121329 6 VGND
port 614 nsew ground input
rlabel viali s 298661 121295 298695 121329 6 VGND
port 614 nsew ground input
rlabel viali s 1317 121295 1340 121329 6 VGND
port 614 nsew ground input
rlabel viali s 1225 121295 1259 121329 6 VGND
port 614 nsew ground input
rlabel viali s 1133 121295 1167 121329 6 VGND
port 614 nsew ground input
rlabel viali s 298753 122383 298787 122417 6 VGND
port 614 nsew ground input
rlabel viali s 298661 122383 298695 122417 6 VGND
port 614 nsew ground input
rlabel viali s 1317 122383 1340 122417 6 VGND
port 614 nsew ground input
rlabel viali s 1225 122383 1259 122417 6 VGND
port 614 nsew ground input
rlabel viali s 1133 122383 1167 122417 6 VGND
port 614 nsew ground input
rlabel viali s 298753 123471 298787 123505 6 VGND
port 614 nsew ground input
rlabel viali s 298661 123471 298695 123505 6 VGND
port 614 nsew ground input
rlabel viali s 1317 123471 1340 123505 6 VGND
port 614 nsew ground input
rlabel viali s 1225 123471 1259 123505 6 VGND
port 614 nsew ground input
rlabel viali s 1133 123471 1167 123505 6 VGND
port 614 nsew ground input
rlabel viali s 298753 124559 298787 124593 6 VGND
port 614 nsew ground input
rlabel viali s 298661 124559 298695 124593 6 VGND
port 614 nsew ground input
rlabel viali s 1317 124559 1340 124593 6 VGND
port 614 nsew ground input
rlabel viali s 1225 124559 1259 124593 6 VGND
port 614 nsew ground input
rlabel viali s 1133 124559 1167 124593 6 VGND
port 614 nsew ground input
rlabel viali s 298753 125647 298787 125681 6 VGND
port 614 nsew ground input
rlabel viali s 298661 125647 298695 125681 6 VGND
port 614 nsew ground input
rlabel viali s 1317 125647 1340 125681 6 VGND
port 614 nsew ground input
rlabel viali s 1225 125647 1259 125681 6 VGND
port 614 nsew ground input
rlabel viali s 1133 125647 1167 125681 6 VGND
port 614 nsew ground input
rlabel viali s 298753 126735 298787 126769 6 VGND
port 614 nsew ground input
rlabel viali s 298661 126735 298695 126769 6 VGND
port 614 nsew ground input
rlabel viali s 1317 126735 1340 126769 6 VGND
port 614 nsew ground input
rlabel viali s 1225 126735 1259 126769 6 VGND
port 614 nsew ground input
rlabel viali s 1133 126735 1167 126769 6 VGND
port 614 nsew ground input
rlabel viali s 298753 127823 298787 127857 6 VGND
port 614 nsew ground input
rlabel viali s 298661 127823 298695 127857 6 VGND
port 614 nsew ground input
rlabel viali s 1317 127823 1340 127857 6 VGND
port 614 nsew ground input
rlabel viali s 1225 127823 1259 127857 6 VGND
port 614 nsew ground input
rlabel viali s 1133 127823 1167 127857 6 VGND
port 614 nsew ground input
rlabel viali s 298753 128911 298787 128945 6 VGND
port 614 nsew ground input
rlabel viali s 298661 128911 298695 128945 6 VGND
port 614 nsew ground input
rlabel viali s 1317 128911 1340 128945 6 VGND
port 614 nsew ground input
rlabel viali s 1225 128911 1259 128945 6 VGND
port 614 nsew ground input
rlabel viali s 1133 128911 1167 128945 6 VGND
port 614 nsew ground input
rlabel viali s 298753 129999 298787 130033 6 VGND
port 614 nsew ground input
rlabel viali s 298661 129999 298695 130033 6 VGND
port 614 nsew ground input
rlabel viali s 1317 129999 1340 130033 6 VGND
port 614 nsew ground input
rlabel viali s 1225 129999 1259 130033 6 VGND
port 614 nsew ground input
rlabel viali s 1133 129999 1167 130033 6 VGND
port 614 nsew ground input
rlabel viali s 298753 131087 298787 131121 6 VGND
port 614 nsew ground input
rlabel viali s 298661 131087 298695 131121 6 VGND
port 614 nsew ground input
rlabel viali s 1317 131087 1340 131121 6 VGND
port 614 nsew ground input
rlabel viali s 1225 131087 1259 131121 6 VGND
port 614 nsew ground input
rlabel viali s 1133 131087 1167 131121 6 VGND
port 614 nsew ground input
rlabel viali s 298753 132175 298787 132209 6 VGND
port 614 nsew ground input
rlabel viali s 298661 132175 298695 132209 6 VGND
port 614 nsew ground input
rlabel viali s 1317 132175 1340 132209 6 VGND
port 614 nsew ground input
rlabel viali s 1225 132175 1259 132209 6 VGND
port 614 nsew ground input
rlabel viali s 1133 132175 1167 132209 6 VGND
port 614 nsew ground input
rlabel viali s 298753 133263 298787 133297 6 VGND
port 614 nsew ground input
rlabel viali s 298661 133263 298695 133297 6 VGND
port 614 nsew ground input
rlabel viali s 1317 133263 1340 133297 6 VGND
port 614 nsew ground input
rlabel viali s 1225 133263 1259 133297 6 VGND
port 614 nsew ground input
rlabel viali s 1133 133263 1167 133297 6 VGND
port 614 nsew ground input
rlabel viali s 298753 134351 298787 134385 6 VGND
port 614 nsew ground input
rlabel viali s 298661 134351 298695 134385 6 VGND
port 614 nsew ground input
rlabel viali s 1317 134351 1340 134385 6 VGND
port 614 nsew ground input
rlabel viali s 1225 134351 1259 134385 6 VGND
port 614 nsew ground input
rlabel viali s 1133 134351 1167 134385 6 VGND
port 614 nsew ground input
rlabel viali s 298753 135439 298787 135473 6 VGND
port 614 nsew ground input
rlabel viali s 298661 135439 298695 135473 6 VGND
port 614 nsew ground input
rlabel viali s 1317 135439 1340 135473 6 VGND
port 614 nsew ground input
rlabel viali s 1225 135439 1259 135473 6 VGND
port 614 nsew ground input
rlabel viali s 1133 135439 1167 135473 6 VGND
port 614 nsew ground input
rlabel viali s 298753 136527 298787 136561 6 VGND
port 614 nsew ground input
rlabel viali s 298661 136527 298695 136561 6 VGND
port 614 nsew ground input
rlabel viali s 1317 136527 1340 136561 6 VGND
port 614 nsew ground input
rlabel viali s 1225 136527 1259 136561 6 VGND
port 614 nsew ground input
rlabel viali s 1133 136527 1167 136561 6 VGND
port 614 nsew ground input
rlabel viali s 298753 137615 298787 137649 6 VGND
port 614 nsew ground input
rlabel viali s 298661 137615 298695 137649 6 VGND
port 614 nsew ground input
rlabel viali s 1317 137615 1340 137649 6 VGND
port 614 nsew ground input
rlabel viali s 1225 137615 1259 137649 6 VGND
port 614 nsew ground input
rlabel viali s 1133 137615 1167 137649 6 VGND
port 614 nsew ground input
rlabel viali s 298753 138703 298787 138737 6 VGND
port 614 nsew ground input
rlabel viali s 298661 138703 298695 138737 6 VGND
port 614 nsew ground input
rlabel viali s 1317 138703 1340 138737 6 VGND
port 614 nsew ground input
rlabel viali s 1225 138703 1259 138737 6 VGND
port 614 nsew ground input
rlabel viali s 1133 138703 1167 138737 6 VGND
port 614 nsew ground input
rlabel viali s 298753 139791 298787 139825 6 VGND
port 614 nsew ground input
rlabel viali s 298661 139791 298695 139825 6 VGND
port 614 nsew ground input
rlabel viali s 1317 139791 1340 139825 6 VGND
port 614 nsew ground input
rlabel viali s 1225 139791 1259 139825 6 VGND
port 614 nsew ground input
rlabel viali s 1133 139791 1167 139825 6 VGND
port 614 nsew ground input
rlabel viali s 298753 140879 298787 140913 6 VGND
port 614 nsew ground input
rlabel viali s 298661 140879 298695 140913 6 VGND
port 614 nsew ground input
rlabel viali s 1317 140879 1340 140913 6 VGND
port 614 nsew ground input
rlabel viali s 1225 140879 1259 140913 6 VGND
port 614 nsew ground input
rlabel viali s 1133 140879 1167 140913 6 VGND
port 614 nsew ground input
rlabel viali s 298753 141967 298787 142001 6 VGND
port 614 nsew ground input
rlabel viali s 298661 141967 298695 142001 6 VGND
port 614 nsew ground input
rlabel viali s 1317 141967 1340 142001 6 VGND
port 614 nsew ground input
rlabel viali s 1225 141967 1259 142001 6 VGND
port 614 nsew ground input
rlabel viali s 1133 141967 1167 142001 6 VGND
port 614 nsew ground input
rlabel viali s 298753 143055 298787 143089 6 VGND
port 614 nsew ground input
rlabel viali s 298661 143055 298695 143089 6 VGND
port 614 nsew ground input
rlabel viali s 1317 143055 1340 143089 6 VGND
port 614 nsew ground input
rlabel viali s 1225 143055 1259 143089 6 VGND
port 614 nsew ground input
rlabel viali s 1133 143055 1167 143089 6 VGND
port 614 nsew ground input
rlabel viali s 298753 144143 298787 144177 6 VGND
port 614 nsew ground input
rlabel viali s 298661 144143 298695 144177 6 VGND
port 614 nsew ground input
rlabel viali s 1317 144143 1340 144177 6 VGND
port 614 nsew ground input
rlabel viali s 1225 144143 1259 144177 6 VGND
port 614 nsew ground input
rlabel viali s 1133 144143 1167 144177 6 VGND
port 614 nsew ground input
rlabel viali s 298753 145231 298787 145265 6 VGND
port 614 nsew ground input
rlabel viali s 298661 145231 298695 145265 6 VGND
port 614 nsew ground input
rlabel viali s 1317 145231 1340 145265 6 VGND
port 614 nsew ground input
rlabel viali s 1225 145231 1259 145265 6 VGND
port 614 nsew ground input
rlabel viali s 1133 145231 1167 145265 6 VGND
port 614 nsew ground input
rlabel viali s 298753 146319 298787 146353 6 VGND
port 614 nsew ground input
rlabel viali s 298661 146319 298695 146353 6 VGND
port 614 nsew ground input
rlabel viali s 1317 146319 1340 146353 6 VGND
port 614 nsew ground input
rlabel viali s 1225 146319 1259 146353 6 VGND
port 614 nsew ground input
rlabel viali s 1133 146319 1167 146353 6 VGND
port 614 nsew ground input
rlabel viali s 298753 147407 298787 147441 6 VGND
port 614 nsew ground input
rlabel viali s 298661 147407 298695 147441 6 VGND
port 614 nsew ground input
rlabel viali s 1317 147407 1340 147441 6 VGND
port 614 nsew ground input
rlabel viali s 1225 147407 1259 147441 6 VGND
port 614 nsew ground input
rlabel viali s 1133 147407 1167 147441 6 VGND
port 614 nsew ground input
rlabel viali s 298753 148495 298787 148529 6 VGND
port 614 nsew ground input
rlabel viali s 298661 148495 298695 148529 6 VGND
port 614 nsew ground input
rlabel viali s 1317 148495 1340 148529 6 VGND
port 614 nsew ground input
rlabel viali s 1225 148495 1259 148529 6 VGND
port 614 nsew ground input
rlabel viali s 1133 148495 1167 148529 6 VGND
port 614 nsew ground input
rlabel viali s 298753 149583 298787 149617 6 VGND
port 614 nsew ground input
rlabel viali s 298661 149583 298695 149617 6 VGND
port 614 nsew ground input
rlabel viali s 1317 149583 1340 149617 6 VGND
port 614 nsew ground input
rlabel viali s 1225 149583 1259 149617 6 VGND
port 614 nsew ground input
rlabel viali s 1133 149583 1167 149617 6 VGND
port 614 nsew ground input
rlabel viali s 298753 150671 298787 150705 6 VGND
port 614 nsew ground input
rlabel viali s 298661 150671 298695 150705 6 VGND
port 614 nsew ground input
rlabel viali s 1317 150671 1340 150705 6 VGND
port 614 nsew ground input
rlabel viali s 1225 150671 1259 150705 6 VGND
port 614 nsew ground input
rlabel viali s 1133 150671 1167 150705 6 VGND
port 614 nsew ground input
rlabel viali s 298753 151759 298787 151793 6 VGND
port 614 nsew ground input
rlabel viali s 298661 151759 298695 151793 6 VGND
port 614 nsew ground input
rlabel viali s 1317 151759 1340 151793 6 VGND
port 614 nsew ground input
rlabel viali s 1225 151759 1259 151793 6 VGND
port 614 nsew ground input
rlabel viali s 1133 151759 1167 151793 6 VGND
port 614 nsew ground input
rlabel viali s 298753 152847 298787 152881 6 VGND
port 614 nsew ground input
rlabel viali s 298661 152847 298695 152881 6 VGND
port 614 nsew ground input
rlabel viali s 1317 152847 1340 152881 6 VGND
port 614 nsew ground input
rlabel viali s 1225 152847 1259 152881 6 VGND
port 614 nsew ground input
rlabel viali s 1133 152847 1167 152881 6 VGND
port 614 nsew ground input
rlabel viali s 298753 153935 298787 153969 6 VGND
port 614 nsew ground input
rlabel viali s 298661 153935 298695 153969 6 VGND
port 614 nsew ground input
rlabel viali s 1317 153935 1340 153969 6 VGND
port 614 nsew ground input
rlabel viali s 1225 153935 1259 153969 6 VGND
port 614 nsew ground input
rlabel viali s 1133 153935 1167 153969 6 VGND
port 614 nsew ground input
rlabel viali s 298753 155023 298787 155057 6 VGND
port 614 nsew ground input
rlabel viali s 298661 155023 298695 155057 6 VGND
port 614 nsew ground input
rlabel viali s 1317 155023 1340 155057 6 VGND
port 614 nsew ground input
rlabel viali s 1225 155023 1259 155057 6 VGND
port 614 nsew ground input
rlabel viali s 1133 155023 1167 155057 6 VGND
port 614 nsew ground input
rlabel viali s 298753 156111 298787 156145 6 VGND
port 614 nsew ground input
rlabel viali s 298661 156111 298695 156145 6 VGND
port 614 nsew ground input
rlabel viali s 1317 156111 1340 156145 6 VGND
port 614 nsew ground input
rlabel viali s 1225 156111 1259 156145 6 VGND
port 614 nsew ground input
rlabel viali s 1133 156111 1167 156145 6 VGND
port 614 nsew ground input
rlabel viali s 298753 157199 298787 157233 6 VGND
port 614 nsew ground input
rlabel viali s 298661 157199 298695 157233 6 VGND
port 614 nsew ground input
rlabel viali s 1317 157199 1340 157233 6 VGND
port 614 nsew ground input
rlabel viali s 1225 157199 1259 157233 6 VGND
port 614 nsew ground input
rlabel viali s 1133 157199 1167 157233 6 VGND
port 614 nsew ground input
rlabel viali s 298753 158287 298787 158321 6 VGND
port 614 nsew ground input
rlabel viali s 298661 158287 298695 158321 6 VGND
port 614 nsew ground input
rlabel viali s 1317 158287 1340 158321 6 VGND
port 614 nsew ground input
rlabel viali s 1225 158287 1259 158321 6 VGND
port 614 nsew ground input
rlabel viali s 1133 158287 1167 158321 6 VGND
port 614 nsew ground input
rlabel viali s 298753 159375 298787 159409 6 VGND
port 614 nsew ground input
rlabel viali s 298661 159375 298695 159409 6 VGND
port 614 nsew ground input
rlabel viali s 1317 159375 1340 159409 6 VGND
port 614 nsew ground input
rlabel viali s 1225 159375 1259 159409 6 VGND
port 614 nsew ground input
rlabel viali s 1133 159375 1167 159409 6 VGND
port 614 nsew ground input
rlabel viali s 298753 160463 298787 160497 6 VGND
port 614 nsew ground input
rlabel viali s 298661 160463 298695 160497 6 VGND
port 614 nsew ground input
rlabel viali s 1317 160463 1340 160497 6 VGND
port 614 nsew ground input
rlabel viali s 1225 160463 1259 160497 6 VGND
port 614 nsew ground input
rlabel viali s 1133 160463 1167 160497 6 VGND
port 614 nsew ground input
rlabel viali s 298753 161551 298787 161585 6 VGND
port 614 nsew ground input
rlabel viali s 298661 161551 298695 161585 6 VGND
port 614 nsew ground input
rlabel viali s 1317 161551 1340 161585 6 VGND
port 614 nsew ground input
rlabel viali s 1225 161551 1259 161585 6 VGND
port 614 nsew ground input
rlabel viali s 1133 161551 1167 161585 6 VGND
port 614 nsew ground input
rlabel viali s 298753 162639 298787 162673 6 VGND
port 614 nsew ground input
rlabel viali s 298661 162639 298695 162673 6 VGND
port 614 nsew ground input
rlabel viali s 1317 162639 1340 162673 6 VGND
port 614 nsew ground input
rlabel viali s 1225 162639 1259 162673 6 VGND
port 614 nsew ground input
rlabel viali s 1133 162639 1167 162673 6 VGND
port 614 nsew ground input
rlabel viali s 298753 163727 298787 163761 6 VGND
port 614 nsew ground input
rlabel viali s 298661 163727 298695 163761 6 VGND
port 614 nsew ground input
rlabel viali s 1317 163727 1340 163761 6 VGND
port 614 nsew ground input
rlabel viali s 1225 163727 1259 163761 6 VGND
port 614 nsew ground input
rlabel viali s 1133 163727 1167 163761 6 VGND
port 614 nsew ground input
rlabel viali s 298753 164815 298787 164849 6 VGND
port 614 nsew ground input
rlabel viali s 298661 164815 298695 164849 6 VGND
port 614 nsew ground input
rlabel viali s 1317 164815 1340 164849 6 VGND
port 614 nsew ground input
rlabel viali s 1225 164815 1259 164849 6 VGND
port 614 nsew ground input
rlabel viali s 1133 164815 1167 164849 6 VGND
port 614 nsew ground input
rlabel viali s 298753 165903 298787 165937 6 VGND
port 614 nsew ground input
rlabel viali s 298661 165903 298695 165937 6 VGND
port 614 nsew ground input
rlabel viali s 1317 165903 1340 165937 6 VGND
port 614 nsew ground input
rlabel viali s 1225 165903 1259 165937 6 VGND
port 614 nsew ground input
rlabel viali s 1133 165903 1167 165937 6 VGND
port 614 nsew ground input
rlabel viali s 298753 166991 298787 167025 6 VGND
port 614 nsew ground input
rlabel viali s 298661 166991 298695 167025 6 VGND
port 614 nsew ground input
rlabel viali s 1317 166991 1340 167025 6 VGND
port 614 nsew ground input
rlabel viali s 1225 166991 1259 167025 6 VGND
port 614 nsew ground input
rlabel viali s 1133 166991 1167 167025 6 VGND
port 614 nsew ground input
rlabel viali s 298753 168079 298787 168113 6 VGND
port 614 nsew ground input
rlabel viali s 298661 168079 298695 168113 6 VGND
port 614 nsew ground input
rlabel viali s 1317 168079 1340 168113 6 VGND
port 614 nsew ground input
rlabel viali s 1225 168079 1259 168113 6 VGND
port 614 nsew ground input
rlabel viali s 1133 168079 1167 168113 6 VGND
port 614 nsew ground input
rlabel viali s 298753 169167 298787 169201 6 VGND
port 614 nsew ground input
rlabel viali s 298661 169167 298695 169201 6 VGND
port 614 nsew ground input
rlabel viali s 1317 169167 1340 169201 6 VGND
port 614 nsew ground input
rlabel viali s 1225 169167 1259 169201 6 VGND
port 614 nsew ground input
rlabel viali s 1133 169167 1167 169201 6 VGND
port 614 nsew ground input
rlabel viali s 298753 170255 298787 170289 6 VGND
port 614 nsew ground input
rlabel viali s 298661 170255 298695 170289 6 VGND
port 614 nsew ground input
rlabel viali s 1317 170255 1340 170289 6 VGND
port 614 nsew ground input
rlabel viali s 1225 170255 1259 170289 6 VGND
port 614 nsew ground input
rlabel viali s 1133 170255 1167 170289 6 VGND
port 614 nsew ground input
rlabel viali s 298753 171343 298787 171377 6 VGND
port 614 nsew ground input
rlabel viali s 298661 171343 298695 171377 6 VGND
port 614 nsew ground input
rlabel viali s 1317 171343 1340 171377 6 VGND
port 614 nsew ground input
rlabel viali s 1225 171343 1259 171377 6 VGND
port 614 nsew ground input
rlabel viali s 1133 171343 1167 171377 6 VGND
port 614 nsew ground input
rlabel viali s 298753 172431 298787 172465 6 VGND
port 614 nsew ground input
rlabel viali s 298661 172431 298695 172465 6 VGND
port 614 nsew ground input
rlabel viali s 1317 172431 1340 172465 6 VGND
port 614 nsew ground input
rlabel viali s 1225 172431 1259 172465 6 VGND
port 614 nsew ground input
rlabel viali s 1133 172431 1167 172465 6 VGND
port 614 nsew ground input
rlabel viali s 298753 173519 298787 173553 6 VGND
port 614 nsew ground input
rlabel viali s 298661 173519 298695 173553 6 VGND
port 614 nsew ground input
rlabel viali s 1317 173519 1340 173553 6 VGND
port 614 nsew ground input
rlabel viali s 1225 173519 1259 173553 6 VGND
port 614 nsew ground input
rlabel viali s 1133 173519 1167 173553 6 VGND
port 614 nsew ground input
rlabel viali s 298753 174607 298787 174641 6 VGND
port 614 nsew ground input
rlabel viali s 298661 174607 298695 174641 6 VGND
port 614 nsew ground input
rlabel viali s 1317 174607 1340 174641 6 VGND
port 614 nsew ground input
rlabel viali s 1225 174607 1259 174641 6 VGND
port 614 nsew ground input
rlabel viali s 1133 174607 1167 174641 6 VGND
port 614 nsew ground input
rlabel viali s 298753 175695 298787 175729 6 VGND
port 614 nsew ground input
rlabel viali s 298661 175695 298695 175729 6 VGND
port 614 nsew ground input
rlabel viali s 1317 175695 1340 175729 6 VGND
port 614 nsew ground input
rlabel viali s 1225 175695 1259 175729 6 VGND
port 614 nsew ground input
rlabel viali s 1133 175695 1167 175729 6 VGND
port 614 nsew ground input
rlabel viali s 298753 176783 298787 176817 6 VGND
port 614 nsew ground input
rlabel viali s 298661 176783 298695 176817 6 VGND
port 614 nsew ground input
rlabel viali s 1317 176783 1340 176817 6 VGND
port 614 nsew ground input
rlabel viali s 1225 176783 1259 176817 6 VGND
port 614 nsew ground input
rlabel viali s 1133 176783 1167 176817 6 VGND
port 614 nsew ground input
rlabel viali s 298753 177871 298787 177905 6 VGND
port 614 nsew ground input
rlabel viali s 298661 177871 298695 177905 6 VGND
port 614 nsew ground input
rlabel viali s 1317 177871 1340 177905 6 VGND
port 614 nsew ground input
rlabel viali s 1225 177871 1259 177905 6 VGND
port 614 nsew ground input
rlabel viali s 1133 177871 1167 177905 6 VGND
port 614 nsew ground input
rlabel viali s 298753 178959 298787 178993 6 VGND
port 614 nsew ground input
rlabel viali s 298661 178959 298695 178993 6 VGND
port 614 nsew ground input
rlabel viali s 1317 178959 1340 178993 6 VGND
port 614 nsew ground input
rlabel viali s 1225 178959 1259 178993 6 VGND
port 614 nsew ground input
rlabel viali s 1133 178959 1167 178993 6 VGND
port 614 nsew ground input
rlabel viali s 298753 180047 298787 180081 6 VGND
port 614 nsew ground input
rlabel viali s 298661 180047 298695 180081 6 VGND
port 614 nsew ground input
rlabel viali s 1317 180047 1340 180081 6 VGND
port 614 nsew ground input
rlabel viali s 1225 180047 1259 180081 6 VGND
port 614 nsew ground input
rlabel viali s 1133 180047 1167 180081 6 VGND
port 614 nsew ground input
rlabel viali s 298753 181135 298787 181169 6 VGND
port 614 nsew ground input
rlabel viali s 298661 181135 298695 181169 6 VGND
port 614 nsew ground input
rlabel viali s 1317 181135 1340 181169 6 VGND
port 614 nsew ground input
rlabel viali s 1225 181135 1259 181169 6 VGND
port 614 nsew ground input
rlabel viali s 1133 181135 1167 181169 6 VGND
port 614 nsew ground input
rlabel viali s 298753 182223 298787 182257 6 VGND
port 614 nsew ground input
rlabel viali s 298661 182223 298695 182257 6 VGND
port 614 nsew ground input
rlabel viali s 1317 182223 1340 182257 6 VGND
port 614 nsew ground input
rlabel viali s 1225 182223 1259 182257 6 VGND
port 614 nsew ground input
rlabel viali s 1133 182223 1167 182257 6 VGND
port 614 nsew ground input
rlabel viali s 298753 183311 298787 183345 6 VGND
port 614 nsew ground input
rlabel viali s 298661 183311 298695 183345 6 VGND
port 614 nsew ground input
rlabel viali s 1317 183311 1340 183345 6 VGND
port 614 nsew ground input
rlabel viali s 1225 183311 1259 183345 6 VGND
port 614 nsew ground input
rlabel viali s 1133 183311 1167 183345 6 VGND
port 614 nsew ground input
rlabel viali s 298753 184399 298787 184433 6 VGND
port 614 nsew ground input
rlabel viali s 298661 184399 298695 184433 6 VGND
port 614 nsew ground input
rlabel viali s 1317 184399 1340 184433 6 VGND
port 614 nsew ground input
rlabel viali s 1225 184399 1259 184433 6 VGND
port 614 nsew ground input
rlabel viali s 1133 184399 1167 184433 6 VGND
port 614 nsew ground input
rlabel viali s 298753 185487 298787 185521 6 VGND
port 614 nsew ground input
rlabel viali s 298661 185487 298695 185521 6 VGND
port 614 nsew ground input
rlabel viali s 1317 185487 1340 185521 6 VGND
port 614 nsew ground input
rlabel viali s 1225 185487 1259 185521 6 VGND
port 614 nsew ground input
rlabel viali s 1133 185487 1167 185521 6 VGND
port 614 nsew ground input
rlabel viali s 298753 186575 298787 186609 6 VGND
port 614 nsew ground input
rlabel viali s 298661 186575 298695 186609 6 VGND
port 614 nsew ground input
rlabel viali s 1317 186575 1340 186609 6 VGND
port 614 nsew ground input
rlabel viali s 1225 186575 1259 186609 6 VGND
port 614 nsew ground input
rlabel viali s 1133 186575 1167 186609 6 VGND
port 614 nsew ground input
rlabel viali s 298753 187663 298787 187697 6 VGND
port 614 nsew ground input
rlabel viali s 298661 187663 298695 187697 6 VGND
port 614 nsew ground input
rlabel viali s 1317 187663 1340 187697 6 VGND
port 614 nsew ground input
rlabel viali s 1225 187663 1259 187697 6 VGND
port 614 nsew ground input
rlabel viali s 1133 187663 1167 187697 6 VGND
port 614 nsew ground input
rlabel viali s 298753 188751 298787 188785 6 VGND
port 614 nsew ground input
rlabel viali s 298661 188751 298695 188785 6 VGND
port 614 nsew ground input
rlabel viali s 1317 188751 1340 188785 6 VGND
port 614 nsew ground input
rlabel viali s 1225 188751 1259 188785 6 VGND
port 614 nsew ground input
rlabel viali s 1133 188751 1167 188785 6 VGND
port 614 nsew ground input
rlabel viali s 298753 189839 298787 189873 6 VGND
port 614 nsew ground input
rlabel viali s 298661 189839 298695 189873 6 VGND
port 614 nsew ground input
rlabel viali s 1317 189839 1340 189873 6 VGND
port 614 nsew ground input
rlabel viali s 1225 189839 1259 189873 6 VGND
port 614 nsew ground input
rlabel viali s 1133 189839 1167 189873 6 VGND
port 614 nsew ground input
rlabel viali s 298753 190927 298787 190961 6 VGND
port 614 nsew ground input
rlabel viali s 298661 190927 298695 190961 6 VGND
port 614 nsew ground input
rlabel viali s 1317 190927 1340 190961 6 VGND
port 614 nsew ground input
rlabel viali s 1225 190927 1259 190961 6 VGND
port 614 nsew ground input
rlabel viali s 1133 190927 1167 190961 6 VGND
port 614 nsew ground input
rlabel viali s 298753 192015 298787 192049 6 VGND
port 614 nsew ground input
rlabel viali s 298661 192015 298695 192049 6 VGND
port 614 nsew ground input
rlabel viali s 1317 192015 1340 192049 6 VGND
port 614 nsew ground input
rlabel viali s 1225 192015 1259 192049 6 VGND
port 614 nsew ground input
rlabel viali s 1133 192015 1167 192049 6 VGND
port 614 nsew ground input
rlabel viali s 298753 193103 298787 193137 6 VGND
port 614 nsew ground input
rlabel viali s 298661 193103 298695 193137 6 VGND
port 614 nsew ground input
rlabel viali s 1317 193103 1340 193137 6 VGND
port 614 nsew ground input
rlabel viali s 1225 193103 1259 193137 6 VGND
port 614 nsew ground input
rlabel viali s 1133 193103 1167 193137 6 VGND
port 614 nsew ground input
rlabel viali s 298753 194191 298787 194225 6 VGND
port 614 nsew ground input
rlabel viali s 298661 194191 298695 194225 6 VGND
port 614 nsew ground input
rlabel viali s 1317 194191 1340 194225 6 VGND
port 614 nsew ground input
rlabel viali s 1225 194191 1259 194225 6 VGND
port 614 nsew ground input
rlabel viali s 1133 194191 1167 194225 6 VGND
port 614 nsew ground input
rlabel viali s 298753 195279 298787 195313 6 VGND
port 614 nsew ground input
rlabel viali s 298661 195279 298695 195313 6 VGND
port 614 nsew ground input
rlabel viali s 1317 195279 1340 195313 6 VGND
port 614 nsew ground input
rlabel viali s 1225 195279 1259 195313 6 VGND
port 614 nsew ground input
rlabel viali s 1133 195279 1167 195313 6 VGND
port 614 nsew ground input
rlabel viali s 298753 196367 298787 196401 6 VGND
port 614 nsew ground input
rlabel viali s 298661 196367 298695 196401 6 VGND
port 614 nsew ground input
rlabel viali s 1317 196367 1340 196401 6 VGND
port 614 nsew ground input
rlabel viali s 1225 196367 1259 196401 6 VGND
port 614 nsew ground input
rlabel viali s 1133 196367 1167 196401 6 VGND
port 614 nsew ground input
rlabel viali s 298753 197455 298787 197489 6 VGND
port 614 nsew ground input
rlabel viali s 298661 197455 298695 197489 6 VGND
port 614 nsew ground input
rlabel viali s 1317 197455 1340 197489 6 VGND
port 614 nsew ground input
rlabel viali s 1225 197455 1259 197489 6 VGND
port 614 nsew ground input
rlabel viali s 1133 197455 1167 197489 6 VGND
port 614 nsew ground input
rlabel viali s 298753 198543 298787 198577 6 VGND
port 614 nsew ground input
rlabel viali s 298661 198543 298695 198577 6 VGND
port 614 nsew ground input
rlabel viali s 1317 198543 1340 198577 6 VGND
port 614 nsew ground input
rlabel viali s 1225 198543 1259 198577 6 VGND
port 614 nsew ground input
rlabel viali s 1133 198543 1167 198577 6 VGND
port 614 nsew ground input
rlabel viali s 298753 199631 298787 199665 6 VGND
port 614 nsew ground input
rlabel viali s 298661 199631 298695 199665 6 VGND
port 614 nsew ground input
rlabel viali s 1317 199631 1340 199665 6 VGND
port 614 nsew ground input
rlabel viali s 1225 199631 1259 199665 6 VGND
port 614 nsew ground input
rlabel viali s 1133 199631 1167 199665 6 VGND
port 614 nsew ground input
rlabel viali s 298753 200719 298787 200753 6 VGND
port 614 nsew ground input
rlabel viali s 298661 200719 298695 200753 6 VGND
port 614 nsew ground input
rlabel viali s 1317 200719 1340 200753 6 VGND
port 614 nsew ground input
rlabel viali s 1225 200719 1259 200753 6 VGND
port 614 nsew ground input
rlabel viali s 1133 200719 1167 200753 6 VGND
port 614 nsew ground input
rlabel viali s 298753 201807 298787 201841 6 VGND
port 614 nsew ground input
rlabel viali s 298661 201807 298695 201841 6 VGND
port 614 nsew ground input
rlabel viali s 1317 201807 1340 201841 6 VGND
port 614 nsew ground input
rlabel viali s 1225 201807 1259 201841 6 VGND
port 614 nsew ground input
rlabel viali s 1133 201807 1167 201841 6 VGND
port 614 nsew ground input
rlabel viali s 298753 202895 298787 202929 6 VGND
port 614 nsew ground input
rlabel viali s 298661 202895 298695 202929 6 VGND
port 614 nsew ground input
rlabel viali s 1317 202895 1340 202929 6 VGND
port 614 nsew ground input
rlabel viali s 1225 202895 1259 202929 6 VGND
port 614 nsew ground input
rlabel viali s 1133 202895 1167 202929 6 VGND
port 614 nsew ground input
rlabel viali s 298753 203983 298787 204017 6 VGND
port 614 nsew ground input
rlabel viali s 298661 203983 298695 204017 6 VGND
port 614 nsew ground input
rlabel viali s 1317 203983 1340 204017 6 VGND
port 614 nsew ground input
rlabel viali s 1225 203983 1259 204017 6 VGND
port 614 nsew ground input
rlabel viali s 1133 203983 1167 204017 6 VGND
port 614 nsew ground input
rlabel viali s 298753 205071 298787 205105 6 VGND
port 614 nsew ground input
rlabel viali s 298661 205071 298695 205105 6 VGND
port 614 nsew ground input
rlabel viali s 1317 205071 1340 205105 6 VGND
port 614 nsew ground input
rlabel viali s 1225 205071 1259 205105 6 VGND
port 614 nsew ground input
rlabel viali s 1133 205071 1167 205105 6 VGND
port 614 nsew ground input
rlabel viali s 298753 206159 298787 206193 6 VGND
port 614 nsew ground input
rlabel viali s 298661 206159 298695 206193 6 VGND
port 614 nsew ground input
rlabel viali s 1317 206159 1340 206193 6 VGND
port 614 nsew ground input
rlabel viali s 1225 206159 1259 206193 6 VGND
port 614 nsew ground input
rlabel viali s 1133 206159 1167 206193 6 VGND
port 614 nsew ground input
rlabel viali s 298753 207247 298787 207281 6 VGND
port 614 nsew ground input
rlabel viali s 298661 207247 298695 207281 6 VGND
port 614 nsew ground input
rlabel viali s 1317 207247 1340 207281 6 VGND
port 614 nsew ground input
rlabel viali s 1225 207247 1259 207281 6 VGND
port 614 nsew ground input
rlabel viali s 1133 207247 1167 207281 6 VGND
port 614 nsew ground input
rlabel viali s 298753 208335 298787 208369 6 VGND
port 614 nsew ground input
rlabel viali s 298661 208335 298695 208369 6 VGND
port 614 nsew ground input
rlabel viali s 1317 208335 1340 208369 6 VGND
port 614 nsew ground input
rlabel viali s 1225 208335 1259 208369 6 VGND
port 614 nsew ground input
rlabel viali s 1133 208335 1167 208369 6 VGND
port 614 nsew ground input
rlabel viali s 298753 209423 298787 209457 6 VGND
port 614 nsew ground input
rlabel viali s 298661 209423 298695 209457 6 VGND
port 614 nsew ground input
rlabel viali s 1317 209423 1340 209457 6 VGND
port 614 nsew ground input
rlabel viali s 1225 209423 1259 209457 6 VGND
port 614 nsew ground input
rlabel viali s 1133 209423 1167 209457 6 VGND
port 614 nsew ground input
rlabel viali s 298753 210511 298787 210545 6 VGND
port 614 nsew ground input
rlabel viali s 298661 210511 298695 210545 6 VGND
port 614 nsew ground input
rlabel viali s 1317 210511 1340 210545 6 VGND
port 614 nsew ground input
rlabel viali s 1225 210511 1259 210545 6 VGND
port 614 nsew ground input
rlabel viali s 1133 210511 1167 210545 6 VGND
port 614 nsew ground input
rlabel viali s 298753 211599 298787 211633 6 VGND
port 614 nsew ground input
rlabel viali s 298661 211599 298695 211633 6 VGND
port 614 nsew ground input
rlabel viali s 1317 211599 1340 211633 6 VGND
port 614 nsew ground input
rlabel viali s 1225 211599 1259 211633 6 VGND
port 614 nsew ground input
rlabel viali s 1133 211599 1167 211633 6 VGND
port 614 nsew ground input
rlabel viali s 298753 212687 298787 212721 6 VGND
port 614 nsew ground input
rlabel viali s 298661 212687 298695 212721 6 VGND
port 614 nsew ground input
rlabel viali s 1317 212687 1340 212721 6 VGND
port 614 nsew ground input
rlabel viali s 1225 212687 1259 212721 6 VGND
port 614 nsew ground input
rlabel viali s 1133 212687 1167 212721 6 VGND
port 614 nsew ground input
rlabel viali s 298753 213775 298787 213809 6 VGND
port 614 nsew ground input
rlabel viali s 298661 213775 298695 213809 6 VGND
port 614 nsew ground input
rlabel viali s 1317 213775 1340 213809 6 VGND
port 614 nsew ground input
rlabel viali s 1225 213775 1259 213809 6 VGND
port 614 nsew ground input
rlabel viali s 1133 213775 1167 213809 6 VGND
port 614 nsew ground input
rlabel viali s 298753 214863 298787 214897 6 VGND
port 614 nsew ground input
rlabel viali s 298661 214863 298695 214897 6 VGND
port 614 nsew ground input
rlabel viali s 1317 214863 1340 214897 6 VGND
port 614 nsew ground input
rlabel viali s 1225 214863 1259 214897 6 VGND
port 614 nsew ground input
rlabel viali s 1133 214863 1167 214897 6 VGND
port 614 nsew ground input
rlabel viali s 298753 215951 298787 215985 6 VGND
port 614 nsew ground input
rlabel viali s 298661 215951 298695 215985 6 VGND
port 614 nsew ground input
rlabel viali s 1317 215951 1340 215985 6 VGND
port 614 nsew ground input
rlabel viali s 1225 215951 1259 215985 6 VGND
port 614 nsew ground input
rlabel viali s 1133 215951 1167 215985 6 VGND
port 614 nsew ground input
rlabel viali s 298753 217039 298787 217073 6 VGND
port 614 nsew ground input
rlabel viali s 298661 217039 298695 217073 6 VGND
port 614 nsew ground input
rlabel viali s 1317 217039 1340 217073 6 VGND
port 614 nsew ground input
rlabel viali s 1225 217039 1259 217073 6 VGND
port 614 nsew ground input
rlabel viali s 1133 217039 1167 217073 6 VGND
port 614 nsew ground input
rlabel viali s 298753 218127 298787 218161 6 VGND
port 614 nsew ground input
rlabel viali s 298661 218127 298695 218161 6 VGND
port 614 nsew ground input
rlabel viali s 1317 218127 1340 218161 6 VGND
port 614 nsew ground input
rlabel viali s 1225 218127 1259 218161 6 VGND
port 614 nsew ground input
rlabel viali s 1133 218127 1167 218161 6 VGND
port 614 nsew ground input
rlabel viali s 298753 219215 298787 219249 6 VGND
port 614 nsew ground input
rlabel viali s 298661 219215 298695 219249 6 VGND
port 614 nsew ground input
rlabel viali s 1317 219215 1340 219249 6 VGND
port 614 nsew ground input
rlabel viali s 1225 219215 1259 219249 6 VGND
port 614 nsew ground input
rlabel viali s 1133 219215 1167 219249 6 VGND
port 614 nsew ground input
rlabel viali s 298753 220303 298787 220337 6 VGND
port 614 nsew ground input
rlabel viali s 298661 220303 298695 220337 6 VGND
port 614 nsew ground input
rlabel viali s 1317 220303 1340 220337 6 VGND
port 614 nsew ground input
rlabel viali s 1225 220303 1259 220337 6 VGND
port 614 nsew ground input
rlabel viali s 1133 220303 1167 220337 6 VGND
port 614 nsew ground input
rlabel viali s 298753 221391 298787 221425 6 VGND
port 614 nsew ground input
rlabel viali s 298661 221391 298695 221425 6 VGND
port 614 nsew ground input
rlabel viali s 1317 221391 1340 221425 6 VGND
port 614 nsew ground input
rlabel viali s 1225 221391 1259 221425 6 VGND
port 614 nsew ground input
rlabel viali s 1133 221391 1167 221425 6 VGND
port 614 nsew ground input
rlabel viali s 298753 222479 298787 222513 6 VGND
port 614 nsew ground input
rlabel viali s 298661 222479 298695 222513 6 VGND
port 614 nsew ground input
rlabel viali s 1317 222479 1340 222513 6 VGND
port 614 nsew ground input
rlabel viali s 1225 222479 1259 222513 6 VGND
port 614 nsew ground input
rlabel viali s 1133 222479 1167 222513 6 VGND
port 614 nsew ground input
rlabel viali s 298753 223567 298787 223601 6 VGND
port 614 nsew ground input
rlabel viali s 298661 223567 298695 223601 6 VGND
port 614 nsew ground input
rlabel viali s 1317 223567 1340 223601 6 VGND
port 614 nsew ground input
rlabel viali s 1225 223567 1259 223601 6 VGND
port 614 nsew ground input
rlabel viali s 1133 223567 1167 223601 6 VGND
port 614 nsew ground input
rlabel viali s 298753 224655 298787 224689 6 VGND
port 614 nsew ground input
rlabel viali s 298661 224655 298695 224689 6 VGND
port 614 nsew ground input
rlabel viali s 1317 224655 1340 224689 6 VGND
port 614 nsew ground input
rlabel viali s 1225 224655 1259 224689 6 VGND
port 614 nsew ground input
rlabel viali s 1133 224655 1167 224689 6 VGND
port 614 nsew ground input
rlabel viali s 298753 225743 298787 225777 6 VGND
port 614 nsew ground input
rlabel viali s 298661 225743 298695 225777 6 VGND
port 614 nsew ground input
rlabel viali s 1317 225743 1340 225777 6 VGND
port 614 nsew ground input
rlabel viali s 1225 225743 1259 225777 6 VGND
port 614 nsew ground input
rlabel viali s 1133 225743 1167 225777 6 VGND
port 614 nsew ground input
rlabel viali s 298753 226831 298787 226865 6 VGND
port 614 nsew ground input
rlabel viali s 298661 226831 298695 226865 6 VGND
port 614 nsew ground input
rlabel viali s 1317 226831 1340 226865 6 VGND
port 614 nsew ground input
rlabel viali s 1225 226831 1259 226865 6 VGND
port 614 nsew ground input
rlabel viali s 1133 226831 1167 226865 6 VGND
port 614 nsew ground input
rlabel viali s 298753 227919 298787 227953 6 VGND
port 614 nsew ground input
rlabel viali s 298661 227919 298695 227953 6 VGND
port 614 nsew ground input
rlabel viali s 1317 227919 1340 227953 6 VGND
port 614 nsew ground input
rlabel viali s 1225 227919 1259 227953 6 VGND
port 614 nsew ground input
rlabel viali s 1133 227919 1167 227953 6 VGND
port 614 nsew ground input
rlabel viali s 298753 229007 298787 229041 6 VGND
port 614 nsew ground input
rlabel viali s 298661 229007 298695 229041 6 VGND
port 614 nsew ground input
rlabel viali s 1317 229007 1340 229041 6 VGND
port 614 nsew ground input
rlabel viali s 1225 229007 1259 229041 6 VGND
port 614 nsew ground input
rlabel viali s 1133 229007 1167 229041 6 VGND
port 614 nsew ground input
rlabel viali s 298753 230095 298787 230129 6 VGND
port 614 nsew ground input
rlabel viali s 298661 230095 298695 230129 6 VGND
port 614 nsew ground input
rlabel viali s 1317 230095 1340 230129 6 VGND
port 614 nsew ground input
rlabel viali s 1225 230095 1259 230129 6 VGND
port 614 nsew ground input
rlabel viali s 1133 230095 1167 230129 6 VGND
port 614 nsew ground input
rlabel viali s 298753 231183 298787 231217 6 VGND
port 614 nsew ground input
rlabel viali s 298661 231183 298695 231217 6 VGND
port 614 nsew ground input
rlabel viali s 1317 231183 1340 231217 6 VGND
port 614 nsew ground input
rlabel viali s 1225 231183 1259 231217 6 VGND
port 614 nsew ground input
rlabel viali s 1133 231183 1167 231217 6 VGND
port 614 nsew ground input
rlabel viali s 298753 232271 298787 232305 6 VGND
port 614 nsew ground input
rlabel viali s 298661 232271 298695 232305 6 VGND
port 614 nsew ground input
rlabel viali s 1317 232271 1340 232305 6 VGND
port 614 nsew ground input
rlabel viali s 1225 232271 1259 232305 6 VGND
port 614 nsew ground input
rlabel viali s 1133 232271 1167 232305 6 VGND
port 614 nsew ground input
rlabel viali s 298753 233359 298787 233393 6 VGND
port 614 nsew ground input
rlabel viali s 298661 233359 298695 233393 6 VGND
port 614 nsew ground input
rlabel viali s 1317 233359 1340 233393 6 VGND
port 614 nsew ground input
rlabel viali s 1225 233359 1259 233393 6 VGND
port 614 nsew ground input
rlabel viali s 1133 233359 1167 233393 6 VGND
port 614 nsew ground input
rlabel viali s 298753 234447 298787 234481 6 VGND
port 614 nsew ground input
rlabel viali s 298661 234447 298695 234481 6 VGND
port 614 nsew ground input
rlabel viali s 1317 234447 1340 234481 6 VGND
port 614 nsew ground input
rlabel viali s 1225 234447 1259 234481 6 VGND
port 614 nsew ground input
rlabel viali s 1133 234447 1167 234481 6 VGND
port 614 nsew ground input
rlabel viali s 298753 235535 298787 235569 6 VGND
port 614 nsew ground input
rlabel viali s 298661 235535 298695 235569 6 VGND
port 614 nsew ground input
rlabel viali s 1317 235535 1340 235569 6 VGND
port 614 nsew ground input
rlabel viali s 1225 235535 1259 235569 6 VGND
port 614 nsew ground input
rlabel viali s 1133 235535 1167 235569 6 VGND
port 614 nsew ground input
rlabel viali s 298753 236623 298787 236657 6 VGND
port 614 nsew ground input
rlabel viali s 298661 236623 298695 236657 6 VGND
port 614 nsew ground input
rlabel viali s 1317 236623 1340 236657 6 VGND
port 614 nsew ground input
rlabel viali s 1225 236623 1259 236657 6 VGND
port 614 nsew ground input
rlabel viali s 1133 236623 1167 236657 6 VGND
port 614 nsew ground input
rlabel viali s 298753 237711 298787 237745 6 VGND
port 614 nsew ground input
rlabel viali s 298661 237711 298695 237745 6 VGND
port 614 nsew ground input
rlabel viali s 1317 237711 1340 237745 6 VGND
port 614 nsew ground input
rlabel viali s 1225 237711 1259 237745 6 VGND
port 614 nsew ground input
rlabel viali s 1133 237711 1167 237745 6 VGND
port 614 nsew ground input
rlabel viali s 298753 238799 298787 238833 6 VGND
port 614 nsew ground input
rlabel viali s 298661 238799 298695 238833 6 VGND
port 614 nsew ground input
rlabel viali s 1317 238799 1340 238833 6 VGND
port 614 nsew ground input
rlabel viali s 1225 238799 1259 238833 6 VGND
port 614 nsew ground input
rlabel viali s 1133 238799 1167 238833 6 VGND
port 614 nsew ground input
rlabel viali s 298753 239887 298787 239921 6 VGND
port 614 nsew ground input
rlabel viali s 298661 239887 298695 239921 6 VGND
port 614 nsew ground input
rlabel viali s 1317 239887 1340 239921 6 VGND
port 614 nsew ground input
rlabel viali s 1225 239887 1259 239921 6 VGND
port 614 nsew ground input
rlabel viali s 1133 239887 1167 239921 6 VGND
port 614 nsew ground input
rlabel viali s 298753 240975 298787 241009 6 VGND
port 614 nsew ground input
rlabel viali s 298661 240975 298695 241009 6 VGND
port 614 nsew ground input
rlabel viali s 1317 240975 1340 241009 6 VGND
port 614 nsew ground input
rlabel viali s 1225 240975 1259 241009 6 VGND
port 614 nsew ground input
rlabel viali s 1133 240975 1167 241009 6 VGND
port 614 nsew ground input
rlabel viali s 298753 242063 298787 242097 6 VGND
port 614 nsew ground input
rlabel viali s 298661 242063 298695 242097 6 VGND
port 614 nsew ground input
rlabel viali s 1317 242063 1340 242097 6 VGND
port 614 nsew ground input
rlabel viali s 1225 242063 1259 242097 6 VGND
port 614 nsew ground input
rlabel viali s 1133 242063 1167 242097 6 VGND
port 614 nsew ground input
rlabel viali s 298753 243151 298787 243185 6 VGND
port 614 nsew ground input
rlabel viali s 298661 243151 298695 243185 6 VGND
port 614 nsew ground input
rlabel viali s 1317 243151 1340 243185 6 VGND
port 614 nsew ground input
rlabel viali s 1225 243151 1259 243185 6 VGND
port 614 nsew ground input
rlabel viali s 1133 243151 1167 243185 6 VGND
port 614 nsew ground input
rlabel viali s 298753 244239 298787 244273 6 VGND
port 614 nsew ground input
rlabel viali s 298661 244239 298695 244273 6 VGND
port 614 nsew ground input
rlabel viali s 1317 244239 1340 244273 6 VGND
port 614 nsew ground input
rlabel viali s 1225 244239 1259 244273 6 VGND
port 614 nsew ground input
rlabel viali s 1133 244239 1167 244273 6 VGND
port 614 nsew ground input
rlabel viali s 298753 245327 298787 245361 6 VGND
port 614 nsew ground input
rlabel viali s 298661 245327 298695 245361 6 VGND
port 614 nsew ground input
rlabel viali s 1317 245327 1340 245361 6 VGND
port 614 nsew ground input
rlabel viali s 1225 245327 1259 245361 6 VGND
port 614 nsew ground input
rlabel viali s 1133 245327 1167 245361 6 VGND
port 614 nsew ground input
rlabel viali s 298753 246415 298787 246449 6 VGND
port 614 nsew ground input
rlabel viali s 298661 246415 298695 246449 6 VGND
port 614 nsew ground input
rlabel viali s 1317 246415 1340 246449 6 VGND
port 614 nsew ground input
rlabel viali s 1225 246415 1259 246449 6 VGND
port 614 nsew ground input
rlabel viali s 1133 246415 1167 246449 6 VGND
port 614 nsew ground input
rlabel viali s 298753 247503 298787 247537 6 VGND
port 614 nsew ground input
rlabel viali s 298661 247503 298695 247537 6 VGND
port 614 nsew ground input
rlabel viali s 1317 247503 1340 247537 6 VGND
port 614 nsew ground input
rlabel viali s 1225 247503 1259 247537 6 VGND
port 614 nsew ground input
rlabel viali s 1133 247503 1167 247537 6 VGND
port 614 nsew ground input
rlabel viali s 298753 248591 298787 248625 6 VGND
port 614 nsew ground input
rlabel viali s 298661 248591 298695 248625 6 VGND
port 614 nsew ground input
rlabel viali s 1317 248591 1340 248625 6 VGND
port 614 nsew ground input
rlabel viali s 1225 248591 1259 248625 6 VGND
port 614 nsew ground input
rlabel viali s 1133 248591 1167 248625 6 VGND
port 614 nsew ground input
rlabel viali s 298753 249679 298787 249713 6 VGND
port 614 nsew ground input
rlabel viali s 298661 249679 298695 249713 6 VGND
port 614 nsew ground input
rlabel viali s 1317 249679 1340 249713 6 VGND
port 614 nsew ground input
rlabel viali s 1225 249679 1259 249713 6 VGND
port 614 nsew ground input
rlabel viali s 1133 249679 1167 249713 6 VGND
port 614 nsew ground input
rlabel viali s 298753 250767 298787 250801 6 VGND
port 614 nsew ground input
rlabel viali s 298661 250767 298695 250801 6 VGND
port 614 nsew ground input
rlabel viali s 1317 250767 1340 250801 6 VGND
port 614 nsew ground input
rlabel viali s 1225 250767 1259 250801 6 VGND
port 614 nsew ground input
rlabel viali s 1133 250767 1167 250801 6 VGND
port 614 nsew ground input
rlabel viali s 298753 251855 298787 251889 6 VGND
port 614 nsew ground input
rlabel viali s 298661 251855 298695 251889 6 VGND
port 614 nsew ground input
rlabel viali s 1317 251855 1340 251889 6 VGND
port 614 nsew ground input
rlabel viali s 1225 251855 1259 251889 6 VGND
port 614 nsew ground input
rlabel viali s 1133 251855 1167 251889 6 VGND
port 614 nsew ground input
rlabel viali s 298753 252943 298787 252977 6 VGND
port 614 nsew ground input
rlabel viali s 298661 252943 298695 252977 6 VGND
port 614 nsew ground input
rlabel viali s 1317 252943 1340 252977 6 VGND
port 614 nsew ground input
rlabel viali s 1225 252943 1259 252977 6 VGND
port 614 nsew ground input
rlabel viali s 1133 252943 1167 252977 6 VGND
port 614 nsew ground input
rlabel viali s 298753 254031 298787 254065 6 VGND
port 614 nsew ground input
rlabel viali s 298661 254031 298695 254065 6 VGND
port 614 nsew ground input
rlabel viali s 1317 254031 1340 254065 6 VGND
port 614 nsew ground input
rlabel viali s 1225 254031 1259 254065 6 VGND
port 614 nsew ground input
rlabel viali s 1133 254031 1167 254065 6 VGND
port 614 nsew ground input
rlabel viali s 298753 255119 298787 255153 6 VGND
port 614 nsew ground input
rlabel viali s 298661 255119 298695 255153 6 VGND
port 614 nsew ground input
rlabel viali s 1317 255119 1340 255153 6 VGND
port 614 nsew ground input
rlabel viali s 1225 255119 1259 255153 6 VGND
port 614 nsew ground input
rlabel viali s 1133 255119 1167 255153 6 VGND
port 614 nsew ground input
rlabel viali s 298753 256207 298787 256241 6 VGND
port 614 nsew ground input
rlabel viali s 298661 256207 298695 256241 6 VGND
port 614 nsew ground input
rlabel viali s 1317 256207 1340 256241 6 VGND
port 614 nsew ground input
rlabel viali s 1225 256207 1259 256241 6 VGND
port 614 nsew ground input
rlabel viali s 1133 256207 1167 256241 6 VGND
port 614 nsew ground input
rlabel viali s 298753 257295 298787 257329 6 VGND
port 614 nsew ground input
rlabel viali s 298661 257295 298695 257329 6 VGND
port 614 nsew ground input
rlabel viali s 1317 257295 1340 257329 6 VGND
port 614 nsew ground input
rlabel viali s 1225 257295 1259 257329 6 VGND
port 614 nsew ground input
rlabel viali s 1133 257295 1167 257329 6 VGND
port 614 nsew ground input
rlabel viali s 298753 258383 298787 258417 6 VGND
port 614 nsew ground input
rlabel viali s 298661 258383 298695 258417 6 VGND
port 614 nsew ground input
rlabel viali s 1317 258383 1340 258417 6 VGND
port 614 nsew ground input
rlabel viali s 1225 258383 1259 258417 6 VGND
port 614 nsew ground input
rlabel viali s 1133 258383 1167 258417 6 VGND
port 614 nsew ground input
rlabel viali s 298753 259471 298787 259505 6 VGND
port 614 nsew ground input
rlabel viali s 298661 259471 298695 259505 6 VGND
port 614 nsew ground input
rlabel viali s 1317 259471 1340 259505 6 VGND
port 614 nsew ground input
rlabel viali s 1225 259471 1259 259505 6 VGND
port 614 nsew ground input
rlabel viali s 1133 259471 1167 259505 6 VGND
port 614 nsew ground input
rlabel viali s 298753 260559 298787 260593 6 VGND
port 614 nsew ground input
rlabel viali s 298661 260559 298695 260593 6 VGND
port 614 nsew ground input
rlabel viali s 1317 260559 1340 260593 6 VGND
port 614 nsew ground input
rlabel viali s 1225 260559 1259 260593 6 VGND
port 614 nsew ground input
rlabel viali s 1133 260559 1167 260593 6 VGND
port 614 nsew ground input
rlabel viali s 298753 261647 298787 261681 6 VGND
port 614 nsew ground input
rlabel viali s 298661 261647 298695 261681 6 VGND
port 614 nsew ground input
rlabel viali s 1317 261647 1340 261681 6 VGND
port 614 nsew ground input
rlabel viali s 1225 261647 1259 261681 6 VGND
port 614 nsew ground input
rlabel viali s 1133 261647 1167 261681 6 VGND
port 614 nsew ground input
rlabel viali s 298753 262735 298787 262769 6 VGND
port 614 nsew ground input
rlabel viali s 298661 262735 298695 262769 6 VGND
port 614 nsew ground input
rlabel viali s 1317 262735 1340 262769 6 VGND
port 614 nsew ground input
rlabel viali s 1225 262735 1259 262769 6 VGND
port 614 nsew ground input
rlabel viali s 1133 262735 1167 262769 6 VGND
port 614 nsew ground input
rlabel viali s 298753 263823 298787 263857 6 VGND
port 614 nsew ground input
rlabel viali s 298661 263823 298695 263857 6 VGND
port 614 nsew ground input
rlabel viali s 1317 263823 1340 263857 6 VGND
port 614 nsew ground input
rlabel viali s 1225 263823 1259 263857 6 VGND
port 614 nsew ground input
rlabel viali s 1133 263823 1167 263857 6 VGND
port 614 nsew ground input
rlabel viali s 298753 264911 298787 264945 6 VGND
port 614 nsew ground input
rlabel viali s 298661 264911 298695 264945 6 VGND
port 614 nsew ground input
rlabel viali s 1317 264911 1340 264945 6 VGND
port 614 nsew ground input
rlabel viali s 1225 264911 1259 264945 6 VGND
port 614 nsew ground input
rlabel viali s 1133 264911 1167 264945 6 VGND
port 614 nsew ground input
rlabel viali s 298753 265999 298787 266033 6 VGND
port 614 nsew ground input
rlabel viali s 298661 265999 298695 266033 6 VGND
port 614 nsew ground input
rlabel viali s 1317 265999 1340 266033 6 VGND
port 614 nsew ground input
rlabel viali s 1225 265999 1259 266033 6 VGND
port 614 nsew ground input
rlabel viali s 1133 265999 1167 266033 6 VGND
port 614 nsew ground input
rlabel viali s 298753 267087 298787 267121 6 VGND
port 614 nsew ground input
rlabel viali s 298661 267087 298695 267121 6 VGND
port 614 nsew ground input
rlabel viali s 1317 267087 1340 267121 6 VGND
port 614 nsew ground input
rlabel viali s 1225 267087 1259 267121 6 VGND
port 614 nsew ground input
rlabel viali s 1133 267087 1167 267121 6 VGND
port 614 nsew ground input
rlabel viali s 298753 268175 298787 268209 6 VGND
port 614 nsew ground input
rlabel viali s 298661 268175 298695 268209 6 VGND
port 614 nsew ground input
rlabel viali s 1317 268175 1340 268209 6 VGND
port 614 nsew ground input
rlabel viali s 1225 268175 1259 268209 6 VGND
port 614 nsew ground input
rlabel viali s 1133 268175 1167 268209 6 VGND
port 614 nsew ground input
rlabel viali s 298753 269263 298787 269297 6 VGND
port 614 nsew ground input
rlabel viali s 298661 269263 298695 269297 6 VGND
port 614 nsew ground input
rlabel viali s 1317 269263 1340 269297 6 VGND
port 614 nsew ground input
rlabel viali s 1225 269263 1259 269297 6 VGND
port 614 nsew ground input
rlabel viali s 1133 269263 1167 269297 6 VGND
port 614 nsew ground input
rlabel viali s 298753 270351 298787 270385 6 VGND
port 614 nsew ground input
rlabel viali s 298661 270351 298695 270385 6 VGND
port 614 nsew ground input
rlabel viali s 1317 270351 1340 270385 6 VGND
port 614 nsew ground input
rlabel viali s 1225 270351 1259 270385 6 VGND
port 614 nsew ground input
rlabel viali s 1133 270351 1167 270385 6 VGND
port 614 nsew ground input
rlabel viali s 298753 271439 298787 271473 6 VGND
port 614 nsew ground input
rlabel viali s 298661 271439 298695 271473 6 VGND
port 614 nsew ground input
rlabel viali s 1317 271439 1340 271473 6 VGND
port 614 nsew ground input
rlabel viali s 1225 271439 1259 271473 6 VGND
port 614 nsew ground input
rlabel viali s 1133 271439 1167 271473 6 VGND
port 614 nsew ground input
rlabel viali s 298753 272527 298787 272561 6 VGND
port 614 nsew ground input
rlabel viali s 298661 272527 298695 272561 6 VGND
port 614 nsew ground input
rlabel viali s 1317 272527 1340 272561 6 VGND
port 614 nsew ground input
rlabel viali s 1225 272527 1259 272561 6 VGND
port 614 nsew ground input
rlabel viali s 1133 272527 1167 272561 6 VGND
port 614 nsew ground input
rlabel viali s 298753 273615 298787 273649 6 VGND
port 614 nsew ground input
rlabel viali s 298661 273615 298695 273649 6 VGND
port 614 nsew ground input
rlabel viali s 1317 273615 1340 273649 6 VGND
port 614 nsew ground input
rlabel viali s 1225 273615 1259 273649 6 VGND
port 614 nsew ground input
rlabel viali s 1133 273615 1167 273649 6 VGND
port 614 nsew ground input
rlabel viali s 298753 274703 298787 274737 6 VGND
port 614 nsew ground input
rlabel viali s 298661 274703 298695 274737 6 VGND
port 614 nsew ground input
rlabel viali s 1317 274703 1340 274737 6 VGND
port 614 nsew ground input
rlabel viali s 1225 274703 1259 274737 6 VGND
port 614 nsew ground input
rlabel viali s 1133 274703 1167 274737 6 VGND
port 614 nsew ground input
rlabel viali s 298753 275791 298787 275825 6 VGND
port 614 nsew ground input
rlabel viali s 298661 275791 298695 275825 6 VGND
port 614 nsew ground input
rlabel viali s 1317 275791 1340 275825 6 VGND
port 614 nsew ground input
rlabel viali s 1225 275791 1259 275825 6 VGND
port 614 nsew ground input
rlabel viali s 1133 275791 1167 275825 6 VGND
port 614 nsew ground input
rlabel viali s 298753 276879 298787 276913 6 VGND
port 614 nsew ground input
rlabel viali s 298661 276879 298695 276913 6 VGND
port 614 nsew ground input
rlabel viali s 1317 276879 1340 276913 6 VGND
port 614 nsew ground input
rlabel viali s 1225 276879 1259 276913 6 VGND
port 614 nsew ground input
rlabel viali s 1133 276879 1167 276913 6 VGND
port 614 nsew ground input
rlabel viali s 298753 277967 298787 278001 6 VGND
port 614 nsew ground input
rlabel viali s 298661 277967 298695 278001 6 VGND
port 614 nsew ground input
rlabel viali s 1317 277967 1340 278001 6 VGND
port 614 nsew ground input
rlabel viali s 1225 277967 1259 278001 6 VGND
port 614 nsew ground input
rlabel viali s 1133 277967 1167 278001 6 VGND
port 614 nsew ground input
rlabel viali s 298753 279055 298787 279089 6 VGND
port 614 nsew ground input
rlabel viali s 298661 279055 298695 279089 6 VGND
port 614 nsew ground input
rlabel viali s 1317 279055 1340 279089 6 VGND
port 614 nsew ground input
rlabel viali s 1225 279055 1259 279089 6 VGND
port 614 nsew ground input
rlabel viali s 1133 279055 1167 279089 6 VGND
port 614 nsew ground input
rlabel viali s 298753 280143 298787 280177 6 VGND
port 614 nsew ground input
rlabel viali s 298661 280143 298695 280177 6 VGND
port 614 nsew ground input
rlabel viali s 1317 280143 1340 280177 6 VGND
port 614 nsew ground input
rlabel viali s 1225 280143 1259 280177 6 VGND
port 614 nsew ground input
rlabel viali s 1133 280143 1167 280177 6 VGND
port 614 nsew ground input
rlabel viali s 298753 281231 298787 281265 6 VGND
port 614 nsew ground input
rlabel viali s 298661 281231 298695 281265 6 VGND
port 614 nsew ground input
rlabel viali s 1317 281231 1340 281265 6 VGND
port 614 nsew ground input
rlabel viali s 1225 281231 1259 281265 6 VGND
port 614 nsew ground input
rlabel viali s 1133 281231 1167 281265 6 VGND
port 614 nsew ground input
rlabel viali s 298753 282319 298787 282353 6 VGND
port 614 nsew ground input
rlabel viali s 298661 282319 298695 282353 6 VGND
port 614 nsew ground input
rlabel viali s 1317 282319 1340 282353 6 VGND
port 614 nsew ground input
rlabel viali s 1225 282319 1259 282353 6 VGND
port 614 nsew ground input
rlabel viali s 1133 282319 1167 282353 6 VGND
port 614 nsew ground input
rlabel viali s 298753 283407 298787 283441 6 VGND
port 614 nsew ground input
rlabel viali s 298661 283407 298695 283441 6 VGND
port 614 nsew ground input
rlabel viali s 1317 283407 1340 283441 6 VGND
port 614 nsew ground input
rlabel viali s 1225 283407 1259 283441 6 VGND
port 614 nsew ground input
rlabel viali s 1133 283407 1167 283441 6 VGND
port 614 nsew ground input
rlabel viali s 298753 284495 298787 284529 6 VGND
port 614 nsew ground input
rlabel viali s 298661 284495 298695 284529 6 VGND
port 614 nsew ground input
rlabel viali s 1317 284495 1340 284529 6 VGND
port 614 nsew ground input
rlabel viali s 1225 284495 1259 284529 6 VGND
port 614 nsew ground input
rlabel viali s 1133 284495 1167 284529 6 VGND
port 614 nsew ground input
rlabel viali s 298753 285583 298787 285617 6 VGND
port 614 nsew ground input
rlabel viali s 298661 285583 298695 285617 6 VGND
port 614 nsew ground input
rlabel viali s 1317 285583 1340 285617 6 VGND
port 614 nsew ground input
rlabel viali s 1225 285583 1259 285617 6 VGND
port 614 nsew ground input
rlabel viali s 1133 285583 1167 285617 6 VGND
port 614 nsew ground input
rlabel viali s 298753 286671 298787 286705 6 VGND
port 614 nsew ground input
rlabel viali s 298661 286671 298695 286705 6 VGND
port 614 nsew ground input
rlabel viali s 1317 286671 1340 286705 6 VGND
port 614 nsew ground input
rlabel viali s 1225 286671 1259 286705 6 VGND
port 614 nsew ground input
rlabel viali s 1133 286671 1167 286705 6 VGND
port 614 nsew ground input
rlabel viali s 298753 287759 298787 287793 6 VGND
port 614 nsew ground input
rlabel viali s 298661 287759 298695 287793 6 VGND
port 614 nsew ground input
rlabel viali s 1317 287759 1340 287793 6 VGND
port 614 nsew ground input
rlabel viali s 1225 287759 1259 287793 6 VGND
port 614 nsew ground input
rlabel viali s 1133 287759 1167 287793 6 VGND
port 614 nsew ground input
rlabel viali s 298753 288847 298787 288881 6 VGND
port 614 nsew ground input
rlabel viali s 298661 288847 298695 288881 6 VGND
port 614 nsew ground input
rlabel viali s 1317 288847 1340 288881 6 VGND
port 614 nsew ground input
rlabel viali s 1225 288847 1259 288881 6 VGND
port 614 nsew ground input
rlabel viali s 1133 288847 1167 288881 6 VGND
port 614 nsew ground input
rlabel viali s 298753 289935 298787 289969 6 VGND
port 614 nsew ground input
rlabel viali s 298661 289935 298695 289969 6 VGND
port 614 nsew ground input
rlabel viali s 1317 289935 1340 289969 6 VGND
port 614 nsew ground input
rlabel viali s 1225 289935 1259 289969 6 VGND
port 614 nsew ground input
rlabel viali s 1133 289935 1167 289969 6 VGND
port 614 nsew ground input
rlabel viali s 298753 291023 298787 291057 6 VGND
port 614 nsew ground input
rlabel viali s 298661 291023 298695 291057 6 VGND
port 614 nsew ground input
rlabel viali s 1317 291023 1340 291057 6 VGND
port 614 nsew ground input
rlabel viali s 1225 291023 1259 291057 6 VGND
port 614 nsew ground input
rlabel viali s 1133 291023 1167 291057 6 VGND
port 614 nsew ground input
rlabel viali s 298753 292111 298787 292145 6 VGND
port 614 nsew ground input
rlabel viali s 298661 292111 298695 292145 6 VGND
port 614 nsew ground input
rlabel viali s 1317 292111 1340 292145 6 VGND
port 614 nsew ground input
rlabel viali s 1225 292111 1259 292145 6 VGND
port 614 nsew ground input
rlabel viali s 1133 292111 1167 292145 6 VGND
port 614 nsew ground input
rlabel viali s 298753 293199 298787 293233 6 VGND
port 614 nsew ground input
rlabel viali s 298661 293199 298695 293233 6 VGND
port 614 nsew ground input
rlabel viali s 1317 293199 1340 293233 6 VGND
port 614 nsew ground input
rlabel viali s 1225 293199 1259 293233 6 VGND
port 614 nsew ground input
rlabel viali s 1133 293199 1167 293233 6 VGND
port 614 nsew ground input
rlabel viali s 298753 294287 298787 294321 6 VGND
port 614 nsew ground input
rlabel viali s 298661 294287 298695 294321 6 VGND
port 614 nsew ground input
rlabel viali s 1317 294287 1340 294321 6 VGND
port 614 nsew ground input
rlabel viali s 1225 294287 1259 294321 6 VGND
port 614 nsew ground input
rlabel viali s 1133 294287 1167 294321 6 VGND
port 614 nsew ground input
rlabel viali s 298753 295375 298787 295409 6 VGND
port 614 nsew ground input
rlabel viali s 298661 295375 298695 295409 6 VGND
port 614 nsew ground input
rlabel viali s 1317 295375 1340 295409 6 VGND
port 614 nsew ground input
rlabel viali s 1225 295375 1259 295409 6 VGND
port 614 nsew ground input
rlabel viali s 1133 295375 1167 295409 6 VGND
port 614 nsew ground input
rlabel viali s 298753 296463 298787 296497 6 VGND
port 614 nsew ground input
rlabel viali s 298661 296463 298695 296497 6 VGND
port 614 nsew ground input
rlabel viali s 1317 296463 1340 296497 6 VGND
port 614 nsew ground input
rlabel viali s 1225 296463 1259 296497 6 VGND
port 614 nsew ground input
rlabel viali s 1133 296463 1167 296497 6 VGND
port 614 nsew ground input
rlabel viali s 298753 297551 298787 297585 6 VGND
port 614 nsew ground input
rlabel viali s 298661 297551 298695 297585 6 VGND
port 614 nsew ground input
rlabel viali s 1317 297551 1340 297585 6 VGND
port 614 nsew ground input
rlabel viali s 1225 297551 1259 297585 6 VGND
port 614 nsew ground input
rlabel viali s 1133 297551 1167 297585 6 VGND
port 614 nsew ground input
rlabel locali s 298695 2445 298799 2553 6 VGND
port 614 nsew ground input
rlabel locali s 1121 2445 1225 2553 6 VGND
port 614 nsew ground input
rlabel locali s 298660 2553 298799 2703 6 VGND
port 614 nsew ground input
rlabel locali s 298660 2703 298816 2737 6 VGND
port 614 nsew ground input
rlabel locali s 298660 2737 298799 2887 6 VGND
port 614 nsew ground input
rlabel locali s 1121 2553 1340 2703 6 VGND
port 614 nsew ground input
rlabel locali s 1104 2703 1340 2737 6 VGND
port 614 nsew ground input
rlabel locali s 1121 2737 1340 2887 6 VGND
port 614 nsew ground input
rlabel locali s 298695 2887 298799 2995 6 VGND
port 614 nsew ground input
rlabel locali s 1121 2887 1225 2995 6 VGND
port 614 nsew ground input
rlabel locali s 298695 3533 298799 3641 6 VGND
port 614 nsew ground input
rlabel locali s 1121 3533 1225 3641 6 VGND
port 614 nsew ground input
rlabel locali s 298660 3641 298799 3791 6 VGND
port 614 nsew ground input
rlabel locali s 298660 3791 298816 3825 6 VGND
port 614 nsew ground input
rlabel locali s 298660 3825 298799 3975 6 VGND
port 614 nsew ground input
rlabel locali s 1121 3641 1340 3791 6 VGND
port 614 nsew ground input
rlabel locali s 1104 3791 1340 3825 6 VGND
port 614 nsew ground input
rlabel locali s 1121 3825 1340 3975 6 VGND
port 614 nsew ground input
rlabel locali s 298695 3975 298799 4083 6 VGND
port 614 nsew ground input
rlabel locali s 1121 3975 1225 4083 6 VGND
port 614 nsew ground input
rlabel locali s 298695 4621 298799 4729 6 VGND
port 614 nsew ground input
rlabel locali s 1121 4621 1225 4729 6 VGND
port 614 nsew ground input
rlabel locali s 298660 4729 298799 4879 6 VGND
port 614 nsew ground input
rlabel locali s 298660 4879 298816 4913 6 VGND
port 614 nsew ground input
rlabel locali s 298660 4913 298799 5063 6 VGND
port 614 nsew ground input
rlabel locali s 1121 4729 1340 4879 6 VGND
port 614 nsew ground input
rlabel locali s 1104 4879 1340 4913 6 VGND
port 614 nsew ground input
rlabel locali s 1121 4913 1340 5063 6 VGND
port 614 nsew ground input
rlabel locali s 298695 5063 298799 5171 6 VGND
port 614 nsew ground input
rlabel locali s 1121 5063 1225 5171 6 VGND
port 614 nsew ground input
rlabel locali s 298695 5709 298799 5817 6 VGND
port 614 nsew ground input
rlabel locali s 1121 5709 1225 5817 6 VGND
port 614 nsew ground input
rlabel locali s 298660 5817 298799 5967 6 VGND
port 614 nsew ground input
rlabel locali s 298660 5967 298816 6001 6 VGND
port 614 nsew ground input
rlabel locali s 298660 6001 298799 6151 6 VGND
port 614 nsew ground input
rlabel locali s 1121 5817 1340 5967 6 VGND
port 614 nsew ground input
rlabel locali s 1104 5967 1340 6001 6 VGND
port 614 nsew ground input
rlabel locali s 1121 6001 1340 6151 6 VGND
port 614 nsew ground input
rlabel locali s 298695 6151 298799 6259 6 VGND
port 614 nsew ground input
rlabel locali s 1121 6151 1225 6259 6 VGND
port 614 nsew ground input
rlabel locali s 298695 6797 298799 6905 6 VGND
port 614 nsew ground input
rlabel locali s 1121 6797 1225 6905 6 VGND
port 614 nsew ground input
rlabel locali s 298660 6905 298799 7055 6 VGND
port 614 nsew ground input
rlabel locali s 298660 7055 298816 7089 6 VGND
port 614 nsew ground input
rlabel locali s 298660 7089 298799 7239 6 VGND
port 614 nsew ground input
rlabel locali s 1121 6905 1340 7055 6 VGND
port 614 nsew ground input
rlabel locali s 1104 7055 1340 7089 6 VGND
port 614 nsew ground input
rlabel locali s 1121 7089 1340 7239 6 VGND
port 614 nsew ground input
rlabel locali s 298695 7239 298799 7347 6 VGND
port 614 nsew ground input
rlabel locali s 1121 7239 1225 7347 6 VGND
port 614 nsew ground input
rlabel locali s 298695 7885 298799 7993 6 VGND
port 614 nsew ground input
rlabel locali s 1121 7885 1225 7993 6 VGND
port 614 nsew ground input
rlabel locali s 298660 7993 298799 8143 6 VGND
port 614 nsew ground input
rlabel locali s 298660 8143 298816 8177 6 VGND
port 614 nsew ground input
rlabel locali s 298660 8177 298799 8327 6 VGND
port 614 nsew ground input
rlabel locali s 1121 7993 1340 8143 6 VGND
port 614 nsew ground input
rlabel locali s 1104 8143 1340 8177 6 VGND
port 614 nsew ground input
rlabel locali s 1121 8177 1340 8327 6 VGND
port 614 nsew ground input
rlabel locali s 298695 8327 298799 8435 6 VGND
port 614 nsew ground input
rlabel locali s 1121 8327 1225 8435 6 VGND
port 614 nsew ground input
rlabel locali s 298695 8973 298799 9081 6 VGND
port 614 nsew ground input
rlabel locali s 1121 8973 1225 9081 6 VGND
port 614 nsew ground input
rlabel locali s 298660 9081 298799 9231 6 VGND
port 614 nsew ground input
rlabel locali s 298660 9231 298816 9265 6 VGND
port 614 nsew ground input
rlabel locali s 298660 9265 298799 9415 6 VGND
port 614 nsew ground input
rlabel locali s 1121 9081 1340 9231 6 VGND
port 614 nsew ground input
rlabel locali s 1104 9231 1340 9265 6 VGND
port 614 nsew ground input
rlabel locali s 1121 9265 1340 9415 6 VGND
port 614 nsew ground input
rlabel locali s 298695 9415 298799 9523 6 VGND
port 614 nsew ground input
rlabel locali s 1121 9415 1225 9523 6 VGND
port 614 nsew ground input
rlabel locali s 298695 10061 298799 10169 6 VGND
port 614 nsew ground input
rlabel locali s 1121 10061 1225 10169 6 VGND
port 614 nsew ground input
rlabel locali s 298660 10169 298799 10319 6 VGND
port 614 nsew ground input
rlabel locali s 298660 10319 298816 10353 6 VGND
port 614 nsew ground input
rlabel locali s 298660 10353 298799 10503 6 VGND
port 614 nsew ground input
rlabel locali s 1121 10169 1340 10319 6 VGND
port 614 nsew ground input
rlabel locali s 1104 10319 1340 10353 6 VGND
port 614 nsew ground input
rlabel locali s 1121 10353 1340 10503 6 VGND
port 614 nsew ground input
rlabel locali s 298695 10503 298799 10611 6 VGND
port 614 nsew ground input
rlabel locali s 1121 10503 1225 10611 6 VGND
port 614 nsew ground input
rlabel locali s 298695 11149 298799 11257 6 VGND
port 614 nsew ground input
rlabel locali s 1121 11149 1225 11257 6 VGND
port 614 nsew ground input
rlabel locali s 298660 11257 298799 11407 6 VGND
port 614 nsew ground input
rlabel locali s 298660 11407 298816 11441 6 VGND
port 614 nsew ground input
rlabel locali s 298660 11441 298799 11591 6 VGND
port 614 nsew ground input
rlabel locali s 1121 11257 1340 11407 6 VGND
port 614 nsew ground input
rlabel locali s 1104 11407 1340 11441 6 VGND
port 614 nsew ground input
rlabel locali s 1121 11441 1340 11591 6 VGND
port 614 nsew ground input
rlabel locali s 298695 11591 298799 11699 6 VGND
port 614 nsew ground input
rlabel locali s 1121 11591 1225 11699 6 VGND
port 614 nsew ground input
rlabel locali s 298695 12237 298799 12345 6 VGND
port 614 nsew ground input
rlabel locali s 1121 12237 1225 12345 6 VGND
port 614 nsew ground input
rlabel locali s 298660 12345 298799 12495 6 VGND
port 614 nsew ground input
rlabel locali s 298660 12495 298816 12529 6 VGND
port 614 nsew ground input
rlabel locali s 298660 12529 298799 12679 6 VGND
port 614 nsew ground input
rlabel locali s 1121 12345 1340 12495 6 VGND
port 614 nsew ground input
rlabel locali s 1104 12495 1340 12529 6 VGND
port 614 nsew ground input
rlabel locali s 1121 12529 1340 12679 6 VGND
port 614 nsew ground input
rlabel locali s 298695 12679 298799 12787 6 VGND
port 614 nsew ground input
rlabel locali s 1121 12679 1225 12787 6 VGND
port 614 nsew ground input
rlabel locali s 298695 13325 298799 13433 6 VGND
port 614 nsew ground input
rlabel locali s 1121 13325 1225 13433 6 VGND
port 614 nsew ground input
rlabel locali s 298660 13433 298799 13583 6 VGND
port 614 nsew ground input
rlabel locali s 298660 13583 298816 13617 6 VGND
port 614 nsew ground input
rlabel locali s 298660 13617 298799 13767 6 VGND
port 614 nsew ground input
rlabel locali s 1121 13433 1340 13583 6 VGND
port 614 nsew ground input
rlabel locali s 1104 13583 1340 13617 6 VGND
port 614 nsew ground input
rlabel locali s 1121 13617 1340 13767 6 VGND
port 614 nsew ground input
rlabel locali s 298695 13767 298799 13875 6 VGND
port 614 nsew ground input
rlabel locali s 1121 13767 1225 13875 6 VGND
port 614 nsew ground input
rlabel locali s 298695 14413 298799 14521 6 VGND
port 614 nsew ground input
rlabel locali s 1121 14413 1225 14521 6 VGND
port 614 nsew ground input
rlabel locali s 298660 14521 298799 14671 6 VGND
port 614 nsew ground input
rlabel locali s 298660 14671 298816 14705 6 VGND
port 614 nsew ground input
rlabel locali s 298660 14705 298799 14855 6 VGND
port 614 nsew ground input
rlabel locali s 1121 14521 1340 14671 6 VGND
port 614 nsew ground input
rlabel locali s 1104 14671 1340 14705 6 VGND
port 614 nsew ground input
rlabel locali s 1121 14705 1340 14855 6 VGND
port 614 nsew ground input
rlabel locali s 298695 14855 298799 14963 6 VGND
port 614 nsew ground input
rlabel locali s 1121 14855 1225 14963 6 VGND
port 614 nsew ground input
rlabel locali s 298695 15501 298799 15609 6 VGND
port 614 nsew ground input
rlabel locali s 1121 15501 1225 15609 6 VGND
port 614 nsew ground input
rlabel locali s 298660 15609 298799 15759 6 VGND
port 614 nsew ground input
rlabel locali s 298660 15759 298816 15793 6 VGND
port 614 nsew ground input
rlabel locali s 298660 15793 298799 15943 6 VGND
port 614 nsew ground input
rlabel locali s 1121 15609 1340 15759 6 VGND
port 614 nsew ground input
rlabel locali s 1104 15759 1340 15793 6 VGND
port 614 nsew ground input
rlabel locali s 1121 15793 1340 15943 6 VGND
port 614 nsew ground input
rlabel locali s 298695 15943 298799 16051 6 VGND
port 614 nsew ground input
rlabel locali s 1121 15943 1225 16051 6 VGND
port 614 nsew ground input
rlabel locali s 298695 16589 298799 16697 6 VGND
port 614 nsew ground input
rlabel locali s 1121 16589 1225 16697 6 VGND
port 614 nsew ground input
rlabel locali s 298660 16697 298799 16847 6 VGND
port 614 nsew ground input
rlabel locali s 298660 16847 298816 16881 6 VGND
port 614 nsew ground input
rlabel locali s 298660 16881 298799 17031 6 VGND
port 614 nsew ground input
rlabel locali s 1121 16697 1340 16847 6 VGND
port 614 nsew ground input
rlabel locali s 1104 16847 1340 16881 6 VGND
port 614 nsew ground input
rlabel locali s 1121 16881 1340 17031 6 VGND
port 614 nsew ground input
rlabel locali s 298695 17031 298799 17139 6 VGND
port 614 nsew ground input
rlabel locali s 1121 17031 1225 17139 6 VGND
port 614 nsew ground input
rlabel locali s 298695 17677 298799 17785 6 VGND
port 614 nsew ground input
rlabel locali s 1121 17677 1225 17785 6 VGND
port 614 nsew ground input
rlabel locali s 298660 17785 298799 17935 6 VGND
port 614 nsew ground input
rlabel locali s 298660 17935 298816 17969 6 VGND
port 614 nsew ground input
rlabel locali s 298660 17969 298799 18119 6 VGND
port 614 nsew ground input
rlabel locali s 1121 17785 1340 17935 6 VGND
port 614 nsew ground input
rlabel locali s 1104 17935 1340 17969 6 VGND
port 614 nsew ground input
rlabel locali s 1121 17969 1340 18119 6 VGND
port 614 nsew ground input
rlabel locali s 298695 18119 298799 18227 6 VGND
port 614 nsew ground input
rlabel locali s 1121 18119 1225 18227 6 VGND
port 614 nsew ground input
rlabel locali s 298695 18765 298799 18873 6 VGND
port 614 nsew ground input
rlabel locali s 1121 18765 1225 18873 6 VGND
port 614 nsew ground input
rlabel locali s 298660 18873 298799 19023 6 VGND
port 614 nsew ground input
rlabel locali s 298660 19023 298816 19057 6 VGND
port 614 nsew ground input
rlabel locali s 298660 19057 298799 19207 6 VGND
port 614 nsew ground input
rlabel locali s 1121 18873 1340 19023 6 VGND
port 614 nsew ground input
rlabel locali s 1104 19023 1340 19057 6 VGND
port 614 nsew ground input
rlabel locali s 1121 19057 1340 19207 6 VGND
port 614 nsew ground input
rlabel locali s 298695 19207 298799 19315 6 VGND
port 614 nsew ground input
rlabel locali s 1121 19207 1225 19315 6 VGND
port 614 nsew ground input
rlabel locali s 298695 19853 298799 19961 6 VGND
port 614 nsew ground input
rlabel locali s 1121 19853 1225 19961 6 VGND
port 614 nsew ground input
rlabel locali s 298660 19961 298799 20111 6 VGND
port 614 nsew ground input
rlabel locali s 298660 20111 298816 20145 6 VGND
port 614 nsew ground input
rlabel locali s 298660 20145 298799 20295 6 VGND
port 614 nsew ground input
rlabel locali s 1121 19961 1340 20111 6 VGND
port 614 nsew ground input
rlabel locali s 1104 20111 1340 20145 6 VGND
port 614 nsew ground input
rlabel locali s 1121 20145 1340 20295 6 VGND
port 614 nsew ground input
rlabel locali s 298695 20295 298799 20403 6 VGND
port 614 nsew ground input
rlabel locali s 1121 20295 1225 20403 6 VGND
port 614 nsew ground input
rlabel locali s 298695 20941 298799 21049 6 VGND
port 614 nsew ground input
rlabel locali s 1121 20941 1225 21049 6 VGND
port 614 nsew ground input
rlabel locali s 298660 21049 298799 21199 6 VGND
port 614 nsew ground input
rlabel locali s 298660 21199 298816 21233 6 VGND
port 614 nsew ground input
rlabel locali s 298660 21233 298799 21383 6 VGND
port 614 nsew ground input
rlabel locali s 1121 21049 1340 21199 6 VGND
port 614 nsew ground input
rlabel locali s 1104 21199 1340 21233 6 VGND
port 614 nsew ground input
rlabel locali s 1121 21233 1340 21383 6 VGND
port 614 nsew ground input
rlabel locali s 298695 21383 298799 21491 6 VGND
port 614 nsew ground input
rlabel locali s 1121 21383 1225 21491 6 VGND
port 614 nsew ground input
rlabel locali s 298695 22029 298799 22137 6 VGND
port 614 nsew ground input
rlabel locali s 1121 22029 1225 22137 6 VGND
port 614 nsew ground input
rlabel locali s 298660 22137 298799 22287 6 VGND
port 614 nsew ground input
rlabel locali s 298660 22287 298816 22321 6 VGND
port 614 nsew ground input
rlabel locali s 298660 22321 298799 22471 6 VGND
port 614 nsew ground input
rlabel locali s 1121 22137 1340 22287 6 VGND
port 614 nsew ground input
rlabel locali s 1104 22287 1340 22321 6 VGND
port 614 nsew ground input
rlabel locali s 1121 22321 1340 22471 6 VGND
port 614 nsew ground input
rlabel locali s 298695 22471 298799 22579 6 VGND
port 614 nsew ground input
rlabel locali s 1121 22471 1225 22579 6 VGND
port 614 nsew ground input
rlabel locali s 298695 23117 298799 23225 6 VGND
port 614 nsew ground input
rlabel locali s 1121 23117 1225 23225 6 VGND
port 614 nsew ground input
rlabel locali s 298660 23225 298799 23375 6 VGND
port 614 nsew ground input
rlabel locali s 298660 23375 298816 23409 6 VGND
port 614 nsew ground input
rlabel locali s 298660 23409 298799 23559 6 VGND
port 614 nsew ground input
rlabel locali s 1121 23225 1340 23375 6 VGND
port 614 nsew ground input
rlabel locali s 1104 23375 1340 23409 6 VGND
port 614 nsew ground input
rlabel locali s 1121 23409 1340 23559 6 VGND
port 614 nsew ground input
rlabel locali s 298695 23559 298799 23667 6 VGND
port 614 nsew ground input
rlabel locali s 1121 23559 1225 23667 6 VGND
port 614 nsew ground input
rlabel locali s 298695 24205 298799 24313 6 VGND
port 614 nsew ground input
rlabel locali s 1121 24205 1225 24313 6 VGND
port 614 nsew ground input
rlabel locali s 298660 24313 298799 24463 6 VGND
port 614 nsew ground input
rlabel locali s 298660 24463 298816 24497 6 VGND
port 614 nsew ground input
rlabel locali s 298660 24497 298799 24647 6 VGND
port 614 nsew ground input
rlabel locali s 1121 24313 1340 24463 6 VGND
port 614 nsew ground input
rlabel locali s 1104 24463 1340 24497 6 VGND
port 614 nsew ground input
rlabel locali s 1121 24497 1340 24647 6 VGND
port 614 nsew ground input
rlabel locali s 298695 24647 298799 24755 6 VGND
port 614 nsew ground input
rlabel locali s 1121 24647 1225 24755 6 VGND
port 614 nsew ground input
rlabel locali s 298695 25293 298799 25401 6 VGND
port 614 nsew ground input
rlabel locali s 1121 25293 1225 25401 6 VGND
port 614 nsew ground input
rlabel locali s 298660 25401 298799 25551 6 VGND
port 614 nsew ground input
rlabel locali s 298660 25551 298816 25585 6 VGND
port 614 nsew ground input
rlabel locali s 298660 25585 298799 25735 6 VGND
port 614 nsew ground input
rlabel locali s 1121 25401 1340 25551 6 VGND
port 614 nsew ground input
rlabel locali s 1104 25551 1340 25585 6 VGND
port 614 nsew ground input
rlabel locali s 1121 25585 1340 25735 6 VGND
port 614 nsew ground input
rlabel locali s 298695 25735 298799 25843 6 VGND
port 614 nsew ground input
rlabel locali s 1121 25735 1225 25843 6 VGND
port 614 nsew ground input
rlabel locali s 298695 26381 298799 26489 6 VGND
port 614 nsew ground input
rlabel locali s 1121 26381 1225 26489 6 VGND
port 614 nsew ground input
rlabel locali s 298660 26489 298799 26639 6 VGND
port 614 nsew ground input
rlabel locali s 298660 26639 298816 26673 6 VGND
port 614 nsew ground input
rlabel locali s 298660 26673 298799 26823 6 VGND
port 614 nsew ground input
rlabel locali s 1121 26489 1340 26639 6 VGND
port 614 nsew ground input
rlabel locali s 1104 26639 1340 26673 6 VGND
port 614 nsew ground input
rlabel locali s 1121 26673 1340 26823 6 VGND
port 614 nsew ground input
rlabel locali s 298695 26823 298799 26931 6 VGND
port 614 nsew ground input
rlabel locali s 1121 26823 1225 26931 6 VGND
port 614 nsew ground input
rlabel locali s 298695 27469 298799 27577 6 VGND
port 614 nsew ground input
rlabel locali s 1121 27469 1225 27577 6 VGND
port 614 nsew ground input
rlabel locali s 298660 27577 298799 27727 6 VGND
port 614 nsew ground input
rlabel locali s 298660 27727 298816 27761 6 VGND
port 614 nsew ground input
rlabel locali s 298660 27761 298799 27911 6 VGND
port 614 nsew ground input
rlabel locali s 1121 27577 1340 27727 6 VGND
port 614 nsew ground input
rlabel locali s 1104 27727 1340 27761 6 VGND
port 614 nsew ground input
rlabel locali s 1121 27761 1340 27911 6 VGND
port 614 nsew ground input
rlabel locali s 298695 27911 298799 28019 6 VGND
port 614 nsew ground input
rlabel locali s 1121 27911 1225 28019 6 VGND
port 614 nsew ground input
rlabel locali s 298695 28557 298799 28665 6 VGND
port 614 nsew ground input
rlabel locali s 1121 28557 1225 28665 6 VGND
port 614 nsew ground input
rlabel locali s 298660 28665 298799 28815 6 VGND
port 614 nsew ground input
rlabel locali s 298660 28815 298816 28849 6 VGND
port 614 nsew ground input
rlabel locali s 298660 28849 298799 28999 6 VGND
port 614 nsew ground input
rlabel locali s 1121 28665 1340 28815 6 VGND
port 614 nsew ground input
rlabel locali s 1104 28815 1340 28849 6 VGND
port 614 nsew ground input
rlabel locali s 1121 28849 1340 28999 6 VGND
port 614 nsew ground input
rlabel locali s 298695 28999 298799 29107 6 VGND
port 614 nsew ground input
rlabel locali s 1121 28999 1225 29107 6 VGND
port 614 nsew ground input
rlabel locali s 298695 29645 298799 29753 6 VGND
port 614 nsew ground input
rlabel locali s 1121 29645 1225 29753 6 VGND
port 614 nsew ground input
rlabel locali s 298660 29753 298799 29903 6 VGND
port 614 nsew ground input
rlabel locali s 298660 29903 298816 29937 6 VGND
port 614 nsew ground input
rlabel locali s 298660 29937 298799 30087 6 VGND
port 614 nsew ground input
rlabel locali s 1121 29753 1340 29903 6 VGND
port 614 nsew ground input
rlabel locali s 1104 29903 1340 29937 6 VGND
port 614 nsew ground input
rlabel locali s 1121 29937 1340 30087 6 VGND
port 614 nsew ground input
rlabel locali s 298695 30087 298799 30195 6 VGND
port 614 nsew ground input
rlabel locali s 1121 30087 1225 30195 6 VGND
port 614 nsew ground input
rlabel locali s 298695 30733 298799 30841 6 VGND
port 614 nsew ground input
rlabel locali s 1121 30733 1225 30841 6 VGND
port 614 nsew ground input
rlabel locali s 298660 30841 298799 30991 6 VGND
port 614 nsew ground input
rlabel locali s 298660 30991 298816 31025 6 VGND
port 614 nsew ground input
rlabel locali s 298660 31025 298799 31175 6 VGND
port 614 nsew ground input
rlabel locali s 1121 30841 1340 30991 6 VGND
port 614 nsew ground input
rlabel locali s 1104 30991 1340 31025 6 VGND
port 614 nsew ground input
rlabel locali s 1121 31025 1340 31175 6 VGND
port 614 nsew ground input
rlabel locali s 298695 31175 298799 31283 6 VGND
port 614 nsew ground input
rlabel locali s 1121 31175 1225 31283 6 VGND
port 614 nsew ground input
rlabel locali s 298695 31821 298799 31929 6 VGND
port 614 nsew ground input
rlabel locali s 1121 31821 1225 31929 6 VGND
port 614 nsew ground input
rlabel locali s 298660 31929 298799 32079 6 VGND
port 614 nsew ground input
rlabel locali s 298660 32079 298816 32113 6 VGND
port 614 nsew ground input
rlabel locali s 298660 32113 298799 32263 6 VGND
port 614 nsew ground input
rlabel locali s 1121 31929 1340 32079 6 VGND
port 614 nsew ground input
rlabel locali s 1104 32079 1340 32113 6 VGND
port 614 nsew ground input
rlabel locali s 1121 32113 1340 32263 6 VGND
port 614 nsew ground input
rlabel locali s 298695 32263 298799 32371 6 VGND
port 614 nsew ground input
rlabel locali s 1121 32263 1225 32371 6 VGND
port 614 nsew ground input
rlabel locali s 298695 32909 298799 33017 6 VGND
port 614 nsew ground input
rlabel locali s 1121 32909 1225 33017 6 VGND
port 614 nsew ground input
rlabel locali s 298660 33017 298799 33167 6 VGND
port 614 nsew ground input
rlabel locali s 298660 33167 298816 33201 6 VGND
port 614 nsew ground input
rlabel locali s 298660 33201 298799 33351 6 VGND
port 614 nsew ground input
rlabel locali s 1121 33017 1340 33167 6 VGND
port 614 nsew ground input
rlabel locali s 1104 33167 1340 33201 6 VGND
port 614 nsew ground input
rlabel locali s 1121 33201 1340 33351 6 VGND
port 614 nsew ground input
rlabel locali s 298695 33351 298799 33459 6 VGND
port 614 nsew ground input
rlabel locali s 1121 33351 1225 33459 6 VGND
port 614 nsew ground input
rlabel locali s 298695 33997 298799 34105 6 VGND
port 614 nsew ground input
rlabel locali s 1121 33997 1225 34105 6 VGND
port 614 nsew ground input
rlabel locali s 298660 34105 298799 34255 6 VGND
port 614 nsew ground input
rlabel locali s 298660 34255 298816 34289 6 VGND
port 614 nsew ground input
rlabel locali s 298660 34289 298799 34439 6 VGND
port 614 nsew ground input
rlabel locali s 1121 34105 1340 34255 6 VGND
port 614 nsew ground input
rlabel locali s 1104 34255 1340 34289 6 VGND
port 614 nsew ground input
rlabel locali s 1121 34289 1340 34439 6 VGND
port 614 nsew ground input
rlabel locali s 298695 34439 298799 34547 6 VGND
port 614 nsew ground input
rlabel locali s 1121 34439 1225 34547 6 VGND
port 614 nsew ground input
rlabel locali s 298695 35085 298799 35193 6 VGND
port 614 nsew ground input
rlabel locali s 1121 35085 1225 35193 6 VGND
port 614 nsew ground input
rlabel locali s 298660 35193 298799 35343 6 VGND
port 614 nsew ground input
rlabel locali s 298660 35343 298816 35377 6 VGND
port 614 nsew ground input
rlabel locali s 298660 35377 298799 35527 6 VGND
port 614 nsew ground input
rlabel locali s 1121 35193 1340 35343 6 VGND
port 614 nsew ground input
rlabel locali s 1104 35343 1340 35377 6 VGND
port 614 nsew ground input
rlabel locali s 1121 35377 1340 35527 6 VGND
port 614 nsew ground input
rlabel locali s 298695 35527 298799 35635 6 VGND
port 614 nsew ground input
rlabel locali s 1121 35527 1225 35635 6 VGND
port 614 nsew ground input
rlabel locali s 298695 36173 298799 36281 6 VGND
port 614 nsew ground input
rlabel locali s 1121 36173 1225 36281 6 VGND
port 614 nsew ground input
rlabel locali s 298660 36281 298799 36431 6 VGND
port 614 nsew ground input
rlabel locali s 298660 36431 298816 36465 6 VGND
port 614 nsew ground input
rlabel locali s 298660 36465 298799 36615 6 VGND
port 614 nsew ground input
rlabel locali s 1121 36281 1340 36431 6 VGND
port 614 nsew ground input
rlabel locali s 1104 36431 1340 36465 6 VGND
port 614 nsew ground input
rlabel locali s 1121 36465 1340 36615 6 VGND
port 614 nsew ground input
rlabel locali s 298695 36615 298799 36723 6 VGND
port 614 nsew ground input
rlabel locali s 1121 36615 1225 36723 6 VGND
port 614 nsew ground input
rlabel locali s 298695 37261 298799 37369 6 VGND
port 614 nsew ground input
rlabel locali s 1121 37261 1225 37369 6 VGND
port 614 nsew ground input
rlabel locali s 298660 37369 298799 37519 6 VGND
port 614 nsew ground input
rlabel locali s 298660 37519 298816 37553 6 VGND
port 614 nsew ground input
rlabel locali s 298660 37553 298799 37703 6 VGND
port 614 nsew ground input
rlabel locali s 1121 37369 1340 37519 6 VGND
port 614 nsew ground input
rlabel locali s 1104 37519 1340 37553 6 VGND
port 614 nsew ground input
rlabel locali s 1121 37553 1340 37703 6 VGND
port 614 nsew ground input
rlabel locali s 298695 37703 298799 37811 6 VGND
port 614 nsew ground input
rlabel locali s 1121 37703 1225 37811 6 VGND
port 614 nsew ground input
rlabel locali s 298695 38349 298799 38457 6 VGND
port 614 nsew ground input
rlabel locali s 1121 38349 1225 38457 6 VGND
port 614 nsew ground input
rlabel locali s 298660 38457 298799 38607 6 VGND
port 614 nsew ground input
rlabel locali s 298660 38607 298816 38641 6 VGND
port 614 nsew ground input
rlabel locali s 298660 38641 298799 38791 6 VGND
port 614 nsew ground input
rlabel locali s 1121 38457 1340 38607 6 VGND
port 614 nsew ground input
rlabel locali s 1104 38607 1340 38641 6 VGND
port 614 nsew ground input
rlabel locali s 1121 38641 1340 38791 6 VGND
port 614 nsew ground input
rlabel locali s 298695 38791 298799 38899 6 VGND
port 614 nsew ground input
rlabel locali s 1121 38791 1225 38899 6 VGND
port 614 nsew ground input
rlabel locali s 298695 39437 298799 39545 6 VGND
port 614 nsew ground input
rlabel locali s 1121 39437 1225 39545 6 VGND
port 614 nsew ground input
rlabel locali s 298660 39545 298799 39695 6 VGND
port 614 nsew ground input
rlabel locali s 298660 39695 298816 39729 6 VGND
port 614 nsew ground input
rlabel locali s 298660 39729 298799 39879 6 VGND
port 614 nsew ground input
rlabel locali s 1121 39545 1340 39695 6 VGND
port 614 nsew ground input
rlabel locali s 1104 39695 1340 39729 6 VGND
port 614 nsew ground input
rlabel locali s 1121 39729 1340 39879 6 VGND
port 614 nsew ground input
rlabel locali s 298695 39879 298799 39987 6 VGND
port 614 nsew ground input
rlabel locali s 1121 39879 1225 39987 6 VGND
port 614 nsew ground input
rlabel locali s 298695 40525 298799 40633 6 VGND
port 614 nsew ground input
rlabel locali s 1121 40525 1225 40633 6 VGND
port 614 nsew ground input
rlabel locali s 298660 40633 298799 40783 6 VGND
port 614 nsew ground input
rlabel locali s 298660 40783 298816 40817 6 VGND
port 614 nsew ground input
rlabel locali s 298660 40817 298799 40967 6 VGND
port 614 nsew ground input
rlabel locali s 1121 40633 1340 40783 6 VGND
port 614 nsew ground input
rlabel locali s 1104 40783 1340 40817 6 VGND
port 614 nsew ground input
rlabel locali s 1121 40817 1340 40967 6 VGND
port 614 nsew ground input
rlabel locali s 298695 40967 298799 41075 6 VGND
port 614 nsew ground input
rlabel locali s 1121 40967 1225 41075 6 VGND
port 614 nsew ground input
rlabel locali s 298695 41613 298799 41721 6 VGND
port 614 nsew ground input
rlabel locali s 1121 41613 1225 41721 6 VGND
port 614 nsew ground input
rlabel locali s 298660 41721 298799 41871 6 VGND
port 614 nsew ground input
rlabel locali s 298660 41871 298816 41905 6 VGND
port 614 nsew ground input
rlabel locali s 298660 41905 298799 42055 6 VGND
port 614 nsew ground input
rlabel locali s 1121 41721 1340 41871 6 VGND
port 614 nsew ground input
rlabel locali s 1104 41871 1340 41905 6 VGND
port 614 nsew ground input
rlabel locali s 1121 41905 1340 42055 6 VGND
port 614 nsew ground input
rlabel locali s 298695 42055 298799 42163 6 VGND
port 614 nsew ground input
rlabel locali s 1121 42055 1225 42163 6 VGND
port 614 nsew ground input
rlabel locali s 298695 42701 298799 42809 6 VGND
port 614 nsew ground input
rlabel locali s 1121 42701 1225 42809 6 VGND
port 614 nsew ground input
rlabel locali s 298660 42809 298799 42959 6 VGND
port 614 nsew ground input
rlabel locali s 298660 42959 298816 42993 6 VGND
port 614 nsew ground input
rlabel locali s 298660 42993 298799 43143 6 VGND
port 614 nsew ground input
rlabel locali s 1121 42809 1340 42959 6 VGND
port 614 nsew ground input
rlabel locali s 1104 42959 1340 42993 6 VGND
port 614 nsew ground input
rlabel locali s 1121 42993 1340 43143 6 VGND
port 614 nsew ground input
rlabel locali s 298695 43143 298799 43251 6 VGND
port 614 nsew ground input
rlabel locali s 1121 43143 1225 43251 6 VGND
port 614 nsew ground input
rlabel locali s 298695 43789 298799 43897 6 VGND
port 614 nsew ground input
rlabel locali s 1121 43789 1225 43897 6 VGND
port 614 nsew ground input
rlabel locali s 298660 43897 298799 44047 6 VGND
port 614 nsew ground input
rlabel locali s 298660 44047 298816 44081 6 VGND
port 614 nsew ground input
rlabel locali s 298660 44081 298799 44231 6 VGND
port 614 nsew ground input
rlabel locali s 1121 43897 1340 44047 6 VGND
port 614 nsew ground input
rlabel locali s 1104 44047 1340 44081 6 VGND
port 614 nsew ground input
rlabel locali s 1121 44081 1340 44231 6 VGND
port 614 nsew ground input
rlabel locali s 298695 44231 298799 44339 6 VGND
port 614 nsew ground input
rlabel locali s 1121 44231 1225 44339 6 VGND
port 614 nsew ground input
rlabel locali s 298695 44877 298799 44985 6 VGND
port 614 nsew ground input
rlabel locali s 1121 44877 1225 44985 6 VGND
port 614 nsew ground input
rlabel locali s 298660 44985 298799 45135 6 VGND
port 614 nsew ground input
rlabel locali s 298660 45135 298816 45169 6 VGND
port 614 nsew ground input
rlabel locali s 298660 45169 298799 45319 6 VGND
port 614 nsew ground input
rlabel locali s 1121 44985 1340 45135 6 VGND
port 614 nsew ground input
rlabel locali s 1104 45135 1340 45169 6 VGND
port 614 nsew ground input
rlabel locali s 1121 45169 1340 45319 6 VGND
port 614 nsew ground input
rlabel locali s 298695 45319 298799 45427 6 VGND
port 614 nsew ground input
rlabel locali s 1121 45319 1225 45427 6 VGND
port 614 nsew ground input
rlabel locali s 298695 45965 298799 46073 6 VGND
port 614 nsew ground input
rlabel locali s 1121 45965 1225 46073 6 VGND
port 614 nsew ground input
rlabel locali s 298660 46073 298799 46223 6 VGND
port 614 nsew ground input
rlabel locali s 298660 46223 298816 46257 6 VGND
port 614 nsew ground input
rlabel locali s 298660 46257 298799 46407 6 VGND
port 614 nsew ground input
rlabel locali s 1121 46073 1340 46223 6 VGND
port 614 nsew ground input
rlabel locali s 1104 46223 1340 46257 6 VGND
port 614 nsew ground input
rlabel locali s 1121 46257 1340 46407 6 VGND
port 614 nsew ground input
rlabel locali s 298695 46407 298799 46515 6 VGND
port 614 nsew ground input
rlabel locali s 1121 46407 1225 46515 6 VGND
port 614 nsew ground input
rlabel locali s 298695 47053 298799 47161 6 VGND
port 614 nsew ground input
rlabel locali s 1121 47053 1225 47161 6 VGND
port 614 nsew ground input
rlabel locali s 298660 47161 298799 47311 6 VGND
port 614 nsew ground input
rlabel locali s 298660 47311 298816 47345 6 VGND
port 614 nsew ground input
rlabel locali s 298660 47345 298799 47495 6 VGND
port 614 nsew ground input
rlabel locali s 1121 47161 1340 47311 6 VGND
port 614 nsew ground input
rlabel locali s 1104 47311 1340 47345 6 VGND
port 614 nsew ground input
rlabel locali s 1121 47345 1340 47495 6 VGND
port 614 nsew ground input
rlabel locali s 298695 47495 298799 47603 6 VGND
port 614 nsew ground input
rlabel locali s 1121 47495 1225 47603 6 VGND
port 614 nsew ground input
rlabel locali s 298695 48141 298799 48249 6 VGND
port 614 nsew ground input
rlabel locali s 1121 48141 1225 48249 6 VGND
port 614 nsew ground input
rlabel locali s 298660 48249 298799 48399 6 VGND
port 614 nsew ground input
rlabel locali s 298660 48399 298816 48433 6 VGND
port 614 nsew ground input
rlabel locali s 298660 48433 298799 48583 6 VGND
port 614 nsew ground input
rlabel locali s 1121 48249 1340 48399 6 VGND
port 614 nsew ground input
rlabel locali s 1104 48399 1340 48433 6 VGND
port 614 nsew ground input
rlabel locali s 1121 48433 1340 48583 6 VGND
port 614 nsew ground input
rlabel locali s 298695 48583 298799 48691 6 VGND
port 614 nsew ground input
rlabel locali s 1121 48583 1225 48691 6 VGND
port 614 nsew ground input
rlabel locali s 298695 49229 298799 49337 6 VGND
port 614 nsew ground input
rlabel locali s 1121 49229 1225 49337 6 VGND
port 614 nsew ground input
rlabel locali s 298660 49337 298799 49487 6 VGND
port 614 nsew ground input
rlabel locali s 298660 49487 298816 49521 6 VGND
port 614 nsew ground input
rlabel locali s 298660 49521 298799 49671 6 VGND
port 614 nsew ground input
rlabel locali s 1121 49337 1340 49487 6 VGND
port 614 nsew ground input
rlabel locali s 1104 49487 1340 49521 6 VGND
port 614 nsew ground input
rlabel locali s 1121 49521 1340 49671 6 VGND
port 614 nsew ground input
rlabel locali s 298695 49671 298799 49779 6 VGND
port 614 nsew ground input
rlabel locali s 1121 49671 1225 49779 6 VGND
port 614 nsew ground input
rlabel locali s 298695 50317 298799 50425 6 VGND
port 614 nsew ground input
rlabel locali s 1121 50317 1225 50425 6 VGND
port 614 nsew ground input
rlabel locali s 298660 50425 298799 50575 6 VGND
port 614 nsew ground input
rlabel locali s 298660 50575 298816 50609 6 VGND
port 614 nsew ground input
rlabel locali s 298660 50609 298799 50759 6 VGND
port 614 nsew ground input
rlabel locali s 1121 50425 1340 50575 6 VGND
port 614 nsew ground input
rlabel locali s 1104 50575 1340 50609 6 VGND
port 614 nsew ground input
rlabel locali s 1121 50609 1340 50759 6 VGND
port 614 nsew ground input
rlabel locali s 298695 50759 298799 50867 6 VGND
port 614 nsew ground input
rlabel locali s 1121 50759 1225 50867 6 VGND
port 614 nsew ground input
rlabel locali s 298695 51405 298799 51513 6 VGND
port 614 nsew ground input
rlabel locali s 1121 51405 1225 51513 6 VGND
port 614 nsew ground input
rlabel locali s 298660 51513 298799 51663 6 VGND
port 614 nsew ground input
rlabel locali s 298660 51663 298816 51697 6 VGND
port 614 nsew ground input
rlabel locali s 298660 51697 298799 51847 6 VGND
port 614 nsew ground input
rlabel locali s 1121 51513 1340 51663 6 VGND
port 614 nsew ground input
rlabel locali s 1104 51663 1340 51697 6 VGND
port 614 nsew ground input
rlabel locali s 1121 51697 1340 51847 6 VGND
port 614 nsew ground input
rlabel locali s 298695 51847 298799 51955 6 VGND
port 614 nsew ground input
rlabel locali s 1121 51847 1225 51955 6 VGND
port 614 nsew ground input
rlabel locali s 298695 52493 298799 52601 6 VGND
port 614 nsew ground input
rlabel locali s 1121 52493 1225 52601 6 VGND
port 614 nsew ground input
rlabel locali s 298660 52601 298799 52751 6 VGND
port 614 nsew ground input
rlabel locali s 298660 52751 298816 52785 6 VGND
port 614 nsew ground input
rlabel locali s 298660 52785 298799 52935 6 VGND
port 614 nsew ground input
rlabel locali s 1121 52601 1340 52751 6 VGND
port 614 nsew ground input
rlabel locali s 1104 52751 1340 52785 6 VGND
port 614 nsew ground input
rlabel locali s 1121 52785 1340 52935 6 VGND
port 614 nsew ground input
rlabel locali s 298695 52935 298799 53043 6 VGND
port 614 nsew ground input
rlabel locali s 1121 52935 1225 53043 6 VGND
port 614 nsew ground input
rlabel locali s 298695 53581 298799 53689 6 VGND
port 614 nsew ground input
rlabel locali s 1121 53581 1225 53689 6 VGND
port 614 nsew ground input
rlabel locali s 298660 53689 298799 53839 6 VGND
port 614 nsew ground input
rlabel locali s 298660 53839 298816 53873 6 VGND
port 614 nsew ground input
rlabel locali s 298660 53873 298799 54023 6 VGND
port 614 nsew ground input
rlabel locali s 1121 53689 1340 53839 6 VGND
port 614 nsew ground input
rlabel locali s 1104 53839 1340 53873 6 VGND
port 614 nsew ground input
rlabel locali s 1121 53873 1340 54023 6 VGND
port 614 nsew ground input
rlabel locali s 298695 54023 298799 54131 6 VGND
port 614 nsew ground input
rlabel locali s 1121 54023 1225 54131 6 VGND
port 614 nsew ground input
rlabel locali s 298695 54669 298799 54777 6 VGND
port 614 nsew ground input
rlabel locali s 1121 54669 1225 54777 6 VGND
port 614 nsew ground input
rlabel locali s 298660 54777 298799 54927 6 VGND
port 614 nsew ground input
rlabel locali s 298660 54927 298816 54961 6 VGND
port 614 nsew ground input
rlabel locali s 298660 54961 298799 55111 6 VGND
port 614 nsew ground input
rlabel locali s 1121 54777 1340 54927 6 VGND
port 614 nsew ground input
rlabel locali s 1104 54927 1340 54961 6 VGND
port 614 nsew ground input
rlabel locali s 1121 54961 1340 55111 6 VGND
port 614 nsew ground input
rlabel locali s 298695 55111 298799 55219 6 VGND
port 614 nsew ground input
rlabel locali s 1121 55111 1225 55219 6 VGND
port 614 nsew ground input
rlabel locali s 298695 55757 298799 55865 6 VGND
port 614 nsew ground input
rlabel locali s 1121 55757 1225 55865 6 VGND
port 614 nsew ground input
rlabel locali s 298660 55865 298799 56015 6 VGND
port 614 nsew ground input
rlabel locali s 298660 56015 298816 56049 6 VGND
port 614 nsew ground input
rlabel locali s 298660 56049 298799 56199 6 VGND
port 614 nsew ground input
rlabel locali s 1121 55865 1340 56015 6 VGND
port 614 nsew ground input
rlabel locali s 1104 56015 1340 56049 6 VGND
port 614 nsew ground input
rlabel locali s 1121 56049 1340 56199 6 VGND
port 614 nsew ground input
rlabel locali s 298695 56199 298799 56307 6 VGND
port 614 nsew ground input
rlabel locali s 1121 56199 1225 56307 6 VGND
port 614 nsew ground input
rlabel locali s 298695 56845 298799 56953 6 VGND
port 614 nsew ground input
rlabel locali s 1121 56845 1225 56953 6 VGND
port 614 nsew ground input
rlabel locali s 298660 56953 298799 57103 6 VGND
port 614 nsew ground input
rlabel locali s 298660 57103 298816 57137 6 VGND
port 614 nsew ground input
rlabel locali s 298660 57137 298799 57287 6 VGND
port 614 nsew ground input
rlabel locali s 1121 56953 1340 57103 6 VGND
port 614 nsew ground input
rlabel locali s 1104 57103 1340 57137 6 VGND
port 614 nsew ground input
rlabel locali s 1121 57137 1340 57287 6 VGND
port 614 nsew ground input
rlabel locali s 298695 57287 298799 57395 6 VGND
port 614 nsew ground input
rlabel locali s 1121 57287 1225 57395 6 VGND
port 614 nsew ground input
rlabel locali s 298695 57933 298799 58041 6 VGND
port 614 nsew ground input
rlabel locali s 1121 57933 1225 58041 6 VGND
port 614 nsew ground input
rlabel locali s 298660 58041 298799 58191 6 VGND
port 614 nsew ground input
rlabel locali s 298660 58191 298816 58225 6 VGND
port 614 nsew ground input
rlabel locali s 298660 58225 298799 58375 6 VGND
port 614 nsew ground input
rlabel locali s 1121 58041 1340 58191 6 VGND
port 614 nsew ground input
rlabel locali s 1104 58191 1340 58225 6 VGND
port 614 nsew ground input
rlabel locali s 1121 58225 1340 58375 6 VGND
port 614 nsew ground input
rlabel locali s 298695 58375 298799 58483 6 VGND
port 614 nsew ground input
rlabel locali s 1121 58375 1225 58483 6 VGND
port 614 nsew ground input
rlabel locali s 298695 59021 298799 59129 6 VGND
port 614 nsew ground input
rlabel locali s 1121 59021 1225 59129 6 VGND
port 614 nsew ground input
rlabel locali s 298660 59129 298799 59279 6 VGND
port 614 nsew ground input
rlabel locali s 298660 59279 298816 59313 6 VGND
port 614 nsew ground input
rlabel locali s 298660 59313 298799 59463 6 VGND
port 614 nsew ground input
rlabel locali s 1121 59129 1340 59279 6 VGND
port 614 nsew ground input
rlabel locali s 1104 59279 1340 59313 6 VGND
port 614 nsew ground input
rlabel locali s 1121 59313 1340 59463 6 VGND
port 614 nsew ground input
rlabel locali s 298695 59463 298799 59571 6 VGND
port 614 nsew ground input
rlabel locali s 1121 59463 1225 59571 6 VGND
port 614 nsew ground input
rlabel locali s 298695 60109 298799 60217 6 VGND
port 614 nsew ground input
rlabel locali s 1121 60109 1225 60217 6 VGND
port 614 nsew ground input
rlabel locali s 298660 60217 298799 60367 6 VGND
port 614 nsew ground input
rlabel locali s 298660 60367 298816 60401 6 VGND
port 614 nsew ground input
rlabel locali s 298660 60401 298799 60551 6 VGND
port 614 nsew ground input
rlabel locali s 1121 60217 1340 60367 6 VGND
port 614 nsew ground input
rlabel locali s 1104 60367 1340 60401 6 VGND
port 614 nsew ground input
rlabel locali s 1121 60401 1340 60551 6 VGND
port 614 nsew ground input
rlabel locali s 298695 60551 298799 60659 6 VGND
port 614 nsew ground input
rlabel locali s 1121 60551 1225 60659 6 VGND
port 614 nsew ground input
rlabel locali s 298695 61197 298799 61305 6 VGND
port 614 nsew ground input
rlabel locali s 1121 61197 1225 61305 6 VGND
port 614 nsew ground input
rlabel locali s 298660 61305 298799 61455 6 VGND
port 614 nsew ground input
rlabel locali s 298660 61455 298816 61489 6 VGND
port 614 nsew ground input
rlabel locali s 298660 61489 298799 61639 6 VGND
port 614 nsew ground input
rlabel locali s 1121 61305 1340 61455 6 VGND
port 614 nsew ground input
rlabel locali s 1104 61455 1340 61489 6 VGND
port 614 nsew ground input
rlabel locali s 1121 61489 1340 61639 6 VGND
port 614 nsew ground input
rlabel locali s 298695 61639 298799 61747 6 VGND
port 614 nsew ground input
rlabel locali s 1121 61639 1225 61747 6 VGND
port 614 nsew ground input
rlabel locali s 298695 62285 298799 62393 6 VGND
port 614 nsew ground input
rlabel locali s 1121 62285 1225 62393 6 VGND
port 614 nsew ground input
rlabel locali s 298660 62393 298799 62543 6 VGND
port 614 nsew ground input
rlabel locali s 298660 62543 298816 62577 6 VGND
port 614 nsew ground input
rlabel locali s 298660 62577 298799 62727 6 VGND
port 614 nsew ground input
rlabel locali s 1121 62393 1340 62543 6 VGND
port 614 nsew ground input
rlabel locali s 1104 62543 1340 62577 6 VGND
port 614 nsew ground input
rlabel locali s 1121 62577 1340 62727 6 VGND
port 614 nsew ground input
rlabel locali s 298695 62727 298799 62835 6 VGND
port 614 nsew ground input
rlabel locali s 1121 62727 1225 62835 6 VGND
port 614 nsew ground input
rlabel locali s 298695 63373 298799 63481 6 VGND
port 614 nsew ground input
rlabel locali s 1121 63373 1225 63481 6 VGND
port 614 nsew ground input
rlabel locali s 298660 63481 298799 63631 6 VGND
port 614 nsew ground input
rlabel locali s 298660 63631 298816 63665 6 VGND
port 614 nsew ground input
rlabel locali s 298660 63665 298799 63815 6 VGND
port 614 nsew ground input
rlabel locali s 1121 63481 1340 63631 6 VGND
port 614 nsew ground input
rlabel locali s 1104 63631 1340 63665 6 VGND
port 614 nsew ground input
rlabel locali s 1121 63665 1340 63815 6 VGND
port 614 nsew ground input
rlabel locali s 298695 63815 298799 63923 6 VGND
port 614 nsew ground input
rlabel locali s 1121 63815 1225 63923 6 VGND
port 614 nsew ground input
rlabel locali s 298695 64461 298799 64569 6 VGND
port 614 nsew ground input
rlabel locali s 1121 64461 1225 64569 6 VGND
port 614 nsew ground input
rlabel locali s 298660 64569 298799 64719 6 VGND
port 614 nsew ground input
rlabel locali s 298660 64719 298816 64753 6 VGND
port 614 nsew ground input
rlabel locali s 298660 64753 298799 64903 6 VGND
port 614 nsew ground input
rlabel locali s 1121 64569 1340 64719 6 VGND
port 614 nsew ground input
rlabel locali s 1104 64719 1340 64753 6 VGND
port 614 nsew ground input
rlabel locali s 1121 64753 1340 64903 6 VGND
port 614 nsew ground input
rlabel locali s 298695 64903 298799 65011 6 VGND
port 614 nsew ground input
rlabel locali s 1121 64903 1225 65011 6 VGND
port 614 nsew ground input
rlabel locali s 298695 65549 298799 65657 6 VGND
port 614 nsew ground input
rlabel locali s 1121 65549 1225 65657 6 VGND
port 614 nsew ground input
rlabel locali s 298660 65657 298799 65807 6 VGND
port 614 nsew ground input
rlabel locali s 298660 65807 298816 65841 6 VGND
port 614 nsew ground input
rlabel locali s 298660 65841 298799 65991 6 VGND
port 614 nsew ground input
rlabel locali s 1121 65657 1340 65807 6 VGND
port 614 nsew ground input
rlabel locali s 1104 65807 1340 65841 6 VGND
port 614 nsew ground input
rlabel locali s 1121 65841 1340 65991 6 VGND
port 614 nsew ground input
rlabel locali s 298695 65991 298799 66099 6 VGND
port 614 nsew ground input
rlabel locali s 1121 65991 1225 66099 6 VGND
port 614 nsew ground input
rlabel locali s 298695 66637 298799 66745 6 VGND
port 614 nsew ground input
rlabel locali s 1121 66637 1225 66745 6 VGND
port 614 nsew ground input
rlabel locali s 298660 66745 298799 66895 6 VGND
port 614 nsew ground input
rlabel locali s 298660 66895 298816 66929 6 VGND
port 614 nsew ground input
rlabel locali s 298660 66929 298799 67079 6 VGND
port 614 nsew ground input
rlabel locali s 1121 66745 1340 66895 6 VGND
port 614 nsew ground input
rlabel locali s 1104 66895 1340 66929 6 VGND
port 614 nsew ground input
rlabel locali s 1121 66929 1340 67079 6 VGND
port 614 nsew ground input
rlabel locali s 298695 67079 298799 67187 6 VGND
port 614 nsew ground input
rlabel locali s 1121 67079 1225 67187 6 VGND
port 614 nsew ground input
rlabel locali s 298695 67725 298799 67833 6 VGND
port 614 nsew ground input
rlabel locali s 1121 67725 1225 67833 6 VGND
port 614 nsew ground input
rlabel locali s 298660 67833 298799 67983 6 VGND
port 614 nsew ground input
rlabel locali s 298660 67983 298816 68017 6 VGND
port 614 nsew ground input
rlabel locali s 298660 68017 298799 68167 6 VGND
port 614 nsew ground input
rlabel locali s 1121 67833 1340 67983 6 VGND
port 614 nsew ground input
rlabel locali s 1104 67983 1340 68017 6 VGND
port 614 nsew ground input
rlabel locali s 1121 68017 1340 68167 6 VGND
port 614 nsew ground input
rlabel locali s 298695 68167 298799 68275 6 VGND
port 614 nsew ground input
rlabel locali s 1121 68167 1225 68275 6 VGND
port 614 nsew ground input
rlabel locali s 298695 68813 298799 68921 6 VGND
port 614 nsew ground input
rlabel locali s 1121 68813 1225 68921 6 VGND
port 614 nsew ground input
rlabel locali s 298660 68921 298799 69071 6 VGND
port 614 nsew ground input
rlabel locali s 298660 69071 298816 69105 6 VGND
port 614 nsew ground input
rlabel locali s 298660 69105 298799 69255 6 VGND
port 614 nsew ground input
rlabel locali s 1121 68921 1340 69071 6 VGND
port 614 nsew ground input
rlabel locali s 1104 69071 1340 69105 6 VGND
port 614 nsew ground input
rlabel locali s 1121 69105 1340 69255 6 VGND
port 614 nsew ground input
rlabel locali s 298695 69255 298799 69363 6 VGND
port 614 nsew ground input
rlabel locali s 1121 69255 1225 69363 6 VGND
port 614 nsew ground input
rlabel locali s 298695 69901 298799 70009 6 VGND
port 614 nsew ground input
rlabel locali s 1121 69901 1225 70009 6 VGND
port 614 nsew ground input
rlabel locali s 298660 70009 298799 70159 6 VGND
port 614 nsew ground input
rlabel locali s 298660 70159 298816 70193 6 VGND
port 614 nsew ground input
rlabel locali s 298660 70193 298799 70343 6 VGND
port 614 nsew ground input
rlabel locali s 1121 70009 1340 70159 6 VGND
port 614 nsew ground input
rlabel locali s 1104 70159 1340 70193 6 VGND
port 614 nsew ground input
rlabel locali s 1121 70193 1340 70343 6 VGND
port 614 nsew ground input
rlabel locali s 298695 70343 298799 70451 6 VGND
port 614 nsew ground input
rlabel locali s 1121 70343 1225 70451 6 VGND
port 614 nsew ground input
rlabel locali s 298695 70989 298799 71097 6 VGND
port 614 nsew ground input
rlabel locali s 1121 70989 1225 71097 6 VGND
port 614 nsew ground input
rlabel locali s 298660 71097 298799 71247 6 VGND
port 614 nsew ground input
rlabel locali s 298660 71247 298816 71281 6 VGND
port 614 nsew ground input
rlabel locali s 298660 71281 298799 71431 6 VGND
port 614 nsew ground input
rlabel locali s 1121 71097 1340 71247 6 VGND
port 614 nsew ground input
rlabel locali s 1104 71247 1340 71281 6 VGND
port 614 nsew ground input
rlabel locali s 1121 71281 1340 71431 6 VGND
port 614 nsew ground input
rlabel locali s 298695 71431 298799 71539 6 VGND
port 614 nsew ground input
rlabel locali s 1121 71431 1225 71539 6 VGND
port 614 nsew ground input
rlabel locali s 298695 72077 298799 72185 6 VGND
port 614 nsew ground input
rlabel locali s 1121 72077 1225 72185 6 VGND
port 614 nsew ground input
rlabel locali s 298660 72185 298799 72335 6 VGND
port 614 nsew ground input
rlabel locali s 298660 72335 298816 72369 6 VGND
port 614 nsew ground input
rlabel locali s 298660 72369 298799 72519 6 VGND
port 614 nsew ground input
rlabel locali s 1121 72185 1340 72335 6 VGND
port 614 nsew ground input
rlabel locali s 1104 72335 1340 72369 6 VGND
port 614 nsew ground input
rlabel locali s 1121 72369 1340 72519 6 VGND
port 614 nsew ground input
rlabel locali s 298695 72519 298799 72627 6 VGND
port 614 nsew ground input
rlabel locali s 1121 72519 1225 72627 6 VGND
port 614 nsew ground input
rlabel locali s 298695 73165 298799 73273 6 VGND
port 614 nsew ground input
rlabel locali s 1121 73165 1225 73273 6 VGND
port 614 nsew ground input
rlabel locali s 298660 73273 298799 73423 6 VGND
port 614 nsew ground input
rlabel locali s 298660 73423 298816 73457 6 VGND
port 614 nsew ground input
rlabel locali s 298660 73457 298799 73607 6 VGND
port 614 nsew ground input
rlabel locali s 1121 73273 1340 73423 6 VGND
port 614 nsew ground input
rlabel locali s 1104 73423 1340 73457 6 VGND
port 614 nsew ground input
rlabel locali s 1121 73457 1340 73607 6 VGND
port 614 nsew ground input
rlabel locali s 298695 73607 298799 73715 6 VGND
port 614 nsew ground input
rlabel locali s 1121 73607 1225 73715 6 VGND
port 614 nsew ground input
rlabel locali s 298695 74253 298799 74361 6 VGND
port 614 nsew ground input
rlabel locali s 1121 74253 1225 74361 6 VGND
port 614 nsew ground input
rlabel locali s 298660 74361 298799 74511 6 VGND
port 614 nsew ground input
rlabel locali s 298660 74511 298816 74545 6 VGND
port 614 nsew ground input
rlabel locali s 298660 74545 298799 74695 6 VGND
port 614 nsew ground input
rlabel locali s 1121 74361 1340 74511 6 VGND
port 614 nsew ground input
rlabel locali s 1104 74511 1340 74545 6 VGND
port 614 nsew ground input
rlabel locali s 1121 74545 1340 74695 6 VGND
port 614 nsew ground input
rlabel locali s 298695 74695 298799 74803 6 VGND
port 614 nsew ground input
rlabel locali s 1121 74695 1225 74803 6 VGND
port 614 nsew ground input
rlabel locali s 298695 75341 298799 75449 6 VGND
port 614 nsew ground input
rlabel locali s 1121 75341 1225 75449 6 VGND
port 614 nsew ground input
rlabel locali s 298660 75449 298799 75599 6 VGND
port 614 nsew ground input
rlabel locali s 298660 75599 298816 75633 6 VGND
port 614 nsew ground input
rlabel locali s 298660 75633 298799 75783 6 VGND
port 614 nsew ground input
rlabel locali s 1121 75449 1340 75599 6 VGND
port 614 nsew ground input
rlabel locali s 1104 75599 1340 75633 6 VGND
port 614 nsew ground input
rlabel locali s 1121 75633 1340 75783 6 VGND
port 614 nsew ground input
rlabel locali s 298695 75783 298799 75891 6 VGND
port 614 nsew ground input
rlabel locali s 1121 75783 1225 75891 6 VGND
port 614 nsew ground input
rlabel locali s 298695 76429 298799 76537 6 VGND
port 614 nsew ground input
rlabel locali s 1121 76429 1225 76537 6 VGND
port 614 nsew ground input
rlabel locali s 298660 76537 298799 76687 6 VGND
port 614 nsew ground input
rlabel locali s 298660 76687 298816 76721 6 VGND
port 614 nsew ground input
rlabel locali s 298660 76721 298799 76871 6 VGND
port 614 nsew ground input
rlabel locali s 1121 76537 1340 76687 6 VGND
port 614 nsew ground input
rlabel locali s 1104 76687 1340 76721 6 VGND
port 614 nsew ground input
rlabel locali s 1121 76721 1340 76871 6 VGND
port 614 nsew ground input
rlabel locali s 298695 76871 298799 76979 6 VGND
port 614 nsew ground input
rlabel locali s 1121 76871 1225 76979 6 VGND
port 614 nsew ground input
rlabel locali s 298695 77517 298799 77625 6 VGND
port 614 nsew ground input
rlabel locali s 1121 77517 1225 77625 6 VGND
port 614 nsew ground input
rlabel locali s 298660 77625 298799 77775 6 VGND
port 614 nsew ground input
rlabel locali s 298660 77775 298816 77809 6 VGND
port 614 nsew ground input
rlabel locali s 298660 77809 298799 77959 6 VGND
port 614 nsew ground input
rlabel locali s 1121 77625 1340 77775 6 VGND
port 614 nsew ground input
rlabel locali s 1104 77775 1340 77809 6 VGND
port 614 nsew ground input
rlabel locali s 1121 77809 1340 77959 6 VGND
port 614 nsew ground input
rlabel locali s 298695 77959 298799 78067 6 VGND
port 614 nsew ground input
rlabel locali s 1121 77959 1225 78067 6 VGND
port 614 nsew ground input
rlabel locali s 298695 78605 298799 78713 6 VGND
port 614 nsew ground input
rlabel locali s 1121 78605 1225 78713 6 VGND
port 614 nsew ground input
rlabel locali s 298660 78713 298799 78863 6 VGND
port 614 nsew ground input
rlabel locali s 298660 78863 298816 78897 6 VGND
port 614 nsew ground input
rlabel locali s 298660 78897 298799 79047 6 VGND
port 614 nsew ground input
rlabel locali s 1121 78713 1340 78863 6 VGND
port 614 nsew ground input
rlabel locali s 1104 78863 1340 78897 6 VGND
port 614 nsew ground input
rlabel locali s 1121 78897 1340 79047 6 VGND
port 614 nsew ground input
rlabel locali s 298695 79047 298799 79155 6 VGND
port 614 nsew ground input
rlabel locali s 1121 79047 1225 79155 6 VGND
port 614 nsew ground input
rlabel locali s 298695 79693 298799 79801 6 VGND
port 614 nsew ground input
rlabel locali s 1121 79693 1225 79801 6 VGND
port 614 nsew ground input
rlabel locali s 298660 79801 298799 79951 6 VGND
port 614 nsew ground input
rlabel locali s 298660 79951 298816 79985 6 VGND
port 614 nsew ground input
rlabel locali s 298660 79985 298799 80135 6 VGND
port 614 nsew ground input
rlabel locali s 1121 79801 1340 79951 6 VGND
port 614 nsew ground input
rlabel locali s 1104 79951 1340 79985 6 VGND
port 614 nsew ground input
rlabel locali s 1121 79985 1340 80135 6 VGND
port 614 nsew ground input
rlabel locali s 298695 80135 298799 80243 6 VGND
port 614 nsew ground input
rlabel locali s 1121 80135 1225 80243 6 VGND
port 614 nsew ground input
rlabel locali s 298695 80781 298799 80889 6 VGND
port 614 nsew ground input
rlabel locali s 1121 80781 1225 80889 6 VGND
port 614 nsew ground input
rlabel locali s 298660 80889 298799 81039 6 VGND
port 614 nsew ground input
rlabel locali s 298660 81039 298816 81073 6 VGND
port 614 nsew ground input
rlabel locali s 298660 81073 298799 81223 6 VGND
port 614 nsew ground input
rlabel locali s 1121 80889 1340 81039 6 VGND
port 614 nsew ground input
rlabel locali s 1104 81039 1340 81073 6 VGND
port 614 nsew ground input
rlabel locali s 1121 81073 1340 81223 6 VGND
port 614 nsew ground input
rlabel locali s 298695 81223 298799 81331 6 VGND
port 614 nsew ground input
rlabel locali s 1121 81223 1225 81331 6 VGND
port 614 nsew ground input
rlabel locali s 298695 81869 298799 81977 6 VGND
port 614 nsew ground input
rlabel locali s 1121 81869 1225 81977 6 VGND
port 614 nsew ground input
rlabel locali s 298660 81977 298799 82127 6 VGND
port 614 nsew ground input
rlabel locali s 298660 82127 298816 82161 6 VGND
port 614 nsew ground input
rlabel locali s 298660 82161 298799 82311 6 VGND
port 614 nsew ground input
rlabel locali s 1121 81977 1340 82127 6 VGND
port 614 nsew ground input
rlabel locali s 1104 82127 1340 82161 6 VGND
port 614 nsew ground input
rlabel locali s 1121 82161 1340 82311 6 VGND
port 614 nsew ground input
rlabel locali s 298695 82311 298799 82419 6 VGND
port 614 nsew ground input
rlabel locali s 1121 82311 1225 82419 6 VGND
port 614 nsew ground input
rlabel locali s 298695 82957 298799 83065 6 VGND
port 614 nsew ground input
rlabel locali s 1121 82957 1225 83065 6 VGND
port 614 nsew ground input
rlabel locali s 298660 83065 298799 83215 6 VGND
port 614 nsew ground input
rlabel locali s 298660 83215 298816 83249 6 VGND
port 614 nsew ground input
rlabel locali s 298660 83249 298799 83399 6 VGND
port 614 nsew ground input
rlabel locali s 1121 83065 1340 83215 6 VGND
port 614 nsew ground input
rlabel locali s 1104 83215 1340 83249 6 VGND
port 614 nsew ground input
rlabel locali s 1121 83249 1340 83399 6 VGND
port 614 nsew ground input
rlabel locali s 298695 83399 298799 83507 6 VGND
port 614 nsew ground input
rlabel locali s 1121 83399 1225 83507 6 VGND
port 614 nsew ground input
rlabel locali s 298695 84045 298799 84153 6 VGND
port 614 nsew ground input
rlabel locali s 1121 84045 1225 84153 6 VGND
port 614 nsew ground input
rlabel locali s 298660 84153 298799 84303 6 VGND
port 614 nsew ground input
rlabel locali s 298660 84303 298816 84337 6 VGND
port 614 nsew ground input
rlabel locali s 298660 84337 298799 84487 6 VGND
port 614 nsew ground input
rlabel locali s 1121 84153 1340 84303 6 VGND
port 614 nsew ground input
rlabel locali s 1104 84303 1340 84337 6 VGND
port 614 nsew ground input
rlabel locali s 1121 84337 1340 84487 6 VGND
port 614 nsew ground input
rlabel locali s 298695 84487 298799 84595 6 VGND
port 614 nsew ground input
rlabel locali s 1121 84487 1225 84595 6 VGND
port 614 nsew ground input
rlabel locali s 298695 85133 298799 85241 6 VGND
port 614 nsew ground input
rlabel locali s 1121 85133 1225 85241 6 VGND
port 614 nsew ground input
rlabel locali s 298660 85241 298799 85391 6 VGND
port 614 nsew ground input
rlabel locali s 298660 85391 298816 85425 6 VGND
port 614 nsew ground input
rlabel locali s 298660 85425 298799 85575 6 VGND
port 614 nsew ground input
rlabel locali s 1121 85241 1340 85391 6 VGND
port 614 nsew ground input
rlabel locali s 1104 85391 1340 85425 6 VGND
port 614 nsew ground input
rlabel locali s 1121 85425 1340 85575 6 VGND
port 614 nsew ground input
rlabel locali s 298695 85575 298799 85683 6 VGND
port 614 nsew ground input
rlabel locali s 1121 85575 1225 85683 6 VGND
port 614 nsew ground input
rlabel locali s 298695 86221 298799 86329 6 VGND
port 614 nsew ground input
rlabel locali s 1121 86221 1225 86329 6 VGND
port 614 nsew ground input
rlabel locali s 298660 86329 298799 86479 6 VGND
port 614 nsew ground input
rlabel locali s 298660 86479 298816 86513 6 VGND
port 614 nsew ground input
rlabel locali s 298660 86513 298799 86663 6 VGND
port 614 nsew ground input
rlabel locali s 1121 86329 1340 86479 6 VGND
port 614 nsew ground input
rlabel locali s 1104 86479 1340 86513 6 VGND
port 614 nsew ground input
rlabel locali s 1121 86513 1340 86663 6 VGND
port 614 nsew ground input
rlabel locali s 298695 86663 298799 86771 6 VGND
port 614 nsew ground input
rlabel locali s 1121 86663 1225 86771 6 VGND
port 614 nsew ground input
rlabel locali s 298695 87309 298799 87417 6 VGND
port 614 nsew ground input
rlabel locali s 1121 87309 1225 87417 6 VGND
port 614 nsew ground input
rlabel locali s 298660 87417 298799 87567 6 VGND
port 614 nsew ground input
rlabel locali s 298660 87567 298816 87601 6 VGND
port 614 nsew ground input
rlabel locali s 298660 87601 298799 87751 6 VGND
port 614 nsew ground input
rlabel locali s 1121 87417 1340 87567 6 VGND
port 614 nsew ground input
rlabel locali s 1104 87567 1340 87601 6 VGND
port 614 nsew ground input
rlabel locali s 1121 87601 1340 87751 6 VGND
port 614 nsew ground input
rlabel locali s 298695 87751 298799 87859 6 VGND
port 614 nsew ground input
rlabel locali s 1121 87751 1225 87859 6 VGND
port 614 nsew ground input
rlabel locali s 298695 88397 298799 88505 6 VGND
port 614 nsew ground input
rlabel locali s 1121 88397 1225 88505 6 VGND
port 614 nsew ground input
rlabel locali s 298660 88505 298799 88655 6 VGND
port 614 nsew ground input
rlabel locali s 298660 88655 298816 88689 6 VGND
port 614 nsew ground input
rlabel locali s 298660 88689 298799 88839 6 VGND
port 614 nsew ground input
rlabel locali s 1121 88505 1340 88655 6 VGND
port 614 nsew ground input
rlabel locali s 1104 88655 1340 88689 6 VGND
port 614 nsew ground input
rlabel locali s 1121 88689 1340 88839 6 VGND
port 614 nsew ground input
rlabel locali s 298695 88839 298799 88947 6 VGND
port 614 nsew ground input
rlabel locali s 1121 88839 1225 88947 6 VGND
port 614 nsew ground input
rlabel locali s 298695 89485 298799 89593 6 VGND
port 614 nsew ground input
rlabel locali s 1121 89485 1225 89593 6 VGND
port 614 nsew ground input
rlabel locali s 298660 89593 298799 89743 6 VGND
port 614 nsew ground input
rlabel locali s 298660 89743 298816 89777 6 VGND
port 614 nsew ground input
rlabel locali s 298660 89777 298799 89927 6 VGND
port 614 nsew ground input
rlabel locali s 1121 89593 1340 89743 6 VGND
port 614 nsew ground input
rlabel locali s 1104 89743 1340 89777 6 VGND
port 614 nsew ground input
rlabel locali s 1121 89777 1340 89927 6 VGND
port 614 nsew ground input
rlabel locali s 298695 89927 298799 90035 6 VGND
port 614 nsew ground input
rlabel locali s 1121 89927 1225 90035 6 VGND
port 614 nsew ground input
rlabel locali s 298695 90573 298799 90681 6 VGND
port 614 nsew ground input
rlabel locali s 1121 90573 1225 90681 6 VGND
port 614 nsew ground input
rlabel locali s 298660 90681 298799 90831 6 VGND
port 614 nsew ground input
rlabel locali s 298660 90831 298816 90865 6 VGND
port 614 nsew ground input
rlabel locali s 298660 90865 298799 91015 6 VGND
port 614 nsew ground input
rlabel locali s 1121 90681 1340 90831 6 VGND
port 614 nsew ground input
rlabel locali s 1104 90831 1340 90865 6 VGND
port 614 nsew ground input
rlabel locali s 1121 90865 1340 91015 6 VGND
port 614 nsew ground input
rlabel locali s 298695 91015 298799 91123 6 VGND
port 614 nsew ground input
rlabel locali s 1121 91015 1225 91123 6 VGND
port 614 nsew ground input
rlabel locali s 298695 91661 298799 91769 6 VGND
port 614 nsew ground input
rlabel locali s 1121 91661 1225 91769 6 VGND
port 614 nsew ground input
rlabel locali s 298660 91769 298799 91919 6 VGND
port 614 nsew ground input
rlabel locali s 298660 91919 298816 91953 6 VGND
port 614 nsew ground input
rlabel locali s 298660 91953 298799 92103 6 VGND
port 614 nsew ground input
rlabel locali s 1121 91769 1340 91919 6 VGND
port 614 nsew ground input
rlabel locali s 1104 91919 1340 91953 6 VGND
port 614 nsew ground input
rlabel locali s 1121 91953 1340 92103 6 VGND
port 614 nsew ground input
rlabel locali s 298695 92103 298799 92211 6 VGND
port 614 nsew ground input
rlabel locali s 1121 92103 1225 92211 6 VGND
port 614 nsew ground input
rlabel locali s 298695 92749 298799 92857 6 VGND
port 614 nsew ground input
rlabel locali s 1121 92749 1225 92857 6 VGND
port 614 nsew ground input
rlabel locali s 298660 92857 298799 93007 6 VGND
port 614 nsew ground input
rlabel locali s 298660 93007 298816 93041 6 VGND
port 614 nsew ground input
rlabel locali s 298660 93041 298799 93191 6 VGND
port 614 nsew ground input
rlabel locali s 1121 92857 1340 93007 6 VGND
port 614 nsew ground input
rlabel locali s 1104 93007 1340 93041 6 VGND
port 614 nsew ground input
rlabel locali s 1121 93041 1340 93191 6 VGND
port 614 nsew ground input
rlabel locali s 298695 93191 298799 93299 6 VGND
port 614 nsew ground input
rlabel locali s 1121 93191 1225 93299 6 VGND
port 614 nsew ground input
rlabel locali s 298695 93837 298799 93945 6 VGND
port 614 nsew ground input
rlabel locali s 1121 93837 1225 93945 6 VGND
port 614 nsew ground input
rlabel locali s 298660 93945 298799 94095 6 VGND
port 614 nsew ground input
rlabel locali s 298660 94095 298816 94129 6 VGND
port 614 nsew ground input
rlabel locali s 298660 94129 298799 94279 6 VGND
port 614 nsew ground input
rlabel locali s 1121 93945 1340 94095 6 VGND
port 614 nsew ground input
rlabel locali s 1104 94095 1340 94129 6 VGND
port 614 nsew ground input
rlabel locali s 1121 94129 1340 94279 6 VGND
port 614 nsew ground input
rlabel locali s 298695 94279 298799 94387 6 VGND
port 614 nsew ground input
rlabel locali s 1121 94279 1225 94387 6 VGND
port 614 nsew ground input
rlabel locali s 298695 94925 298799 95033 6 VGND
port 614 nsew ground input
rlabel locali s 1121 94925 1225 95033 6 VGND
port 614 nsew ground input
rlabel locali s 298660 95033 298799 95183 6 VGND
port 614 nsew ground input
rlabel locali s 298660 95183 298816 95217 6 VGND
port 614 nsew ground input
rlabel locali s 298660 95217 298799 95367 6 VGND
port 614 nsew ground input
rlabel locali s 1121 95033 1340 95183 6 VGND
port 614 nsew ground input
rlabel locali s 1104 95183 1340 95217 6 VGND
port 614 nsew ground input
rlabel locali s 1121 95217 1340 95367 6 VGND
port 614 nsew ground input
rlabel locali s 298695 95367 298799 95475 6 VGND
port 614 nsew ground input
rlabel locali s 1121 95367 1225 95475 6 VGND
port 614 nsew ground input
rlabel locali s 298695 96013 298799 96121 6 VGND
port 614 nsew ground input
rlabel locali s 1121 96013 1225 96121 6 VGND
port 614 nsew ground input
rlabel locali s 298660 96121 298799 96271 6 VGND
port 614 nsew ground input
rlabel locali s 298660 96271 298816 96305 6 VGND
port 614 nsew ground input
rlabel locali s 298660 96305 298799 96455 6 VGND
port 614 nsew ground input
rlabel locali s 1121 96121 1340 96271 6 VGND
port 614 nsew ground input
rlabel locali s 1104 96271 1340 96305 6 VGND
port 614 nsew ground input
rlabel locali s 1121 96305 1340 96455 6 VGND
port 614 nsew ground input
rlabel locali s 298695 96455 298799 96563 6 VGND
port 614 nsew ground input
rlabel locali s 1121 96455 1225 96563 6 VGND
port 614 nsew ground input
rlabel locali s 298695 97101 298799 97209 6 VGND
port 614 nsew ground input
rlabel locali s 1121 97101 1225 97209 6 VGND
port 614 nsew ground input
rlabel locali s 298660 97209 298799 97359 6 VGND
port 614 nsew ground input
rlabel locali s 298660 97359 298816 97393 6 VGND
port 614 nsew ground input
rlabel locali s 298660 97393 298799 97543 6 VGND
port 614 nsew ground input
rlabel locali s 1121 97209 1340 97359 6 VGND
port 614 nsew ground input
rlabel locali s 1104 97359 1340 97393 6 VGND
port 614 nsew ground input
rlabel locali s 1121 97393 1340 97543 6 VGND
port 614 nsew ground input
rlabel locali s 298695 97543 298799 97651 6 VGND
port 614 nsew ground input
rlabel locali s 1121 97543 1225 97651 6 VGND
port 614 nsew ground input
rlabel locali s 298695 98189 298799 98297 6 VGND
port 614 nsew ground input
rlabel locali s 1121 98189 1225 98297 6 VGND
port 614 nsew ground input
rlabel locali s 298660 98297 298799 98447 6 VGND
port 614 nsew ground input
rlabel locali s 298660 98447 298816 98481 6 VGND
port 614 nsew ground input
rlabel locali s 298660 98481 298799 98631 6 VGND
port 614 nsew ground input
rlabel locali s 1121 98297 1340 98447 6 VGND
port 614 nsew ground input
rlabel locali s 1104 98447 1340 98481 6 VGND
port 614 nsew ground input
rlabel locali s 1121 98481 1340 98631 6 VGND
port 614 nsew ground input
rlabel locali s 298695 98631 298799 98739 6 VGND
port 614 nsew ground input
rlabel locali s 1121 98631 1225 98739 6 VGND
port 614 nsew ground input
rlabel locali s 298695 99277 298799 99385 6 VGND
port 614 nsew ground input
rlabel locali s 1121 99277 1225 99385 6 VGND
port 614 nsew ground input
rlabel locali s 298660 99385 298799 99535 6 VGND
port 614 nsew ground input
rlabel locali s 298660 99535 298816 99569 6 VGND
port 614 nsew ground input
rlabel locali s 298660 99569 298799 99719 6 VGND
port 614 nsew ground input
rlabel locali s 1121 99385 1340 99535 6 VGND
port 614 nsew ground input
rlabel locali s 1104 99535 1340 99569 6 VGND
port 614 nsew ground input
rlabel locali s 1121 99569 1340 99719 6 VGND
port 614 nsew ground input
rlabel locali s 298695 99719 298799 99827 6 VGND
port 614 nsew ground input
rlabel locali s 1121 99719 1225 99827 6 VGND
port 614 nsew ground input
rlabel locali s 298695 100365 298799 100473 6 VGND
port 614 nsew ground input
rlabel locali s 1121 100365 1225 100473 6 VGND
port 614 nsew ground input
rlabel locali s 298660 100473 298799 100623 6 VGND
port 614 nsew ground input
rlabel locali s 298660 100623 298816 100657 6 VGND
port 614 nsew ground input
rlabel locali s 298660 100657 298799 100807 6 VGND
port 614 nsew ground input
rlabel locali s 1121 100473 1340 100623 6 VGND
port 614 nsew ground input
rlabel locali s 1104 100623 1340 100657 6 VGND
port 614 nsew ground input
rlabel locali s 1121 100657 1340 100807 6 VGND
port 614 nsew ground input
rlabel locali s 298695 100807 298799 100915 6 VGND
port 614 nsew ground input
rlabel locali s 1121 100807 1225 100915 6 VGND
port 614 nsew ground input
rlabel locali s 298695 101453 298799 101561 6 VGND
port 614 nsew ground input
rlabel locali s 1121 101453 1225 101561 6 VGND
port 614 nsew ground input
rlabel locali s 298660 101561 298799 101711 6 VGND
port 614 nsew ground input
rlabel locali s 298660 101711 298816 101745 6 VGND
port 614 nsew ground input
rlabel locali s 298660 101745 298799 101895 6 VGND
port 614 nsew ground input
rlabel locali s 1121 101561 1340 101711 6 VGND
port 614 nsew ground input
rlabel locali s 1104 101711 1340 101745 6 VGND
port 614 nsew ground input
rlabel locali s 1121 101745 1340 101895 6 VGND
port 614 nsew ground input
rlabel locali s 298695 101895 298799 102003 6 VGND
port 614 nsew ground input
rlabel locali s 1121 101895 1225 102003 6 VGND
port 614 nsew ground input
rlabel locali s 298695 102541 298799 102649 6 VGND
port 614 nsew ground input
rlabel locali s 1121 102541 1225 102649 6 VGND
port 614 nsew ground input
rlabel locali s 298660 102649 298799 102799 6 VGND
port 614 nsew ground input
rlabel locali s 298660 102799 298816 102833 6 VGND
port 614 nsew ground input
rlabel locali s 298660 102833 298799 102983 6 VGND
port 614 nsew ground input
rlabel locali s 1121 102649 1340 102799 6 VGND
port 614 nsew ground input
rlabel locali s 1104 102799 1340 102833 6 VGND
port 614 nsew ground input
rlabel locali s 1121 102833 1340 102983 6 VGND
port 614 nsew ground input
rlabel locali s 298695 102983 298799 103091 6 VGND
port 614 nsew ground input
rlabel locali s 1121 102983 1225 103091 6 VGND
port 614 nsew ground input
rlabel locali s 298695 103629 298799 103737 6 VGND
port 614 nsew ground input
rlabel locali s 1121 103629 1225 103737 6 VGND
port 614 nsew ground input
rlabel locali s 298660 103737 298799 103887 6 VGND
port 614 nsew ground input
rlabel locali s 298660 103887 298816 103921 6 VGND
port 614 nsew ground input
rlabel locali s 298660 103921 298799 104071 6 VGND
port 614 nsew ground input
rlabel locali s 1121 103737 1340 103887 6 VGND
port 614 nsew ground input
rlabel locali s 1104 103887 1340 103921 6 VGND
port 614 nsew ground input
rlabel locali s 1121 103921 1340 104071 6 VGND
port 614 nsew ground input
rlabel locali s 298695 104071 298799 104179 6 VGND
port 614 nsew ground input
rlabel locali s 1121 104071 1225 104179 6 VGND
port 614 nsew ground input
rlabel locali s 298695 104717 298799 104825 6 VGND
port 614 nsew ground input
rlabel locali s 1121 104717 1225 104825 6 VGND
port 614 nsew ground input
rlabel locali s 298660 104825 298799 104975 6 VGND
port 614 nsew ground input
rlabel locali s 298660 104975 298816 105009 6 VGND
port 614 nsew ground input
rlabel locali s 298660 105009 298799 105159 6 VGND
port 614 nsew ground input
rlabel locali s 1121 104825 1340 104975 6 VGND
port 614 nsew ground input
rlabel locali s 1104 104975 1340 105009 6 VGND
port 614 nsew ground input
rlabel locali s 1121 105009 1340 105159 6 VGND
port 614 nsew ground input
rlabel locali s 298695 105159 298799 105267 6 VGND
port 614 nsew ground input
rlabel locali s 1121 105159 1225 105267 6 VGND
port 614 nsew ground input
rlabel locali s 298695 105805 298799 105913 6 VGND
port 614 nsew ground input
rlabel locali s 1121 105805 1225 105913 6 VGND
port 614 nsew ground input
rlabel locali s 298660 105913 298799 106063 6 VGND
port 614 nsew ground input
rlabel locali s 298660 106063 298816 106097 6 VGND
port 614 nsew ground input
rlabel locali s 298660 106097 298799 106247 6 VGND
port 614 nsew ground input
rlabel locali s 1121 105913 1340 106063 6 VGND
port 614 nsew ground input
rlabel locali s 1104 106063 1340 106097 6 VGND
port 614 nsew ground input
rlabel locali s 1121 106097 1340 106247 6 VGND
port 614 nsew ground input
rlabel locali s 298695 106247 298799 106355 6 VGND
port 614 nsew ground input
rlabel locali s 1121 106247 1225 106355 6 VGND
port 614 nsew ground input
rlabel locali s 298695 106893 298799 107001 6 VGND
port 614 nsew ground input
rlabel locali s 1121 106893 1225 107001 6 VGND
port 614 nsew ground input
rlabel locali s 298660 107001 298799 107151 6 VGND
port 614 nsew ground input
rlabel locali s 298660 107151 298816 107185 6 VGND
port 614 nsew ground input
rlabel locali s 298660 107185 298799 107335 6 VGND
port 614 nsew ground input
rlabel locali s 1121 107001 1340 107151 6 VGND
port 614 nsew ground input
rlabel locali s 1104 107151 1340 107185 6 VGND
port 614 nsew ground input
rlabel locali s 1121 107185 1340 107335 6 VGND
port 614 nsew ground input
rlabel locali s 298695 107335 298799 107443 6 VGND
port 614 nsew ground input
rlabel locali s 1121 107335 1225 107443 6 VGND
port 614 nsew ground input
rlabel locali s 298695 107981 298799 108089 6 VGND
port 614 nsew ground input
rlabel locali s 1121 107981 1225 108089 6 VGND
port 614 nsew ground input
rlabel locali s 298660 108089 298799 108239 6 VGND
port 614 nsew ground input
rlabel locali s 298660 108239 298816 108273 6 VGND
port 614 nsew ground input
rlabel locali s 298660 108273 298799 108423 6 VGND
port 614 nsew ground input
rlabel locali s 1121 108089 1340 108239 6 VGND
port 614 nsew ground input
rlabel locali s 1104 108239 1340 108273 6 VGND
port 614 nsew ground input
rlabel locali s 1121 108273 1340 108423 6 VGND
port 614 nsew ground input
rlabel locali s 298695 108423 298799 108531 6 VGND
port 614 nsew ground input
rlabel locali s 1121 108423 1225 108531 6 VGND
port 614 nsew ground input
rlabel locali s 298695 109069 298799 109177 6 VGND
port 614 nsew ground input
rlabel locali s 1121 109069 1225 109177 6 VGND
port 614 nsew ground input
rlabel locali s 298660 109177 298799 109327 6 VGND
port 614 nsew ground input
rlabel locali s 298660 109327 298816 109361 6 VGND
port 614 nsew ground input
rlabel locali s 298660 109361 298799 109511 6 VGND
port 614 nsew ground input
rlabel locali s 1121 109177 1340 109327 6 VGND
port 614 nsew ground input
rlabel locali s 1104 109327 1340 109361 6 VGND
port 614 nsew ground input
rlabel locali s 1121 109361 1340 109511 6 VGND
port 614 nsew ground input
rlabel locali s 298695 109511 298799 109619 6 VGND
port 614 nsew ground input
rlabel locali s 1121 109511 1225 109619 6 VGND
port 614 nsew ground input
rlabel locali s 298695 110157 298799 110265 6 VGND
port 614 nsew ground input
rlabel locali s 1121 110157 1225 110265 6 VGND
port 614 nsew ground input
rlabel locali s 298660 110265 298799 110415 6 VGND
port 614 nsew ground input
rlabel locali s 298660 110415 298816 110449 6 VGND
port 614 nsew ground input
rlabel locali s 298660 110449 298799 110599 6 VGND
port 614 nsew ground input
rlabel locali s 1121 110265 1340 110415 6 VGND
port 614 nsew ground input
rlabel locali s 1104 110415 1340 110449 6 VGND
port 614 nsew ground input
rlabel locali s 1121 110449 1340 110599 6 VGND
port 614 nsew ground input
rlabel locali s 298695 110599 298799 110707 6 VGND
port 614 nsew ground input
rlabel locali s 1121 110599 1225 110707 6 VGND
port 614 nsew ground input
rlabel locali s 298695 111245 298799 111353 6 VGND
port 614 nsew ground input
rlabel locali s 1121 111245 1225 111353 6 VGND
port 614 nsew ground input
rlabel locali s 298660 111353 298799 111503 6 VGND
port 614 nsew ground input
rlabel locali s 298660 111503 298816 111537 6 VGND
port 614 nsew ground input
rlabel locali s 298660 111537 298799 111687 6 VGND
port 614 nsew ground input
rlabel locali s 1121 111353 1340 111503 6 VGND
port 614 nsew ground input
rlabel locali s 1104 111503 1340 111537 6 VGND
port 614 nsew ground input
rlabel locali s 1121 111537 1340 111687 6 VGND
port 614 nsew ground input
rlabel locali s 298695 111687 298799 111795 6 VGND
port 614 nsew ground input
rlabel locali s 1121 111687 1225 111795 6 VGND
port 614 nsew ground input
rlabel locali s 298695 112333 298799 112441 6 VGND
port 614 nsew ground input
rlabel locali s 1121 112333 1225 112441 6 VGND
port 614 nsew ground input
rlabel locali s 298660 112441 298799 112591 6 VGND
port 614 nsew ground input
rlabel locali s 298660 112591 298816 112625 6 VGND
port 614 nsew ground input
rlabel locali s 298660 112625 298799 112775 6 VGND
port 614 nsew ground input
rlabel locali s 1121 112441 1340 112591 6 VGND
port 614 nsew ground input
rlabel locali s 1104 112591 1340 112625 6 VGND
port 614 nsew ground input
rlabel locali s 1121 112625 1340 112775 6 VGND
port 614 nsew ground input
rlabel locali s 298695 112775 298799 112883 6 VGND
port 614 nsew ground input
rlabel locali s 1121 112775 1225 112883 6 VGND
port 614 nsew ground input
rlabel locali s 298695 113421 298799 113529 6 VGND
port 614 nsew ground input
rlabel locali s 1121 113421 1225 113529 6 VGND
port 614 nsew ground input
rlabel locali s 298660 113529 298799 113679 6 VGND
port 614 nsew ground input
rlabel locali s 298660 113679 298816 113713 6 VGND
port 614 nsew ground input
rlabel locali s 298660 113713 298799 113863 6 VGND
port 614 nsew ground input
rlabel locali s 1121 113529 1340 113679 6 VGND
port 614 nsew ground input
rlabel locali s 1104 113679 1340 113713 6 VGND
port 614 nsew ground input
rlabel locali s 1121 113713 1340 113863 6 VGND
port 614 nsew ground input
rlabel locali s 298695 113863 298799 113971 6 VGND
port 614 nsew ground input
rlabel locali s 1121 113863 1225 113971 6 VGND
port 614 nsew ground input
rlabel locali s 298695 114509 298799 114617 6 VGND
port 614 nsew ground input
rlabel locali s 1121 114509 1225 114617 6 VGND
port 614 nsew ground input
rlabel locali s 298660 114617 298799 114767 6 VGND
port 614 nsew ground input
rlabel locali s 298660 114767 298816 114801 6 VGND
port 614 nsew ground input
rlabel locali s 298660 114801 298799 114951 6 VGND
port 614 nsew ground input
rlabel locali s 1121 114617 1340 114767 6 VGND
port 614 nsew ground input
rlabel locali s 1104 114767 1340 114801 6 VGND
port 614 nsew ground input
rlabel locali s 1121 114801 1340 114951 6 VGND
port 614 nsew ground input
rlabel locali s 298695 114951 298799 115059 6 VGND
port 614 nsew ground input
rlabel locali s 1121 114951 1225 115059 6 VGND
port 614 nsew ground input
rlabel locali s 298695 115597 298799 115705 6 VGND
port 614 nsew ground input
rlabel locali s 1121 115597 1225 115705 6 VGND
port 614 nsew ground input
rlabel locali s 298660 115705 298799 115855 6 VGND
port 614 nsew ground input
rlabel locali s 298660 115855 298816 115889 6 VGND
port 614 nsew ground input
rlabel locali s 298660 115889 298799 116039 6 VGND
port 614 nsew ground input
rlabel locali s 1121 115705 1340 115855 6 VGND
port 614 nsew ground input
rlabel locali s 1104 115855 1340 115889 6 VGND
port 614 nsew ground input
rlabel locali s 1121 115889 1340 116039 6 VGND
port 614 nsew ground input
rlabel locali s 298695 116039 298799 116147 6 VGND
port 614 nsew ground input
rlabel locali s 1121 116039 1225 116147 6 VGND
port 614 nsew ground input
rlabel locali s 298695 116685 298799 116793 6 VGND
port 614 nsew ground input
rlabel locali s 1121 116685 1225 116793 6 VGND
port 614 nsew ground input
rlabel locali s 298660 116793 298799 116943 6 VGND
port 614 nsew ground input
rlabel locali s 298660 116943 298816 116977 6 VGND
port 614 nsew ground input
rlabel locali s 298660 116977 298799 117127 6 VGND
port 614 nsew ground input
rlabel locali s 1121 116793 1340 116943 6 VGND
port 614 nsew ground input
rlabel locali s 1104 116943 1340 116977 6 VGND
port 614 nsew ground input
rlabel locali s 1121 116977 1340 117127 6 VGND
port 614 nsew ground input
rlabel locali s 298695 117127 298799 117235 6 VGND
port 614 nsew ground input
rlabel locali s 1121 117127 1225 117235 6 VGND
port 614 nsew ground input
rlabel locali s 298695 117773 298799 117881 6 VGND
port 614 nsew ground input
rlabel locali s 1121 117773 1225 117881 6 VGND
port 614 nsew ground input
rlabel locali s 298660 117881 298799 118031 6 VGND
port 614 nsew ground input
rlabel locali s 298660 118031 298816 118065 6 VGND
port 614 nsew ground input
rlabel locali s 298660 118065 298799 118215 6 VGND
port 614 nsew ground input
rlabel locali s 1121 117881 1340 118031 6 VGND
port 614 nsew ground input
rlabel locali s 1104 118031 1340 118065 6 VGND
port 614 nsew ground input
rlabel locali s 1121 118065 1340 118215 6 VGND
port 614 nsew ground input
rlabel locali s 298695 118215 298799 118323 6 VGND
port 614 nsew ground input
rlabel locali s 1121 118215 1225 118323 6 VGND
port 614 nsew ground input
rlabel locali s 298695 118861 298799 118969 6 VGND
port 614 nsew ground input
rlabel locali s 1121 118861 1225 118969 6 VGND
port 614 nsew ground input
rlabel locali s 298660 118969 298799 119119 6 VGND
port 614 nsew ground input
rlabel locali s 298660 119119 298816 119153 6 VGND
port 614 nsew ground input
rlabel locali s 298660 119153 298799 119303 6 VGND
port 614 nsew ground input
rlabel locali s 1121 118969 1340 119119 6 VGND
port 614 nsew ground input
rlabel locali s 1104 119119 1340 119153 6 VGND
port 614 nsew ground input
rlabel locali s 1121 119153 1340 119303 6 VGND
port 614 nsew ground input
rlabel locali s 298695 119303 298799 119411 6 VGND
port 614 nsew ground input
rlabel locali s 1121 119303 1225 119411 6 VGND
port 614 nsew ground input
rlabel locali s 298695 119949 298799 120057 6 VGND
port 614 nsew ground input
rlabel locali s 1121 119949 1225 120057 6 VGND
port 614 nsew ground input
rlabel locali s 298660 120057 298799 120207 6 VGND
port 614 nsew ground input
rlabel locali s 298660 120207 298816 120241 6 VGND
port 614 nsew ground input
rlabel locali s 298660 120241 298799 120391 6 VGND
port 614 nsew ground input
rlabel locali s 1121 120057 1340 120207 6 VGND
port 614 nsew ground input
rlabel locali s 1104 120207 1340 120241 6 VGND
port 614 nsew ground input
rlabel locali s 1121 120241 1340 120391 6 VGND
port 614 nsew ground input
rlabel locali s 298695 120391 298799 120499 6 VGND
port 614 nsew ground input
rlabel locali s 1121 120391 1225 120499 6 VGND
port 614 nsew ground input
rlabel locali s 298695 121037 298799 121145 6 VGND
port 614 nsew ground input
rlabel locali s 1121 121037 1225 121145 6 VGND
port 614 nsew ground input
rlabel locali s 298660 121145 298799 121295 6 VGND
port 614 nsew ground input
rlabel locali s 298660 121295 298816 121329 6 VGND
port 614 nsew ground input
rlabel locali s 298660 121329 298799 121479 6 VGND
port 614 nsew ground input
rlabel locali s 1121 121145 1340 121295 6 VGND
port 614 nsew ground input
rlabel locali s 1104 121295 1340 121329 6 VGND
port 614 nsew ground input
rlabel locali s 1121 121329 1340 121479 6 VGND
port 614 nsew ground input
rlabel locali s 298695 121479 298799 121587 6 VGND
port 614 nsew ground input
rlabel locali s 1121 121479 1225 121587 6 VGND
port 614 nsew ground input
rlabel locali s 298695 122125 298799 122233 6 VGND
port 614 nsew ground input
rlabel locali s 1121 122125 1225 122233 6 VGND
port 614 nsew ground input
rlabel locali s 298660 122233 298799 122383 6 VGND
port 614 nsew ground input
rlabel locali s 298660 122383 298816 122417 6 VGND
port 614 nsew ground input
rlabel locali s 298660 122417 298799 122567 6 VGND
port 614 nsew ground input
rlabel locali s 1121 122233 1340 122383 6 VGND
port 614 nsew ground input
rlabel locali s 1104 122383 1340 122417 6 VGND
port 614 nsew ground input
rlabel locali s 1121 122417 1340 122567 6 VGND
port 614 nsew ground input
rlabel locali s 298695 122567 298799 122675 6 VGND
port 614 nsew ground input
rlabel locali s 1121 122567 1225 122675 6 VGND
port 614 nsew ground input
rlabel locali s 298695 123213 298799 123321 6 VGND
port 614 nsew ground input
rlabel locali s 1121 123213 1225 123321 6 VGND
port 614 nsew ground input
rlabel locali s 298660 123321 298799 123471 6 VGND
port 614 nsew ground input
rlabel locali s 298660 123471 298816 123505 6 VGND
port 614 nsew ground input
rlabel locali s 298660 123505 298799 123655 6 VGND
port 614 nsew ground input
rlabel locali s 1121 123321 1340 123471 6 VGND
port 614 nsew ground input
rlabel locali s 1104 123471 1340 123505 6 VGND
port 614 nsew ground input
rlabel locali s 1121 123505 1340 123655 6 VGND
port 614 nsew ground input
rlabel locali s 298695 123655 298799 123763 6 VGND
port 614 nsew ground input
rlabel locali s 1121 123655 1225 123763 6 VGND
port 614 nsew ground input
rlabel locali s 298695 124301 298799 124409 6 VGND
port 614 nsew ground input
rlabel locali s 1121 124301 1225 124409 6 VGND
port 614 nsew ground input
rlabel locali s 298660 124409 298799 124559 6 VGND
port 614 nsew ground input
rlabel locali s 298660 124559 298816 124593 6 VGND
port 614 nsew ground input
rlabel locali s 298660 124593 298799 124743 6 VGND
port 614 nsew ground input
rlabel locali s 1121 124409 1340 124559 6 VGND
port 614 nsew ground input
rlabel locali s 1104 124559 1340 124593 6 VGND
port 614 nsew ground input
rlabel locali s 1121 124593 1340 124743 6 VGND
port 614 nsew ground input
rlabel locali s 298695 124743 298799 124851 6 VGND
port 614 nsew ground input
rlabel locali s 1121 124743 1225 124851 6 VGND
port 614 nsew ground input
rlabel locali s 298695 125389 298799 125497 6 VGND
port 614 nsew ground input
rlabel locali s 1121 125389 1225 125497 6 VGND
port 614 nsew ground input
rlabel locali s 298660 125497 298799 125647 6 VGND
port 614 nsew ground input
rlabel locali s 298660 125647 298816 125681 6 VGND
port 614 nsew ground input
rlabel locali s 298660 125681 298799 125831 6 VGND
port 614 nsew ground input
rlabel locali s 1121 125497 1340 125647 6 VGND
port 614 nsew ground input
rlabel locali s 1104 125647 1340 125681 6 VGND
port 614 nsew ground input
rlabel locali s 1121 125681 1340 125831 6 VGND
port 614 nsew ground input
rlabel locali s 298695 125831 298799 125939 6 VGND
port 614 nsew ground input
rlabel locali s 1121 125831 1225 125939 6 VGND
port 614 nsew ground input
rlabel locali s 298695 126477 298799 126585 6 VGND
port 614 nsew ground input
rlabel locali s 1121 126477 1225 126585 6 VGND
port 614 nsew ground input
rlabel locali s 298660 126585 298799 126735 6 VGND
port 614 nsew ground input
rlabel locali s 298660 126735 298816 126769 6 VGND
port 614 nsew ground input
rlabel locali s 298660 126769 298799 126919 6 VGND
port 614 nsew ground input
rlabel locali s 1121 126585 1340 126735 6 VGND
port 614 nsew ground input
rlabel locali s 1104 126735 1340 126769 6 VGND
port 614 nsew ground input
rlabel locali s 1121 126769 1340 126919 6 VGND
port 614 nsew ground input
rlabel locali s 298695 126919 298799 127027 6 VGND
port 614 nsew ground input
rlabel locali s 1121 126919 1225 127027 6 VGND
port 614 nsew ground input
rlabel locali s 298695 127565 298799 127673 6 VGND
port 614 nsew ground input
rlabel locali s 1121 127565 1225 127673 6 VGND
port 614 nsew ground input
rlabel locali s 298660 127673 298799 127823 6 VGND
port 614 nsew ground input
rlabel locali s 298660 127823 298816 127857 6 VGND
port 614 nsew ground input
rlabel locali s 298660 127857 298799 128007 6 VGND
port 614 nsew ground input
rlabel locali s 1121 127673 1340 127823 6 VGND
port 614 nsew ground input
rlabel locali s 1104 127823 1340 127857 6 VGND
port 614 nsew ground input
rlabel locali s 1121 127857 1340 128007 6 VGND
port 614 nsew ground input
rlabel locali s 298695 128007 298799 128115 6 VGND
port 614 nsew ground input
rlabel locali s 1121 128007 1225 128115 6 VGND
port 614 nsew ground input
rlabel locali s 298695 128653 298799 128761 6 VGND
port 614 nsew ground input
rlabel locali s 1121 128653 1225 128761 6 VGND
port 614 nsew ground input
rlabel locali s 298660 128761 298799 128911 6 VGND
port 614 nsew ground input
rlabel locali s 298660 128911 298816 128945 6 VGND
port 614 nsew ground input
rlabel locali s 298660 128945 298799 129095 6 VGND
port 614 nsew ground input
rlabel locali s 1121 128761 1340 128911 6 VGND
port 614 nsew ground input
rlabel locali s 1104 128911 1340 128945 6 VGND
port 614 nsew ground input
rlabel locali s 1121 128945 1340 129095 6 VGND
port 614 nsew ground input
rlabel locali s 298695 129095 298799 129203 6 VGND
port 614 nsew ground input
rlabel locali s 1121 129095 1225 129203 6 VGND
port 614 nsew ground input
rlabel locali s 298695 129741 298799 129849 6 VGND
port 614 nsew ground input
rlabel locali s 1121 129741 1225 129849 6 VGND
port 614 nsew ground input
rlabel locali s 298660 129849 298799 129999 6 VGND
port 614 nsew ground input
rlabel locali s 298660 129999 298816 130033 6 VGND
port 614 nsew ground input
rlabel locali s 298660 130033 298799 130183 6 VGND
port 614 nsew ground input
rlabel locali s 1121 129849 1340 129999 6 VGND
port 614 nsew ground input
rlabel locali s 1104 129999 1340 130033 6 VGND
port 614 nsew ground input
rlabel locali s 1121 130033 1340 130183 6 VGND
port 614 nsew ground input
rlabel locali s 298695 130183 298799 130291 6 VGND
port 614 nsew ground input
rlabel locali s 1121 130183 1225 130291 6 VGND
port 614 nsew ground input
rlabel locali s 298695 130829 298799 130937 6 VGND
port 614 nsew ground input
rlabel locali s 1121 130829 1225 130937 6 VGND
port 614 nsew ground input
rlabel locali s 298660 130937 298799 131087 6 VGND
port 614 nsew ground input
rlabel locali s 298660 131087 298816 131121 6 VGND
port 614 nsew ground input
rlabel locali s 298660 131121 298799 131271 6 VGND
port 614 nsew ground input
rlabel locali s 1121 130937 1340 131087 6 VGND
port 614 nsew ground input
rlabel locali s 1104 131087 1340 131121 6 VGND
port 614 nsew ground input
rlabel locali s 1121 131121 1340 131271 6 VGND
port 614 nsew ground input
rlabel locali s 298695 131271 298799 131379 6 VGND
port 614 nsew ground input
rlabel locali s 1121 131271 1225 131379 6 VGND
port 614 nsew ground input
rlabel locali s 298695 131917 298799 132025 6 VGND
port 614 nsew ground input
rlabel locali s 1121 131917 1225 132025 6 VGND
port 614 nsew ground input
rlabel locali s 298660 132025 298799 132175 6 VGND
port 614 nsew ground input
rlabel locali s 298660 132175 298816 132209 6 VGND
port 614 nsew ground input
rlabel locali s 298660 132209 298799 132359 6 VGND
port 614 nsew ground input
rlabel locali s 1121 132025 1340 132175 6 VGND
port 614 nsew ground input
rlabel locali s 1104 132175 1340 132209 6 VGND
port 614 nsew ground input
rlabel locali s 1121 132209 1340 132359 6 VGND
port 614 nsew ground input
rlabel locali s 298695 132359 298799 132467 6 VGND
port 614 nsew ground input
rlabel locali s 1121 132359 1225 132467 6 VGND
port 614 nsew ground input
rlabel locali s 298695 133005 298799 133113 6 VGND
port 614 nsew ground input
rlabel locali s 1121 133005 1225 133113 6 VGND
port 614 nsew ground input
rlabel locali s 298660 133113 298799 133263 6 VGND
port 614 nsew ground input
rlabel locali s 298660 133263 298816 133297 6 VGND
port 614 nsew ground input
rlabel locali s 298660 133297 298799 133447 6 VGND
port 614 nsew ground input
rlabel locali s 1121 133113 1340 133263 6 VGND
port 614 nsew ground input
rlabel locali s 1104 133263 1340 133297 6 VGND
port 614 nsew ground input
rlabel locali s 1121 133297 1340 133447 6 VGND
port 614 nsew ground input
rlabel locali s 298695 133447 298799 133555 6 VGND
port 614 nsew ground input
rlabel locali s 1121 133447 1225 133555 6 VGND
port 614 nsew ground input
rlabel locali s 298695 134093 298799 134201 6 VGND
port 614 nsew ground input
rlabel locali s 1121 134093 1225 134201 6 VGND
port 614 nsew ground input
rlabel locali s 298660 134201 298799 134351 6 VGND
port 614 nsew ground input
rlabel locali s 298660 134351 298816 134385 6 VGND
port 614 nsew ground input
rlabel locali s 298660 134385 298799 134535 6 VGND
port 614 nsew ground input
rlabel locali s 1121 134201 1340 134351 6 VGND
port 614 nsew ground input
rlabel locali s 1104 134351 1340 134385 6 VGND
port 614 nsew ground input
rlabel locali s 1121 134385 1340 134535 6 VGND
port 614 nsew ground input
rlabel locali s 298695 134535 298799 134643 6 VGND
port 614 nsew ground input
rlabel locali s 1121 134535 1225 134643 6 VGND
port 614 nsew ground input
rlabel locali s 298695 135181 298799 135289 6 VGND
port 614 nsew ground input
rlabel locali s 1121 135181 1225 135289 6 VGND
port 614 nsew ground input
rlabel locali s 298660 135289 298799 135439 6 VGND
port 614 nsew ground input
rlabel locali s 298660 135439 298816 135473 6 VGND
port 614 nsew ground input
rlabel locali s 298660 135473 298799 135623 6 VGND
port 614 nsew ground input
rlabel locali s 1121 135289 1340 135439 6 VGND
port 614 nsew ground input
rlabel locali s 1104 135439 1340 135473 6 VGND
port 614 nsew ground input
rlabel locali s 1121 135473 1340 135623 6 VGND
port 614 nsew ground input
rlabel locali s 298695 135623 298799 135731 6 VGND
port 614 nsew ground input
rlabel locali s 1121 135623 1225 135731 6 VGND
port 614 nsew ground input
rlabel locali s 298695 136269 298799 136377 6 VGND
port 614 nsew ground input
rlabel locali s 1121 136269 1225 136377 6 VGND
port 614 nsew ground input
rlabel locali s 298660 136377 298799 136527 6 VGND
port 614 nsew ground input
rlabel locali s 298660 136527 298816 136561 6 VGND
port 614 nsew ground input
rlabel locali s 298660 136561 298799 136711 6 VGND
port 614 nsew ground input
rlabel locali s 1121 136377 1340 136527 6 VGND
port 614 nsew ground input
rlabel locali s 1104 136527 1340 136561 6 VGND
port 614 nsew ground input
rlabel locali s 1121 136561 1340 136711 6 VGND
port 614 nsew ground input
rlabel locali s 298695 136711 298799 136819 6 VGND
port 614 nsew ground input
rlabel locali s 1121 136711 1225 136819 6 VGND
port 614 nsew ground input
rlabel locali s 298695 137357 298799 137465 6 VGND
port 614 nsew ground input
rlabel locali s 1121 137357 1225 137465 6 VGND
port 614 nsew ground input
rlabel locali s 298660 137465 298799 137615 6 VGND
port 614 nsew ground input
rlabel locali s 298660 137615 298816 137649 6 VGND
port 614 nsew ground input
rlabel locali s 298660 137649 298799 137799 6 VGND
port 614 nsew ground input
rlabel locali s 1121 137465 1340 137615 6 VGND
port 614 nsew ground input
rlabel locali s 1104 137615 1340 137649 6 VGND
port 614 nsew ground input
rlabel locali s 1121 137649 1340 137799 6 VGND
port 614 nsew ground input
rlabel locali s 298695 137799 298799 137907 6 VGND
port 614 nsew ground input
rlabel locali s 1121 137799 1225 137907 6 VGND
port 614 nsew ground input
rlabel locali s 298695 138445 298799 138553 6 VGND
port 614 nsew ground input
rlabel locali s 1121 138445 1225 138553 6 VGND
port 614 nsew ground input
rlabel locali s 298660 138553 298799 138703 6 VGND
port 614 nsew ground input
rlabel locali s 298660 138703 298816 138737 6 VGND
port 614 nsew ground input
rlabel locali s 298660 138737 298799 138887 6 VGND
port 614 nsew ground input
rlabel locali s 1121 138553 1340 138703 6 VGND
port 614 nsew ground input
rlabel locali s 1104 138703 1340 138737 6 VGND
port 614 nsew ground input
rlabel locali s 1121 138737 1340 138887 6 VGND
port 614 nsew ground input
rlabel locali s 298695 138887 298799 138995 6 VGND
port 614 nsew ground input
rlabel locali s 1121 138887 1225 138995 6 VGND
port 614 nsew ground input
rlabel locali s 298695 139533 298799 139641 6 VGND
port 614 nsew ground input
rlabel locali s 1121 139533 1225 139641 6 VGND
port 614 nsew ground input
rlabel locali s 298660 139641 298799 139791 6 VGND
port 614 nsew ground input
rlabel locali s 298660 139791 298816 139825 6 VGND
port 614 nsew ground input
rlabel locali s 298660 139825 298799 139975 6 VGND
port 614 nsew ground input
rlabel locali s 1121 139641 1340 139791 6 VGND
port 614 nsew ground input
rlabel locali s 1104 139791 1340 139825 6 VGND
port 614 nsew ground input
rlabel locali s 1121 139825 1340 139975 6 VGND
port 614 nsew ground input
rlabel locali s 298695 139975 298799 140083 6 VGND
port 614 nsew ground input
rlabel locali s 1121 139975 1225 140083 6 VGND
port 614 nsew ground input
rlabel locali s 298695 140621 298799 140729 6 VGND
port 614 nsew ground input
rlabel locali s 1121 140621 1225 140729 6 VGND
port 614 nsew ground input
rlabel locali s 298660 140729 298799 140879 6 VGND
port 614 nsew ground input
rlabel locali s 298660 140879 298816 140913 6 VGND
port 614 nsew ground input
rlabel locali s 298660 140913 298799 141063 6 VGND
port 614 nsew ground input
rlabel locali s 1121 140729 1340 140879 6 VGND
port 614 nsew ground input
rlabel locali s 1104 140879 1340 140913 6 VGND
port 614 nsew ground input
rlabel locali s 1121 140913 1340 141063 6 VGND
port 614 nsew ground input
rlabel locali s 298695 141063 298799 141171 6 VGND
port 614 nsew ground input
rlabel locali s 1121 141063 1225 141171 6 VGND
port 614 nsew ground input
rlabel locali s 298695 141709 298799 141817 6 VGND
port 614 nsew ground input
rlabel locali s 1121 141709 1225 141817 6 VGND
port 614 nsew ground input
rlabel locali s 298660 141817 298799 141967 6 VGND
port 614 nsew ground input
rlabel locali s 298660 141967 298816 142001 6 VGND
port 614 nsew ground input
rlabel locali s 298660 142001 298799 142151 6 VGND
port 614 nsew ground input
rlabel locali s 1121 141817 1340 141967 6 VGND
port 614 nsew ground input
rlabel locali s 1104 141967 1340 142001 6 VGND
port 614 nsew ground input
rlabel locali s 1121 142001 1340 142151 6 VGND
port 614 nsew ground input
rlabel locali s 298695 142151 298799 142259 6 VGND
port 614 nsew ground input
rlabel locali s 1121 142151 1225 142259 6 VGND
port 614 nsew ground input
rlabel locali s 298695 142797 298799 142905 6 VGND
port 614 nsew ground input
rlabel locali s 1121 142797 1225 142905 6 VGND
port 614 nsew ground input
rlabel locali s 298660 142905 298799 143055 6 VGND
port 614 nsew ground input
rlabel locali s 298660 143055 298816 143089 6 VGND
port 614 nsew ground input
rlabel locali s 298660 143089 298799 143239 6 VGND
port 614 nsew ground input
rlabel locali s 1121 142905 1340 143055 6 VGND
port 614 nsew ground input
rlabel locali s 1104 143055 1340 143089 6 VGND
port 614 nsew ground input
rlabel locali s 1121 143089 1340 143239 6 VGND
port 614 nsew ground input
rlabel locali s 298695 143239 298799 143347 6 VGND
port 614 nsew ground input
rlabel locali s 1121 143239 1225 143347 6 VGND
port 614 nsew ground input
rlabel locali s 298695 143885 298799 143993 6 VGND
port 614 nsew ground input
rlabel locali s 1121 143885 1225 143993 6 VGND
port 614 nsew ground input
rlabel locali s 298660 143993 298799 144143 6 VGND
port 614 nsew ground input
rlabel locali s 298660 144143 298816 144177 6 VGND
port 614 nsew ground input
rlabel locali s 298660 144177 298799 144327 6 VGND
port 614 nsew ground input
rlabel locali s 1121 143993 1340 144143 6 VGND
port 614 nsew ground input
rlabel locali s 1104 144143 1340 144177 6 VGND
port 614 nsew ground input
rlabel locali s 1121 144177 1340 144327 6 VGND
port 614 nsew ground input
rlabel locali s 298695 144327 298799 144435 6 VGND
port 614 nsew ground input
rlabel locali s 1121 144327 1225 144435 6 VGND
port 614 nsew ground input
rlabel locali s 298695 144973 298799 145081 6 VGND
port 614 nsew ground input
rlabel locali s 1121 144973 1225 145081 6 VGND
port 614 nsew ground input
rlabel locali s 298660 145081 298799 145231 6 VGND
port 614 nsew ground input
rlabel locali s 298660 145231 298816 145265 6 VGND
port 614 nsew ground input
rlabel locali s 298660 145265 298799 145415 6 VGND
port 614 nsew ground input
rlabel locali s 1121 145081 1340 145231 6 VGND
port 614 nsew ground input
rlabel locali s 1104 145231 1340 145265 6 VGND
port 614 nsew ground input
rlabel locali s 1121 145265 1340 145415 6 VGND
port 614 nsew ground input
rlabel locali s 298695 145415 298799 145523 6 VGND
port 614 nsew ground input
rlabel locali s 1121 145415 1225 145523 6 VGND
port 614 nsew ground input
rlabel locali s 298695 146061 298799 146169 6 VGND
port 614 nsew ground input
rlabel locali s 1121 146061 1225 146169 6 VGND
port 614 nsew ground input
rlabel locali s 298660 146169 298799 146319 6 VGND
port 614 nsew ground input
rlabel locali s 298660 146319 298816 146353 6 VGND
port 614 nsew ground input
rlabel locali s 298660 146353 298799 146503 6 VGND
port 614 nsew ground input
rlabel locali s 1121 146169 1340 146319 6 VGND
port 614 nsew ground input
rlabel locali s 1104 146319 1340 146353 6 VGND
port 614 nsew ground input
rlabel locali s 1121 146353 1340 146503 6 VGND
port 614 nsew ground input
rlabel locali s 298695 146503 298799 146611 6 VGND
port 614 nsew ground input
rlabel locali s 1121 146503 1225 146611 6 VGND
port 614 nsew ground input
rlabel locali s 298695 147149 298799 147257 6 VGND
port 614 nsew ground input
rlabel locali s 1121 147149 1225 147257 6 VGND
port 614 nsew ground input
rlabel locali s 298660 147257 298799 147407 6 VGND
port 614 nsew ground input
rlabel locali s 298660 147407 298816 147441 6 VGND
port 614 nsew ground input
rlabel locali s 298660 147441 298799 147591 6 VGND
port 614 nsew ground input
rlabel locali s 1121 147257 1340 147407 6 VGND
port 614 nsew ground input
rlabel locali s 1104 147407 1340 147441 6 VGND
port 614 nsew ground input
rlabel locali s 1121 147441 1340 147591 6 VGND
port 614 nsew ground input
rlabel locali s 298695 147591 298799 147699 6 VGND
port 614 nsew ground input
rlabel locali s 1121 147591 1225 147699 6 VGND
port 614 nsew ground input
rlabel locali s 298695 148237 298799 148345 6 VGND
port 614 nsew ground input
rlabel locali s 1121 148237 1225 148345 6 VGND
port 614 nsew ground input
rlabel locali s 298660 148345 298799 148495 6 VGND
port 614 nsew ground input
rlabel locali s 298660 148495 298816 148529 6 VGND
port 614 nsew ground input
rlabel locali s 298660 148529 298799 148679 6 VGND
port 614 nsew ground input
rlabel locali s 1121 148345 1340 148495 6 VGND
port 614 nsew ground input
rlabel locali s 1104 148495 1340 148529 6 VGND
port 614 nsew ground input
rlabel locali s 1121 148529 1340 148679 6 VGND
port 614 nsew ground input
rlabel locali s 298695 148679 298799 148787 6 VGND
port 614 nsew ground input
rlabel locali s 1121 148679 1225 148787 6 VGND
port 614 nsew ground input
rlabel locali s 298695 149325 298799 149433 6 VGND
port 614 nsew ground input
rlabel locali s 1121 149325 1225 149433 6 VGND
port 614 nsew ground input
rlabel locali s 298660 149433 298799 149583 6 VGND
port 614 nsew ground input
rlabel locali s 298660 149583 298816 149617 6 VGND
port 614 nsew ground input
rlabel locali s 298660 149617 298799 149767 6 VGND
port 614 nsew ground input
rlabel locali s 1121 149433 1340 149583 6 VGND
port 614 nsew ground input
rlabel locali s 1104 149583 1340 149617 6 VGND
port 614 nsew ground input
rlabel locali s 1121 149617 1340 149767 6 VGND
port 614 nsew ground input
rlabel locali s 298695 149767 298799 149875 6 VGND
port 614 nsew ground input
rlabel locali s 1121 149767 1225 149875 6 VGND
port 614 nsew ground input
rlabel locali s 298695 150413 298799 150521 6 VGND
port 614 nsew ground input
rlabel locali s 1121 150413 1225 150521 6 VGND
port 614 nsew ground input
rlabel locali s 298660 150521 298799 150671 6 VGND
port 614 nsew ground input
rlabel locali s 298660 150671 298816 150705 6 VGND
port 614 nsew ground input
rlabel locali s 298660 150705 298799 150855 6 VGND
port 614 nsew ground input
rlabel locali s 1121 150521 1340 150671 6 VGND
port 614 nsew ground input
rlabel locali s 1104 150671 1340 150705 6 VGND
port 614 nsew ground input
rlabel locali s 1121 150705 1340 150855 6 VGND
port 614 nsew ground input
rlabel locali s 298695 150855 298799 150963 6 VGND
port 614 nsew ground input
rlabel locali s 1121 150855 1225 150963 6 VGND
port 614 nsew ground input
rlabel locali s 298695 151501 298799 151609 6 VGND
port 614 nsew ground input
rlabel locali s 1121 151501 1225 151609 6 VGND
port 614 nsew ground input
rlabel locali s 298660 151609 298799 151759 6 VGND
port 614 nsew ground input
rlabel locali s 298660 151759 298816 151793 6 VGND
port 614 nsew ground input
rlabel locali s 298660 151793 298799 151943 6 VGND
port 614 nsew ground input
rlabel locali s 1121 151609 1340 151759 6 VGND
port 614 nsew ground input
rlabel locali s 1104 151759 1340 151793 6 VGND
port 614 nsew ground input
rlabel locali s 1121 151793 1340 151943 6 VGND
port 614 nsew ground input
rlabel locali s 298695 151943 298799 152051 6 VGND
port 614 nsew ground input
rlabel locali s 1121 151943 1225 152051 6 VGND
port 614 nsew ground input
rlabel locali s 298695 152589 298799 152697 6 VGND
port 614 nsew ground input
rlabel locali s 1121 152589 1225 152697 6 VGND
port 614 nsew ground input
rlabel locali s 298660 152697 298799 152847 6 VGND
port 614 nsew ground input
rlabel locali s 298660 152847 298816 152881 6 VGND
port 614 nsew ground input
rlabel locali s 298660 152881 298799 153031 6 VGND
port 614 nsew ground input
rlabel locali s 1121 152697 1340 152847 6 VGND
port 614 nsew ground input
rlabel locali s 1104 152847 1340 152881 6 VGND
port 614 nsew ground input
rlabel locali s 1121 152881 1340 153031 6 VGND
port 614 nsew ground input
rlabel locali s 298695 153031 298799 153139 6 VGND
port 614 nsew ground input
rlabel locali s 1121 153031 1225 153139 6 VGND
port 614 nsew ground input
rlabel locali s 298695 153677 298799 153785 6 VGND
port 614 nsew ground input
rlabel locali s 1121 153677 1225 153785 6 VGND
port 614 nsew ground input
rlabel locali s 298660 153785 298799 153935 6 VGND
port 614 nsew ground input
rlabel locali s 298660 153935 298816 153969 6 VGND
port 614 nsew ground input
rlabel locali s 298660 153969 298799 154119 6 VGND
port 614 nsew ground input
rlabel locali s 1121 153785 1340 153935 6 VGND
port 614 nsew ground input
rlabel locali s 1104 153935 1340 153969 6 VGND
port 614 nsew ground input
rlabel locali s 1121 153969 1340 154119 6 VGND
port 614 nsew ground input
rlabel locali s 298695 154119 298799 154227 6 VGND
port 614 nsew ground input
rlabel locali s 1121 154119 1225 154227 6 VGND
port 614 nsew ground input
rlabel locali s 298695 154765 298799 154873 6 VGND
port 614 nsew ground input
rlabel locali s 1121 154765 1225 154873 6 VGND
port 614 nsew ground input
rlabel locali s 298660 154873 298799 155023 6 VGND
port 614 nsew ground input
rlabel locali s 298660 155023 298816 155057 6 VGND
port 614 nsew ground input
rlabel locali s 298660 155057 298799 155207 6 VGND
port 614 nsew ground input
rlabel locali s 1121 154873 1340 155023 6 VGND
port 614 nsew ground input
rlabel locali s 1104 155023 1340 155057 6 VGND
port 614 nsew ground input
rlabel locali s 1121 155057 1340 155207 6 VGND
port 614 nsew ground input
rlabel locali s 298695 155207 298799 155315 6 VGND
port 614 nsew ground input
rlabel locali s 1121 155207 1225 155315 6 VGND
port 614 nsew ground input
rlabel locali s 298695 155853 298799 155961 6 VGND
port 614 nsew ground input
rlabel locali s 1121 155853 1225 155961 6 VGND
port 614 nsew ground input
rlabel locali s 298660 155961 298799 156111 6 VGND
port 614 nsew ground input
rlabel locali s 298660 156111 298816 156145 6 VGND
port 614 nsew ground input
rlabel locali s 298660 156145 298799 156295 6 VGND
port 614 nsew ground input
rlabel locali s 1121 155961 1340 156111 6 VGND
port 614 nsew ground input
rlabel locali s 1104 156111 1340 156145 6 VGND
port 614 nsew ground input
rlabel locali s 1121 156145 1340 156295 6 VGND
port 614 nsew ground input
rlabel locali s 298695 156295 298799 156403 6 VGND
port 614 nsew ground input
rlabel locali s 1121 156295 1225 156403 6 VGND
port 614 nsew ground input
rlabel locali s 298695 156941 298799 157049 6 VGND
port 614 nsew ground input
rlabel locali s 1121 156941 1225 157049 6 VGND
port 614 nsew ground input
rlabel locali s 298660 157049 298799 157199 6 VGND
port 614 nsew ground input
rlabel locali s 298660 157199 298816 157233 6 VGND
port 614 nsew ground input
rlabel locali s 298660 157233 298799 157383 6 VGND
port 614 nsew ground input
rlabel locali s 1121 157049 1340 157199 6 VGND
port 614 nsew ground input
rlabel locali s 1104 157199 1340 157233 6 VGND
port 614 nsew ground input
rlabel locali s 1121 157233 1340 157383 6 VGND
port 614 nsew ground input
rlabel locali s 298695 157383 298799 157491 6 VGND
port 614 nsew ground input
rlabel locali s 1121 157383 1225 157491 6 VGND
port 614 nsew ground input
rlabel locali s 298695 158029 298799 158137 6 VGND
port 614 nsew ground input
rlabel locali s 1121 158029 1225 158137 6 VGND
port 614 nsew ground input
rlabel locali s 298660 158137 298799 158287 6 VGND
port 614 nsew ground input
rlabel locali s 298660 158287 298816 158321 6 VGND
port 614 nsew ground input
rlabel locali s 298660 158321 298799 158471 6 VGND
port 614 nsew ground input
rlabel locali s 1121 158137 1340 158287 6 VGND
port 614 nsew ground input
rlabel locali s 1104 158287 1340 158321 6 VGND
port 614 nsew ground input
rlabel locali s 1121 158321 1340 158471 6 VGND
port 614 nsew ground input
rlabel locali s 298695 158471 298799 158579 6 VGND
port 614 nsew ground input
rlabel locali s 1121 158471 1225 158579 6 VGND
port 614 nsew ground input
rlabel locali s 298695 159117 298799 159225 6 VGND
port 614 nsew ground input
rlabel locali s 1121 159117 1225 159225 6 VGND
port 614 nsew ground input
rlabel locali s 298660 159225 298799 159375 6 VGND
port 614 nsew ground input
rlabel locali s 298660 159375 298816 159409 6 VGND
port 614 nsew ground input
rlabel locali s 298660 159409 298799 159559 6 VGND
port 614 nsew ground input
rlabel locali s 1121 159225 1340 159375 6 VGND
port 614 nsew ground input
rlabel locali s 1104 159375 1340 159409 6 VGND
port 614 nsew ground input
rlabel locali s 1121 159409 1340 159559 6 VGND
port 614 nsew ground input
rlabel locali s 298695 159559 298799 159667 6 VGND
port 614 nsew ground input
rlabel locali s 1121 159559 1225 159667 6 VGND
port 614 nsew ground input
rlabel locali s 298695 160205 298799 160313 6 VGND
port 614 nsew ground input
rlabel locali s 1121 160205 1225 160313 6 VGND
port 614 nsew ground input
rlabel locali s 298660 160313 298799 160463 6 VGND
port 614 nsew ground input
rlabel locali s 298660 160463 298816 160497 6 VGND
port 614 nsew ground input
rlabel locali s 298660 160497 298799 160647 6 VGND
port 614 nsew ground input
rlabel locali s 1121 160313 1340 160463 6 VGND
port 614 nsew ground input
rlabel locali s 1104 160463 1340 160497 6 VGND
port 614 nsew ground input
rlabel locali s 1121 160497 1340 160647 6 VGND
port 614 nsew ground input
rlabel locali s 298695 160647 298799 160755 6 VGND
port 614 nsew ground input
rlabel locali s 1121 160647 1225 160755 6 VGND
port 614 nsew ground input
rlabel locali s 298695 161293 298799 161401 6 VGND
port 614 nsew ground input
rlabel locali s 1121 161293 1225 161401 6 VGND
port 614 nsew ground input
rlabel locali s 298660 161401 298799 161551 6 VGND
port 614 nsew ground input
rlabel locali s 298660 161551 298816 161585 6 VGND
port 614 nsew ground input
rlabel locali s 298660 161585 298799 161735 6 VGND
port 614 nsew ground input
rlabel locali s 1121 161401 1340 161551 6 VGND
port 614 nsew ground input
rlabel locali s 1104 161551 1340 161585 6 VGND
port 614 nsew ground input
rlabel locali s 1121 161585 1340 161735 6 VGND
port 614 nsew ground input
rlabel locali s 298695 161735 298799 161843 6 VGND
port 614 nsew ground input
rlabel locali s 1121 161735 1225 161843 6 VGND
port 614 nsew ground input
rlabel locali s 298695 162381 298799 162489 6 VGND
port 614 nsew ground input
rlabel locali s 1121 162381 1225 162489 6 VGND
port 614 nsew ground input
rlabel locali s 298660 162489 298799 162639 6 VGND
port 614 nsew ground input
rlabel locali s 298660 162639 298816 162673 6 VGND
port 614 nsew ground input
rlabel locali s 298660 162673 298799 162823 6 VGND
port 614 nsew ground input
rlabel locali s 1121 162489 1340 162639 6 VGND
port 614 nsew ground input
rlabel locali s 1104 162639 1340 162673 6 VGND
port 614 nsew ground input
rlabel locali s 1121 162673 1340 162823 6 VGND
port 614 nsew ground input
rlabel locali s 298695 162823 298799 162931 6 VGND
port 614 nsew ground input
rlabel locali s 1121 162823 1225 162931 6 VGND
port 614 nsew ground input
rlabel locali s 298695 163469 298799 163577 6 VGND
port 614 nsew ground input
rlabel locali s 1121 163469 1225 163577 6 VGND
port 614 nsew ground input
rlabel locali s 298660 163577 298799 163727 6 VGND
port 614 nsew ground input
rlabel locali s 298660 163727 298816 163761 6 VGND
port 614 nsew ground input
rlabel locali s 298660 163761 298799 163911 6 VGND
port 614 nsew ground input
rlabel locali s 1121 163577 1340 163727 6 VGND
port 614 nsew ground input
rlabel locali s 1104 163727 1340 163761 6 VGND
port 614 nsew ground input
rlabel locali s 1121 163761 1340 163911 6 VGND
port 614 nsew ground input
rlabel locali s 298695 163911 298799 164019 6 VGND
port 614 nsew ground input
rlabel locali s 1121 163911 1225 164019 6 VGND
port 614 nsew ground input
rlabel locali s 298695 164557 298799 164665 6 VGND
port 614 nsew ground input
rlabel locali s 1121 164557 1225 164665 6 VGND
port 614 nsew ground input
rlabel locali s 298660 164665 298799 164815 6 VGND
port 614 nsew ground input
rlabel locali s 298660 164815 298816 164849 6 VGND
port 614 nsew ground input
rlabel locali s 298660 164849 298799 164999 6 VGND
port 614 nsew ground input
rlabel locali s 1121 164665 1340 164815 6 VGND
port 614 nsew ground input
rlabel locali s 1104 164815 1340 164849 6 VGND
port 614 nsew ground input
rlabel locali s 1121 164849 1340 164999 6 VGND
port 614 nsew ground input
rlabel locali s 298695 164999 298799 165107 6 VGND
port 614 nsew ground input
rlabel locali s 1121 164999 1225 165107 6 VGND
port 614 nsew ground input
rlabel locali s 298695 165645 298799 165753 6 VGND
port 614 nsew ground input
rlabel locali s 1121 165645 1225 165753 6 VGND
port 614 nsew ground input
rlabel locali s 298660 165753 298799 165903 6 VGND
port 614 nsew ground input
rlabel locali s 298660 165903 298816 165937 6 VGND
port 614 nsew ground input
rlabel locali s 298660 165937 298799 166087 6 VGND
port 614 nsew ground input
rlabel locali s 1121 165753 1340 165903 6 VGND
port 614 nsew ground input
rlabel locali s 1104 165903 1340 165937 6 VGND
port 614 nsew ground input
rlabel locali s 1121 165937 1340 166087 6 VGND
port 614 nsew ground input
rlabel locali s 298695 166087 298799 166195 6 VGND
port 614 nsew ground input
rlabel locali s 1121 166087 1225 166195 6 VGND
port 614 nsew ground input
rlabel locali s 298695 166733 298799 166841 6 VGND
port 614 nsew ground input
rlabel locali s 1121 166733 1225 166841 6 VGND
port 614 nsew ground input
rlabel locali s 298660 166841 298799 166991 6 VGND
port 614 nsew ground input
rlabel locali s 298660 166991 298816 167025 6 VGND
port 614 nsew ground input
rlabel locali s 298660 167025 298799 167175 6 VGND
port 614 nsew ground input
rlabel locali s 1121 166841 1340 166991 6 VGND
port 614 nsew ground input
rlabel locali s 1104 166991 1340 167025 6 VGND
port 614 nsew ground input
rlabel locali s 1121 167025 1340 167175 6 VGND
port 614 nsew ground input
rlabel locali s 298695 167175 298799 167283 6 VGND
port 614 nsew ground input
rlabel locali s 1121 167175 1225 167283 6 VGND
port 614 nsew ground input
rlabel locali s 298695 167821 298799 167929 6 VGND
port 614 nsew ground input
rlabel locali s 1121 167821 1225 167929 6 VGND
port 614 nsew ground input
rlabel locali s 298660 167929 298799 168079 6 VGND
port 614 nsew ground input
rlabel locali s 298660 168079 298816 168113 6 VGND
port 614 nsew ground input
rlabel locali s 298660 168113 298799 168263 6 VGND
port 614 nsew ground input
rlabel locali s 1121 167929 1340 168079 6 VGND
port 614 nsew ground input
rlabel locali s 1104 168079 1340 168113 6 VGND
port 614 nsew ground input
rlabel locali s 1121 168113 1340 168263 6 VGND
port 614 nsew ground input
rlabel locali s 298695 168263 298799 168371 6 VGND
port 614 nsew ground input
rlabel locali s 1121 168263 1225 168371 6 VGND
port 614 nsew ground input
rlabel locali s 298695 168909 298799 169017 6 VGND
port 614 nsew ground input
rlabel locali s 1121 168909 1225 169017 6 VGND
port 614 nsew ground input
rlabel locali s 298660 169017 298799 169167 6 VGND
port 614 nsew ground input
rlabel locali s 298660 169167 298816 169201 6 VGND
port 614 nsew ground input
rlabel locali s 298660 169201 298799 169351 6 VGND
port 614 nsew ground input
rlabel locali s 1121 169017 1340 169167 6 VGND
port 614 nsew ground input
rlabel locali s 1104 169167 1340 169201 6 VGND
port 614 nsew ground input
rlabel locali s 1121 169201 1340 169351 6 VGND
port 614 nsew ground input
rlabel locali s 298695 169351 298799 169459 6 VGND
port 614 nsew ground input
rlabel locali s 1121 169351 1225 169459 6 VGND
port 614 nsew ground input
rlabel locali s 298695 169997 298799 170105 6 VGND
port 614 nsew ground input
rlabel locali s 1121 169997 1225 170105 6 VGND
port 614 nsew ground input
rlabel locali s 298660 170105 298799 170255 6 VGND
port 614 nsew ground input
rlabel locali s 298660 170255 298816 170289 6 VGND
port 614 nsew ground input
rlabel locali s 298660 170289 298799 170439 6 VGND
port 614 nsew ground input
rlabel locali s 1121 170105 1340 170255 6 VGND
port 614 nsew ground input
rlabel locali s 1104 170255 1340 170289 6 VGND
port 614 nsew ground input
rlabel locali s 1121 170289 1340 170439 6 VGND
port 614 nsew ground input
rlabel locali s 298695 170439 298799 170547 6 VGND
port 614 nsew ground input
rlabel locali s 1121 170439 1225 170547 6 VGND
port 614 nsew ground input
rlabel locali s 298695 171085 298799 171193 6 VGND
port 614 nsew ground input
rlabel locali s 1121 171085 1225 171193 6 VGND
port 614 nsew ground input
rlabel locali s 298660 171193 298799 171343 6 VGND
port 614 nsew ground input
rlabel locali s 298660 171343 298816 171377 6 VGND
port 614 nsew ground input
rlabel locali s 298660 171377 298799 171527 6 VGND
port 614 nsew ground input
rlabel locali s 1121 171193 1340 171343 6 VGND
port 614 nsew ground input
rlabel locali s 1104 171343 1340 171377 6 VGND
port 614 nsew ground input
rlabel locali s 1121 171377 1340 171527 6 VGND
port 614 nsew ground input
rlabel locali s 298695 171527 298799 171635 6 VGND
port 614 nsew ground input
rlabel locali s 1121 171527 1225 171635 6 VGND
port 614 nsew ground input
rlabel locali s 298695 172173 298799 172281 6 VGND
port 614 nsew ground input
rlabel locali s 1121 172173 1225 172281 6 VGND
port 614 nsew ground input
rlabel locali s 298660 172281 298799 172431 6 VGND
port 614 nsew ground input
rlabel locali s 298660 172431 298816 172465 6 VGND
port 614 nsew ground input
rlabel locali s 298660 172465 298799 172615 6 VGND
port 614 nsew ground input
rlabel locali s 1121 172281 1340 172431 6 VGND
port 614 nsew ground input
rlabel locali s 1104 172431 1340 172465 6 VGND
port 614 nsew ground input
rlabel locali s 1121 172465 1340 172615 6 VGND
port 614 nsew ground input
rlabel locali s 298695 172615 298799 172723 6 VGND
port 614 nsew ground input
rlabel locali s 1121 172615 1225 172723 6 VGND
port 614 nsew ground input
rlabel locali s 298695 173261 298799 173369 6 VGND
port 614 nsew ground input
rlabel locali s 1121 173261 1225 173369 6 VGND
port 614 nsew ground input
rlabel locali s 298660 173369 298799 173519 6 VGND
port 614 nsew ground input
rlabel locali s 298660 173519 298816 173553 6 VGND
port 614 nsew ground input
rlabel locali s 298660 173553 298799 173703 6 VGND
port 614 nsew ground input
rlabel locali s 1121 173369 1340 173519 6 VGND
port 614 nsew ground input
rlabel locali s 1104 173519 1340 173553 6 VGND
port 614 nsew ground input
rlabel locali s 1121 173553 1340 173703 6 VGND
port 614 nsew ground input
rlabel locali s 298695 173703 298799 173811 6 VGND
port 614 nsew ground input
rlabel locali s 1121 173703 1225 173811 6 VGND
port 614 nsew ground input
rlabel locali s 298695 174349 298799 174457 6 VGND
port 614 nsew ground input
rlabel locali s 1121 174349 1225 174457 6 VGND
port 614 nsew ground input
rlabel locali s 298660 174457 298799 174607 6 VGND
port 614 nsew ground input
rlabel locali s 298660 174607 298816 174641 6 VGND
port 614 nsew ground input
rlabel locali s 298660 174641 298799 174791 6 VGND
port 614 nsew ground input
rlabel locali s 1121 174457 1340 174607 6 VGND
port 614 nsew ground input
rlabel locali s 1104 174607 1340 174641 6 VGND
port 614 nsew ground input
rlabel locali s 1121 174641 1340 174791 6 VGND
port 614 nsew ground input
rlabel locali s 298695 174791 298799 174899 6 VGND
port 614 nsew ground input
rlabel locali s 1121 174791 1225 174899 6 VGND
port 614 nsew ground input
rlabel locali s 298695 175437 298799 175545 6 VGND
port 614 nsew ground input
rlabel locali s 1121 175437 1225 175545 6 VGND
port 614 nsew ground input
rlabel locali s 298660 175545 298799 175695 6 VGND
port 614 nsew ground input
rlabel locali s 298660 175695 298816 175729 6 VGND
port 614 nsew ground input
rlabel locali s 298660 175729 298799 175879 6 VGND
port 614 nsew ground input
rlabel locali s 1121 175545 1340 175695 6 VGND
port 614 nsew ground input
rlabel locali s 1104 175695 1340 175729 6 VGND
port 614 nsew ground input
rlabel locali s 1121 175729 1340 175879 6 VGND
port 614 nsew ground input
rlabel locali s 298695 175879 298799 175987 6 VGND
port 614 nsew ground input
rlabel locali s 1121 175879 1225 175987 6 VGND
port 614 nsew ground input
rlabel locali s 298695 176525 298799 176633 6 VGND
port 614 nsew ground input
rlabel locali s 1121 176525 1225 176633 6 VGND
port 614 nsew ground input
rlabel locali s 298660 176633 298799 176783 6 VGND
port 614 nsew ground input
rlabel locali s 298660 176783 298816 176817 6 VGND
port 614 nsew ground input
rlabel locali s 298660 176817 298799 176967 6 VGND
port 614 nsew ground input
rlabel locali s 1121 176633 1340 176783 6 VGND
port 614 nsew ground input
rlabel locali s 1104 176783 1340 176817 6 VGND
port 614 nsew ground input
rlabel locali s 1121 176817 1340 176967 6 VGND
port 614 nsew ground input
rlabel locali s 298695 176967 298799 177075 6 VGND
port 614 nsew ground input
rlabel locali s 1121 176967 1225 177075 6 VGND
port 614 nsew ground input
rlabel locali s 298695 177613 298799 177721 6 VGND
port 614 nsew ground input
rlabel locali s 1121 177613 1225 177721 6 VGND
port 614 nsew ground input
rlabel locali s 298660 177721 298799 177871 6 VGND
port 614 nsew ground input
rlabel locali s 298660 177871 298816 177905 6 VGND
port 614 nsew ground input
rlabel locali s 298660 177905 298799 178055 6 VGND
port 614 nsew ground input
rlabel locali s 1121 177721 1340 177871 6 VGND
port 614 nsew ground input
rlabel locali s 1104 177871 1340 177905 6 VGND
port 614 nsew ground input
rlabel locali s 1121 177905 1340 178055 6 VGND
port 614 nsew ground input
rlabel locali s 298695 178055 298799 178163 6 VGND
port 614 nsew ground input
rlabel locali s 1121 178055 1225 178163 6 VGND
port 614 nsew ground input
rlabel locali s 298695 178701 298799 178809 6 VGND
port 614 nsew ground input
rlabel locali s 1121 178701 1225 178809 6 VGND
port 614 nsew ground input
rlabel locali s 298660 178809 298799 178959 6 VGND
port 614 nsew ground input
rlabel locali s 298660 178959 298816 178993 6 VGND
port 614 nsew ground input
rlabel locali s 298660 178993 298799 179143 6 VGND
port 614 nsew ground input
rlabel locali s 1121 178809 1340 178959 6 VGND
port 614 nsew ground input
rlabel locali s 1104 178959 1340 178993 6 VGND
port 614 nsew ground input
rlabel locali s 1121 178993 1340 179143 6 VGND
port 614 nsew ground input
rlabel locali s 298695 179143 298799 179251 6 VGND
port 614 nsew ground input
rlabel locali s 1121 179143 1225 179251 6 VGND
port 614 nsew ground input
rlabel locali s 298695 179789 298799 179897 6 VGND
port 614 nsew ground input
rlabel locali s 1121 179789 1225 179897 6 VGND
port 614 nsew ground input
rlabel locali s 298660 179897 298799 180047 6 VGND
port 614 nsew ground input
rlabel locali s 298660 180047 298816 180081 6 VGND
port 614 nsew ground input
rlabel locali s 298660 180081 298799 180231 6 VGND
port 614 nsew ground input
rlabel locali s 1121 179897 1340 180047 6 VGND
port 614 nsew ground input
rlabel locali s 1104 180047 1340 180081 6 VGND
port 614 nsew ground input
rlabel locali s 1121 180081 1340 180231 6 VGND
port 614 nsew ground input
rlabel locali s 298695 180231 298799 180339 6 VGND
port 614 nsew ground input
rlabel locali s 1121 180231 1225 180339 6 VGND
port 614 nsew ground input
rlabel locali s 298695 180877 298799 180985 6 VGND
port 614 nsew ground input
rlabel locali s 1121 180877 1225 180985 6 VGND
port 614 nsew ground input
rlabel locali s 298660 180985 298799 181135 6 VGND
port 614 nsew ground input
rlabel locali s 298660 181135 298816 181169 6 VGND
port 614 nsew ground input
rlabel locali s 298660 181169 298799 181319 6 VGND
port 614 nsew ground input
rlabel locali s 1121 180985 1340 181135 6 VGND
port 614 nsew ground input
rlabel locali s 1104 181135 1340 181169 6 VGND
port 614 nsew ground input
rlabel locali s 1121 181169 1340 181319 6 VGND
port 614 nsew ground input
rlabel locali s 298695 181319 298799 181427 6 VGND
port 614 nsew ground input
rlabel locali s 1121 181319 1225 181427 6 VGND
port 614 nsew ground input
rlabel locali s 298695 181965 298799 182073 6 VGND
port 614 nsew ground input
rlabel locali s 1121 181965 1225 182073 6 VGND
port 614 nsew ground input
rlabel locali s 298660 182073 298799 182223 6 VGND
port 614 nsew ground input
rlabel locali s 298660 182223 298816 182257 6 VGND
port 614 nsew ground input
rlabel locali s 298660 182257 298799 182407 6 VGND
port 614 nsew ground input
rlabel locali s 1121 182073 1340 182223 6 VGND
port 614 nsew ground input
rlabel locali s 1104 182223 1340 182257 6 VGND
port 614 nsew ground input
rlabel locali s 1121 182257 1340 182407 6 VGND
port 614 nsew ground input
rlabel locali s 298695 182407 298799 182515 6 VGND
port 614 nsew ground input
rlabel locali s 1121 182407 1225 182515 6 VGND
port 614 nsew ground input
rlabel locali s 298695 183053 298799 183161 6 VGND
port 614 nsew ground input
rlabel locali s 1121 183053 1225 183161 6 VGND
port 614 nsew ground input
rlabel locali s 298660 183161 298799 183311 6 VGND
port 614 nsew ground input
rlabel locali s 298660 183311 298816 183345 6 VGND
port 614 nsew ground input
rlabel locali s 298660 183345 298799 183495 6 VGND
port 614 nsew ground input
rlabel locali s 1121 183161 1340 183311 6 VGND
port 614 nsew ground input
rlabel locali s 1104 183311 1340 183345 6 VGND
port 614 nsew ground input
rlabel locali s 1121 183345 1340 183495 6 VGND
port 614 nsew ground input
rlabel locali s 298695 183495 298799 183603 6 VGND
port 614 nsew ground input
rlabel locali s 1121 183495 1225 183603 6 VGND
port 614 nsew ground input
rlabel locali s 298695 184141 298799 184249 6 VGND
port 614 nsew ground input
rlabel locali s 1121 184141 1225 184249 6 VGND
port 614 nsew ground input
rlabel locali s 298660 184249 298799 184399 6 VGND
port 614 nsew ground input
rlabel locali s 298660 184399 298816 184433 6 VGND
port 614 nsew ground input
rlabel locali s 298660 184433 298799 184583 6 VGND
port 614 nsew ground input
rlabel locali s 1121 184249 1340 184399 6 VGND
port 614 nsew ground input
rlabel locali s 1104 184399 1340 184433 6 VGND
port 614 nsew ground input
rlabel locali s 1121 184433 1340 184583 6 VGND
port 614 nsew ground input
rlabel locali s 298695 184583 298799 184691 6 VGND
port 614 nsew ground input
rlabel locali s 1121 184583 1225 184691 6 VGND
port 614 nsew ground input
rlabel locali s 298695 185229 298799 185337 6 VGND
port 614 nsew ground input
rlabel locali s 1121 185229 1225 185337 6 VGND
port 614 nsew ground input
rlabel locali s 298660 185337 298799 185487 6 VGND
port 614 nsew ground input
rlabel locali s 298660 185487 298816 185521 6 VGND
port 614 nsew ground input
rlabel locali s 298660 185521 298799 185671 6 VGND
port 614 nsew ground input
rlabel locali s 1121 185337 1340 185487 6 VGND
port 614 nsew ground input
rlabel locali s 1104 185487 1340 185521 6 VGND
port 614 nsew ground input
rlabel locali s 1121 185521 1340 185671 6 VGND
port 614 nsew ground input
rlabel locali s 298695 185671 298799 185779 6 VGND
port 614 nsew ground input
rlabel locali s 1121 185671 1225 185779 6 VGND
port 614 nsew ground input
rlabel locali s 298695 186317 298799 186425 6 VGND
port 614 nsew ground input
rlabel locali s 1121 186317 1225 186425 6 VGND
port 614 nsew ground input
rlabel locali s 298660 186425 298799 186575 6 VGND
port 614 nsew ground input
rlabel locali s 298660 186575 298816 186609 6 VGND
port 614 nsew ground input
rlabel locali s 298660 186609 298799 186759 6 VGND
port 614 nsew ground input
rlabel locali s 1121 186425 1340 186575 6 VGND
port 614 nsew ground input
rlabel locali s 1104 186575 1340 186609 6 VGND
port 614 nsew ground input
rlabel locali s 1121 186609 1340 186759 6 VGND
port 614 nsew ground input
rlabel locali s 298695 186759 298799 186867 6 VGND
port 614 nsew ground input
rlabel locali s 1121 186759 1225 186867 6 VGND
port 614 nsew ground input
rlabel locali s 298695 187405 298799 187513 6 VGND
port 614 nsew ground input
rlabel locali s 1121 187405 1225 187513 6 VGND
port 614 nsew ground input
rlabel locali s 298660 187513 298799 187663 6 VGND
port 614 nsew ground input
rlabel locali s 298660 187663 298816 187697 6 VGND
port 614 nsew ground input
rlabel locali s 298660 187697 298799 187847 6 VGND
port 614 nsew ground input
rlabel locali s 1121 187513 1340 187663 6 VGND
port 614 nsew ground input
rlabel locali s 1104 187663 1340 187697 6 VGND
port 614 nsew ground input
rlabel locali s 1121 187697 1340 187847 6 VGND
port 614 nsew ground input
rlabel locali s 298695 187847 298799 187955 6 VGND
port 614 nsew ground input
rlabel locali s 1121 187847 1225 187955 6 VGND
port 614 nsew ground input
rlabel locali s 298695 188493 298799 188601 6 VGND
port 614 nsew ground input
rlabel locali s 1121 188493 1225 188601 6 VGND
port 614 nsew ground input
rlabel locali s 298660 188601 298799 188751 6 VGND
port 614 nsew ground input
rlabel locali s 298660 188751 298816 188785 6 VGND
port 614 nsew ground input
rlabel locali s 298660 188785 298799 188935 6 VGND
port 614 nsew ground input
rlabel locali s 1121 188601 1340 188751 6 VGND
port 614 nsew ground input
rlabel locali s 1104 188751 1340 188785 6 VGND
port 614 nsew ground input
rlabel locali s 1121 188785 1340 188935 6 VGND
port 614 nsew ground input
rlabel locali s 298695 188935 298799 189043 6 VGND
port 614 nsew ground input
rlabel locali s 1121 188935 1225 189043 6 VGND
port 614 nsew ground input
rlabel locali s 298695 189581 298799 189689 6 VGND
port 614 nsew ground input
rlabel locali s 1121 189581 1225 189689 6 VGND
port 614 nsew ground input
rlabel locali s 298660 189689 298799 189839 6 VGND
port 614 nsew ground input
rlabel locali s 298660 189839 298816 189873 6 VGND
port 614 nsew ground input
rlabel locali s 298660 189873 298799 190023 6 VGND
port 614 nsew ground input
rlabel locali s 1121 189689 1340 189839 6 VGND
port 614 nsew ground input
rlabel locali s 1104 189839 1340 189873 6 VGND
port 614 nsew ground input
rlabel locali s 1121 189873 1340 190023 6 VGND
port 614 nsew ground input
rlabel locali s 298695 190023 298799 190131 6 VGND
port 614 nsew ground input
rlabel locali s 1121 190023 1225 190131 6 VGND
port 614 nsew ground input
rlabel locali s 298695 190669 298799 190777 6 VGND
port 614 nsew ground input
rlabel locali s 1121 190669 1225 190777 6 VGND
port 614 nsew ground input
rlabel locali s 298660 190777 298799 190927 6 VGND
port 614 nsew ground input
rlabel locali s 298660 190927 298816 190961 6 VGND
port 614 nsew ground input
rlabel locali s 298660 190961 298799 191111 6 VGND
port 614 nsew ground input
rlabel locali s 1121 190777 1340 190927 6 VGND
port 614 nsew ground input
rlabel locali s 1104 190927 1340 190961 6 VGND
port 614 nsew ground input
rlabel locali s 1121 190961 1340 191111 6 VGND
port 614 nsew ground input
rlabel locali s 298695 191111 298799 191219 6 VGND
port 614 nsew ground input
rlabel locali s 1121 191111 1225 191219 6 VGND
port 614 nsew ground input
rlabel locali s 298695 191757 298799 191865 6 VGND
port 614 nsew ground input
rlabel locali s 1121 191757 1225 191865 6 VGND
port 614 nsew ground input
rlabel locali s 298660 191865 298799 192015 6 VGND
port 614 nsew ground input
rlabel locali s 298660 192015 298816 192049 6 VGND
port 614 nsew ground input
rlabel locali s 298660 192049 298799 192199 6 VGND
port 614 nsew ground input
rlabel locali s 1121 191865 1340 192015 6 VGND
port 614 nsew ground input
rlabel locali s 1104 192015 1340 192049 6 VGND
port 614 nsew ground input
rlabel locali s 1121 192049 1340 192199 6 VGND
port 614 nsew ground input
rlabel locali s 298695 192199 298799 192307 6 VGND
port 614 nsew ground input
rlabel locali s 1121 192199 1225 192307 6 VGND
port 614 nsew ground input
rlabel locali s 298695 192845 298799 192953 6 VGND
port 614 nsew ground input
rlabel locali s 1121 192845 1225 192953 6 VGND
port 614 nsew ground input
rlabel locali s 298660 192953 298799 193103 6 VGND
port 614 nsew ground input
rlabel locali s 298660 193103 298816 193137 6 VGND
port 614 nsew ground input
rlabel locali s 298660 193137 298799 193287 6 VGND
port 614 nsew ground input
rlabel locali s 1121 192953 1340 193103 6 VGND
port 614 nsew ground input
rlabel locali s 1104 193103 1340 193137 6 VGND
port 614 nsew ground input
rlabel locali s 1121 193137 1340 193287 6 VGND
port 614 nsew ground input
rlabel locali s 298695 193287 298799 193395 6 VGND
port 614 nsew ground input
rlabel locali s 1121 193287 1225 193395 6 VGND
port 614 nsew ground input
rlabel locali s 298695 193933 298799 194041 6 VGND
port 614 nsew ground input
rlabel locali s 1121 193933 1225 194041 6 VGND
port 614 nsew ground input
rlabel locali s 298660 194041 298799 194191 6 VGND
port 614 nsew ground input
rlabel locali s 298660 194191 298816 194225 6 VGND
port 614 nsew ground input
rlabel locali s 298660 194225 298799 194375 6 VGND
port 614 nsew ground input
rlabel locali s 1121 194041 1340 194191 6 VGND
port 614 nsew ground input
rlabel locali s 1104 194191 1340 194225 6 VGND
port 614 nsew ground input
rlabel locali s 1121 194225 1340 194375 6 VGND
port 614 nsew ground input
rlabel locali s 298695 194375 298799 194483 6 VGND
port 614 nsew ground input
rlabel locali s 1121 194375 1225 194483 6 VGND
port 614 nsew ground input
rlabel locali s 298695 195021 298799 195129 6 VGND
port 614 nsew ground input
rlabel locali s 1121 195021 1225 195129 6 VGND
port 614 nsew ground input
rlabel locali s 298660 195129 298799 195279 6 VGND
port 614 nsew ground input
rlabel locali s 298660 195279 298816 195313 6 VGND
port 614 nsew ground input
rlabel locali s 298660 195313 298799 195463 6 VGND
port 614 nsew ground input
rlabel locali s 1121 195129 1340 195279 6 VGND
port 614 nsew ground input
rlabel locali s 1104 195279 1340 195313 6 VGND
port 614 nsew ground input
rlabel locali s 1121 195313 1340 195463 6 VGND
port 614 nsew ground input
rlabel locali s 298695 195463 298799 195571 6 VGND
port 614 nsew ground input
rlabel locali s 1121 195463 1225 195571 6 VGND
port 614 nsew ground input
rlabel locali s 298695 196109 298799 196217 6 VGND
port 614 nsew ground input
rlabel locali s 1121 196109 1225 196217 6 VGND
port 614 nsew ground input
rlabel locali s 298660 196217 298799 196367 6 VGND
port 614 nsew ground input
rlabel locali s 298660 196367 298816 196401 6 VGND
port 614 nsew ground input
rlabel locali s 298660 196401 298799 196551 6 VGND
port 614 nsew ground input
rlabel locali s 1121 196217 1340 196367 6 VGND
port 614 nsew ground input
rlabel locali s 1104 196367 1340 196401 6 VGND
port 614 nsew ground input
rlabel locali s 1121 196401 1340 196551 6 VGND
port 614 nsew ground input
rlabel locali s 298695 196551 298799 196659 6 VGND
port 614 nsew ground input
rlabel locali s 1121 196551 1225 196659 6 VGND
port 614 nsew ground input
rlabel locali s 298695 197197 298799 197305 6 VGND
port 614 nsew ground input
rlabel locali s 1121 197197 1225 197305 6 VGND
port 614 nsew ground input
rlabel locali s 298660 197305 298799 197455 6 VGND
port 614 nsew ground input
rlabel locali s 298660 197455 298816 197489 6 VGND
port 614 nsew ground input
rlabel locali s 298660 197489 298799 197639 6 VGND
port 614 nsew ground input
rlabel locali s 1121 197305 1340 197455 6 VGND
port 614 nsew ground input
rlabel locali s 1104 197455 1340 197489 6 VGND
port 614 nsew ground input
rlabel locali s 1121 197489 1340 197639 6 VGND
port 614 nsew ground input
rlabel locali s 298695 197639 298799 197747 6 VGND
port 614 nsew ground input
rlabel locali s 1121 197639 1225 197747 6 VGND
port 614 nsew ground input
rlabel locali s 298695 198285 298799 198393 6 VGND
port 614 nsew ground input
rlabel locali s 1121 198285 1225 198393 6 VGND
port 614 nsew ground input
rlabel locali s 298660 198393 298799 198543 6 VGND
port 614 nsew ground input
rlabel locali s 298660 198543 298816 198577 6 VGND
port 614 nsew ground input
rlabel locali s 298660 198577 298799 198727 6 VGND
port 614 nsew ground input
rlabel locali s 1121 198393 1340 198543 6 VGND
port 614 nsew ground input
rlabel locali s 1104 198543 1340 198577 6 VGND
port 614 nsew ground input
rlabel locali s 1121 198577 1340 198727 6 VGND
port 614 nsew ground input
rlabel locali s 298695 198727 298799 198835 6 VGND
port 614 nsew ground input
rlabel locali s 1121 198727 1225 198835 6 VGND
port 614 nsew ground input
rlabel locali s 298695 199373 298799 199481 6 VGND
port 614 nsew ground input
rlabel locali s 1121 199373 1225 199481 6 VGND
port 614 nsew ground input
rlabel locali s 298660 199481 298799 199631 6 VGND
port 614 nsew ground input
rlabel locali s 298660 199631 298816 199665 6 VGND
port 614 nsew ground input
rlabel locali s 298660 199665 298799 199815 6 VGND
port 614 nsew ground input
rlabel locali s 1121 199481 1340 199631 6 VGND
port 614 nsew ground input
rlabel locali s 1104 199631 1340 199665 6 VGND
port 614 nsew ground input
rlabel locali s 1121 199665 1340 199815 6 VGND
port 614 nsew ground input
rlabel locali s 298695 199815 298799 199923 6 VGND
port 614 nsew ground input
rlabel locali s 1121 199815 1225 199923 6 VGND
port 614 nsew ground input
rlabel locali s 298695 200461 298799 200569 6 VGND
port 614 nsew ground input
rlabel locali s 1121 200461 1225 200569 6 VGND
port 614 nsew ground input
rlabel locali s 298660 200569 298799 200719 6 VGND
port 614 nsew ground input
rlabel locali s 298660 200719 298816 200753 6 VGND
port 614 nsew ground input
rlabel locali s 298660 200753 298799 200903 6 VGND
port 614 nsew ground input
rlabel locali s 1121 200569 1340 200719 6 VGND
port 614 nsew ground input
rlabel locali s 1104 200719 1340 200753 6 VGND
port 614 nsew ground input
rlabel locali s 1121 200753 1340 200903 6 VGND
port 614 nsew ground input
rlabel locali s 298695 200903 298799 201011 6 VGND
port 614 nsew ground input
rlabel locali s 1121 200903 1225 201011 6 VGND
port 614 nsew ground input
rlabel locali s 298695 201549 298799 201657 6 VGND
port 614 nsew ground input
rlabel locali s 1121 201549 1225 201657 6 VGND
port 614 nsew ground input
rlabel locali s 298660 201657 298799 201807 6 VGND
port 614 nsew ground input
rlabel locali s 298660 201807 298816 201841 6 VGND
port 614 nsew ground input
rlabel locali s 298660 201841 298799 201991 6 VGND
port 614 nsew ground input
rlabel locali s 1121 201657 1340 201807 6 VGND
port 614 nsew ground input
rlabel locali s 1104 201807 1340 201841 6 VGND
port 614 nsew ground input
rlabel locali s 1121 201841 1340 201991 6 VGND
port 614 nsew ground input
rlabel locali s 298695 201991 298799 202099 6 VGND
port 614 nsew ground input
rlabel locali s 1121 201991 1225 202099 6 VGND
port 614 nsew ground input
rlabel locali s 298695 202637 298799 202745 6 VGND
port 614 nsew ground input
rlabel locali s 1121 202637 1225 202745 6 VGND
port 614 nsew ground input
rlabel locali s 298660 202745 298799 202895 6 VGND
port 614 nsew ground input
rlabel locali s 298660 202895 298816 202929 6 VGND
port 614 nsew ground input
rlabel locali s 298660 202929 298799 203079 6 VGND
port 614 nsew ground input
rlabel locali s 1121 202745 1340 202895 6 VGND
port 614 nsew ground input
rlabel locali s 1104 202895 1340 202929 6 VGND
port 614 nsew ground input
rlabel locali s 1121 202929 1340 203079 6 VGND
port 614 nsew ground input
rlabel locali s 298695 203079 298799 203187 6 VGND
port 614 nsew ground input
rlabel locali s 1121 203079 1225 203187 6 VGND
port 614 nsew ground input
rlabel locali s 298695 203725 298799 203833 6 VGND
port 614 nsew ground input
rlabel locali s 1121 203725 1225 203833 6 VGND
port 614 nsew ground input
rlabel locali s 298660 203833 298799 203983 6 VGND
port 614 nsew ground input
rlabel locali s 298660 203983 298816 204017 6 VGND
port 614 nsew ground input
rlabel locali s 298660 204017 298799 204167 6 VGND
port 614 nsew ground input
rlabel locali s 1121 203833 1340 203983 6 VGND
port 614 nsew ground input
rlabel locali s 1104 203983 1340 204017 6 VGND
port 614 nsew ground input
rlabel locali s 1121 204017 1340 204167 6 VGND
port 614 nsew ground input
rlabel locali s 298695 204167 298799 204275 6 VGND
port 614 nsew ground input
rlabel locali s 1121 204167 1225 204275 6 VGND
port 614 nsew ground input
rlabel locali s 298695 204813 298799 204921 6 VGND
port 614 nsew ground input
rlabel locali s 1121 204813 1225 204921 6 VGND
port 614 nsew ground input
rlabel locali s 298660 204921 298799 205071 6 VGND
port 614 nsew ground input
rlabel locali s 298660 205071 298816 205105 6 VGND
port 614 nsew ground input
rlabel locali s 298660 205105 298799 205255 6 VGND
port 614 nsew ground input
rlabel locali s 1121 204921 1340 205071 6 VGND
port 614 nsew ground input
rlabel locali s 1104 205071 1340 205105 6 VGND
port 614 nsew ground input
rlabel locali s 1121 205105 1340 205255 6 VGND
port 614 nsew ground input
rlabel locali s 298695 205255 298799 205363 6 VGND
port 614 nsew ground input
rlabel locali s 1121 205255 1225 205363 6 VGND
port 614 nsew ground input
rlabel locali s 298695 205901 298799 206009 6 VGND
port 614 nsew ground input
rlabel locali s 1121 205901 1225 206009 6 VGND
port 614 nsew ground input
rlabel locali s 298660 206009 298799 206159 6 VGND
port 614 nsew ground input
rlabel locali s 298660 206159 298816 206193 6 VGND
port 614 nsew ground input
rlabel locali s 298660 206193 298799 206343 6 VGND
port 614 nsew ground input
rlabel locali s 1121 206009 1340 206159 6 VGND
port 614 nsew ground input
rlabel locali s 1104 206159 1340 206193 6 VGND
port 614 nsew ground input
rlabel locali s 1121 206193 1340 206343 6 VGND
port 614 nsew ground input
rlabel locali s 298695 206343 298799 206451 6 VGND
port 614 nsew ground input
rlabel locali s 1121 206343 1225 206451 6 VGND
port 614 nsew ground input
rlabel locali s 298695 206989 298799 207097 6 VGND
port 614 nsew ground input
rlabel locali s 1121 206989 1225 207097 6 VGND
port 614 nsew ground input
rlabel locali s 298660 207097 298799 207247 6 VGND
port 614 nsew ground input
rlabel locali s 298660 207247 298816 207281 6 VGND
port 614 nsew ground input
rlabel locali s 298660 207281 298799 207431 6 VGND
port 614 nsew ground input
rlabel locali s 1121 207097 1340 207247 6 VGND
port 614 nsew ground input
rlabel locali s 1104 207247 1340 207281 6 VGND
port 614 nsew ground input
rlabel locali s 1121 207281 1340 207431 6 VGND
port 614 nsew ground input
rlabel locali s 298695 207431 298799 207539 6 VGND
port 614 nsew ground input
rlabel locali s 1121 207431 1225 207539 6 VGND
port 614 nsew ground input
rlabel locali s 298695 208077 298799 208185 6 VGND
port 614 nsew ground input
rlabel locali s 1121 208077 1225 208185 6 VGND
port 614 nsew ground input
rlabel locali s 298660 208185 298799 208335 6 VGND
port 614 nsew ground input
rlabel locali s 298660 208335 298816 208369 6 VGND
port 614 nsew ground input
rlabel locali s 298660 208369 298799 208519 6 VGND
port 614 nsew ground input
rlabel locali s 1121 208185 1340 208335 6 VGND
port 614 nsew ground input
rlabel locali s 1104 208335 1340 208369 6 VGND
port 614 nsew ground input
rlabel locali s 1121 208369 1340 208519 6 VGND
port 614 nsew ground input
rlabel locali s 298695 208519 298799 208627 6 VGND
port 614 nsew ground input
rlabel locali s 1121 208519 1225 208627 6 VGND
port 614 nsew ground input
rlabel locali s 298695 209165 298799 209273 6 VGND
port 614 nsew ground input
rlabel locali s 1121 209165 1225 209273 6 VGND
port 614 nsew ground input
rlabel locali s 298660 209273 298799 209423 6 VGND
port 614 nsew ground input
rlabel locali s 298660 209423 298816 209457 6 VGND
port 614 nsew ground input
rlabel locali s 298660 209457 298799 209607 6 VGND
port 614 nsew ground input
rlabel locali s 1121 209273 1340 209423 6 VGND
port 614 nsew ground input
rlabel locali s 1104 209423 1340 209457 6 VGND
port 614 nsew ground input
rlabel locali s 1121 209457 1340 209607 6 VGND
port 614 nsew ground input
rlabel locali s 298695 209607 298799 209715 6 VGND
port 614 nsew ground input
rlabel locali s 1121 209607 1225 209715 6 VGND
port 614 nsew ground input
rlabel locali s 298695 210253 298799 210361 6 VGND
port 614 nsew ground input
rlabel locali s 1121 210253 1225 210361 6 VGND
port 614 nsew ground input
rlabel locali s 298660 210361 298799 210511 6 VGND
port 614 nsew ground input
rlabel locali s 298660 210511 298816 210545 6 VGND
port 614 nsew ground input
rlabel locali s 298660 210545 298799 210695 6 VGND
port 614 nsew ground input
rlabel locali s 1121 210361 1340 210511 6 VGND
port 614 nsew ground input
rlabel locali s 1104 210511 1340 210545 6 VGND
port 614 nsew ground input
rlabel locali s 1121 210545 1340 210695 6 VGND
port 614 nsew ground input
rlabel locali s 298695 210695 298799 210803 6 VGND
port 614 nsew ground input
rlabel locali s 1121 210695 1225 210803 6 VGND
port 614 nsew ground input
rlabel locali s 298695 211341 298799 211449 6 VGND
port 614 nsew ground input
rlabel locali s 1121 211341 1225 211449 6 VGND
port 614 nsew ground input
rlabel locali s 298660 211449 298799 211599 6 VGND
port 614 nsew ground input
rlabel locali s 298660 211599 298816 211633 6 VGND
port 614 nsew ground input
rlabel locali s 298660 211633 298799 211783 6 VGND
port 614 nsew ground input
rlabel locali s 1121 211449 1340 211599 6 VGND
port 614 nsew ground input
rlabel locali s 1104 211599 1340 211633 6 VGND
port 614 nsew ground input
rlabel locali s 1121 211633 1340 211783 6 VGND
port 614 nsew ground input
rlabel locali s 298695 211783 298799 211891 6 VGND
port 614 nsew ground input
rlabel locali s 1121 211783 1225 211891 6 VGND
port 614 nsew ground input
rlabel locali s 298695 212429 298799 212537 6 VGND
port 614 nsew ground input
rlabel locali s 1121 212429 1225 212537 6 VGND
port 614 nsew ground input
rlabel locali s 298660 212537 298799 212687 6 VGND
port 614 nsew ground input
rlabel locali s 298660 212687 298816 212721 6 VGND
port 614 nsew ground input
rlabel locali s 298660 212721 298799 212871 6 VGND
port 614 nsew ground input
rlabel locali s 1121 212537 1340 212687 6 VGND
port 614 nsew ground input
rlabel locali s 1104 212687 1340 212721 6 VGND
port 614 nsew ground input
rlabel locali s 1121 212721 1340 212871 6 VGND
port 614 nsew ground input
rlabel locali s 298695 212871 298799 212979 6 VGND
port 614 nsew ground input
rlabel locali s 1121 212871 1225 212979 6 VGND
port 614 nsew ground input
rlabel locali s 298695 213517 298799 213625 6 VGND
port 614 nsew ground input
rlabel locali s 1121 213517 1225 213625 6 VGND
port 614 nsew ground input
rlabel locali s 298660 213625 298799 213775 6 VGND
port 614 nsew ground input
rlabel locali s 298660 213775 298816 213809 6 VGND
port 614 nsew ground input
rlabel locali s 298660 213809 298799 213959 6 VGND
port 614 nsew ground input
rlabel locali s 1121 213625 1340 213775 6 VGND
port 614 nsew ground input
rlabel locali s 1104 213775 1340 213809 6 VGND
port 614 nsew ground input
rlabel locali s 1121 213809 1340 213959 6 VGND
port 614 nsew ground input
rlabel locali s 298695 213959 298799 214067 6 VGND
port 614 nsew ground input
rlabel locali s 1121 213959 1225 214067 6 VGND
port 614 nsew ground input
rlabel locali s 298695 214605 298799 214713 6 VGND
port 614 nsew ground input
rlabel locali s 1121 214605 1225 214713 6 VGND
port 614 nsew ground input
rlabel locali s 298660 214713 298799 214863 6 VGND
port 614 nsew ground input
rlabel locali s 298660 214863 298816 214897 6 VGND
port 614 nsew ground input
rlabel locali s 298660 214897 298799 215047 6 VGND
port 614 nsew ground input
rlabel locali s 1121 214713 1340 214863 6 VGND
port 614 nsew ground input
rlabel locali s 1104 214863 1340 214897 6 VGND
port 614 nsew ground input
rlabel locali s 1121 214897 1340 215047 6 VGND
port 614 nsew ground input
rlabel locali s 298695 215047 298799 215155 6 VGND
port 614 nsew ground input
rlabel locali s 1121 215047 1225 215155 6 VGND
port 614 nsew ground input
rlabel locali s 298695 215693 298799 215801 6 VGND
port 614 nsew ground input
rlabel locali s 1121 215693 1225 215801 6 VGND
port 614 nsew ground input
rlabel locali s 298660 215801 298799 215951 6 VGND
port 614 nsew ground input
rlabel locali s 298660 215951 298816 215985 6 VGND
port 614 nsew ground input
rlabel locali s 298660 215985 298799 216135 6 VGND
port 614 nsew ground input
rlabel locali s 1121 215801 1340 215951 6 VGND
port 614 nsew ground input
rlabel locali s 1104 215951 1340 215985 6 VGND
port 614 nsew ground input
rlabel locali s 1121 215985 1340 216135 6 VGND
port 614 nsew ground input
rlabel locali s 298695 216135 298799 216243 6 VGND
port 614 nsew ground input
rlabel locali s 1121 216135 1225 216243 6 VGND
port 614 nsew ground input
rlabel locali s 298695 216781 298799 216889 6 VGND
port 614 nsew ground input
rlabel locali s 1121 216781 1225 216889 6 VGND
port 614 nsew ground input
rlabel locali s 298660 216889 298799 217039 6 VGND
port 614 nsew ground input
rlabel locali s 298660 217039 298816 217073 6 VGND
port 614 nsew ground input
rlabel locali s 298660 217073 298799 217223 6 VGND
port 614 nsew ground input
rlabel locali s 1121 216889 1340 217039 6 VGND
port 614 nsew ground input
rlabel locali s 1104 217039 1340 217073 6 VGND
port 614 nsew ground input
rlabel locali s 1121 217073 1340 217223 6 VGND
port 614 nsew ground input
rlabel locali s 298695 217223 298799 217331 6 VGND
port 614 nsew ground input
rlabel locali s 1121 217223 1225 217331 6 VGND
port 614 nsew ground input
rlabel locali s 298695 217869 298799 217977 6 VGND
port 614 nsew ground input
rlabel locali s 1121 217869 1225 217977 6 VGND
port 614 nsew ground input
rlabel locali s 298660 217977 298799 218127 6 VGND
port 614 nsew ground input
rlabel locali s 298660 218127 298816 218161 6 VGND
port 614 nsew ground input
rlabel locali s 298660 218161 298799 218311 6 VGND
port 614 nsew ground input
rlabel locali s 1121 217977 1340 218127 6 VGND
port 614 nsew ground input
rlabel locali s 1104 218127 1340 218161 6 VGND
port 614 nsew ground input
rlabel locali s 1121 218161 1340 218311 6 VGND
port 614 nsew ground input
rlabel locali s 298695 218311 298799 218419 6 VGND
port 614 nsew ground input
rlabel locali s 1121 218311 1225 218419 6 VGND
port 614 nsew ground input
rlabel locali s 298695 218957 298799 219065 6 VGND
port 614 nsew ground input
rlabel locali s 1121 218957 1225 219065 6 VGND
port 614 nsew ground input
rlabel locali s 298660 219065 298799 219215 6 VGND
port 614 nsew ground input
rlabel locali s 298660 219215 298816 219249 6 VGND
port 614 nsew ground input
rlabel locali s 298660 219249 298799 219399 6 VGND
port 614 nsew ground input
rlabel locali s 1121 219065 1340 219215 6 VGND
port 614 nsew ground input
rlabel locali s 1104 219215 1340 219249 6 VGND
port 614 nsew ground input
rlabel locali s 1121 219249 1340 219399 6 VGND
port 614 nsew ground input
rlabel locali s 298695 219399 298799 219507 6 VGND
port 614 nsew ground input
rlabel locali s 1121 219399 1225 219507 6 VGND
port 614 nsew ground input
rlabel locali s 298695 220045 298799 220153 6 VGND
port 614 nsew ground input
rlabel locali s 1121 220045 1225 220153 6 VGND
port 614 nsew ground input
rlabel locali s 298660 220153 298799 220303 6 VGND
port 614 nsew ground input
rlabel locali s 298660 220303 298816 220337 6 VGND
port 614 nsew ground input
rlabel locali s 298660 220337 298799 220487 6 VGND
port 614 nsew ground input
rlabel locali s 1121 220153 1340 220303 6 VGND
port 614 nsew ground input
rlabel locali s 1104 220303 1340 220337 6 VGND
port 614 nsew ground input
rlabel locali s 1121 220337 1340 220487 6 VGND
port 614 nsew ground input
rlabel locali s 298695 220487 298799 220595 6 VGND
port 614 nsew ground input
rlabel locali s 1121 220487 1225 220595 6 VGND
port 614 nsew ground input
rlabel locali s 298695 221133 298799 221241 6 VGND
port 614 nsew ground input
rlabel locali s 1121 221133 1225 221241 6 VGND
port 614 nsew ground input
rlabel locali s 298660 221241 298799 221391 6 VGND
port 614 nsew ground input
rlabel locali s 298660 221391 298816 221425 6 VGND
port 614 nsew ground input
rlabel locali s 298660 221425 298799 221575 6 VGND
port 614 nsew ground input
rlabel locali s 1121 221241 1340 221391 6 VGND
port 614 nsew ground input
rlabel locali s 1104 221391 1340 221425 6 VGND
port 614 nsew ground input
rlabel locali s 1121 221425 1340 221575 6 VGND
port 614 nsew ground input
rlabel locali s 298695 221575 298799 221683 6 VGND
port 614 nsew ground input
rlabel locali s 1121 221575 1225 221683 6 VGND
port 614 nsew ground input
rlabel locali s 298695 222221 298799 222329 6 VGND
port 614 nsew ground input
rlabel locali s 1121 222221 1225 222329 6 VGND
port 614 nsew ground input
rlabel locali s 298660 222329 298799 222479 6 VGND
port 614 nsew ground input
rlabel locali s 298660 222479 298816 222513 6 VGND
port 614 nsew ground input
rlabel locali s 298660 222513 298799 222663 6 VGND
port 614 nsew ground input
rlabel locali s 1121 222329 1340 222479 6 VGND
port 614 nsew ground input
rlabel locali s 1104 222479 1340 222513 6 VGND
port 614 nsew ground input
rlabel locali s 1121 222513 1340 222663 6 VGND
port 614 nsew ground input
rlabel locali s 298695 222663 298799 222771 6 VGND
port 614 nsew ground input
rlabel locali s 1121 222663 1225 222771 6 VGND
port 614 nsew ground input
rlabel locali s 298695 223309 298799 223417 6 VGND
port 614 nsew ground input
rlabel locali s 1121 223309 1225 223417 6 VGND
port 614 nsew ground input
rlabel locali s 298660 223417 298799 223567 6 VGND
port 614 nsew ground input
rlabel locali s 298660 223567 298816 223601 6 VGND
port 614 nsew ground input
rlabel locali s 298660 223601 298799 223751 6 VGND
port 614 nsew ground input
rlabel locali s 1121 223417 1340 223567 6 VGND
port 614 nsew ground input
rlabel locali s 1104 223567 1340 223601 6 VGND
port 614 nsew ground input
rlabel locali s 1121 223601 1340 223751 6 VGND
port 614 nsew ground input
rlabel locali s 298695 223751 298799 223859 6 VGND
port 614 nsew ground input
rlabel locali s 1121 223751 1225 223859 6 VGND
port 614 nsew ground input
rlabel locali s 298695 224397 298799 224505 6 VGND
port 614 nsew ground input
rlabel locali s 1121 224397 1225 224505 6 VGND
port 614 nsew ground input
rlabel locali s 298660 224505 298799 224655 6 VGND
port 614 nsew ground input
rlabel locali s 298660 224655 298816 224689 6 VGND
port 614 nsew ground input
rlabel locali s 298660 224689 298799 224839 6 VGND
port 614 nsew ground input
rlabel locali s 1121 224505 1340 224655 6 VGND
port 614 nsew ground input
rlabel locali s 1104 224655 1340 224689 6 VGND
port 614 nsew ground input
rlabel locali s 1121 224689 1340 224839 6 VGND
port 614 nsew ground input
rlabel locali s 298695 224839 298799 224947 6 VGND
port 614 nsew ground input
rlabel locali s 1121 224839 1225 224947 6 VGND
port 614 nsew ground input
rlabel locali s 298695 225485 298799 225593 6 VGND
port 614 nsew ground input
rlabel locali s 1121 225485 1225 225593 6 VGND
port 614 nsew ground input
rlabel locali s 298660 225593 298799 225743 6 VGND
port 614 nsew ground input
rlabel locali s 298660 225743 298816 225777 6 VGND
port 614 nsew ground input
rlabel locali s 298660 225777 298799 225927 6 VGND
port 614 nsew ground input
rlabel locali s 1121 225593 1340 225743 6 VGND
port 614 nsew ground input
rlabel locali s 1104 225743 1340 225777 6 VGND
port 614 nsew ground input
rlabel locali s 1121 225777 1340 225927 6 VGND
port 614 nsew ground input
rlabel locali s 298695 225927 298799 226035 6 VGND
port 614 nsew ground input
rlabel locali s 1121 225927 1225 226035 6 VGND
port 614 nsew ground input
rlabel locali s 298695 226573 298799 226681 6 VGND
port 614 nsew ground input
rlabel locali s 1121 226573 1225 226681 6 VGND
port 614 nsew ground input
rlabel locali s 298660 226681 298799 226831 6 VGND
port 614 nsew ground input
rlabel locali s 298660 226831 298816 226865 6 VGND
port 614 nsew ground input
rlabel locali s 298660 226865 298799 227015 6 VGND
port 614 nsew ground input
rlabel locali s 1121 226681 1340 226831 6 VGND
port 614 nsew ground input
rlabel locali s 1104 226831 1340 226865 6 VGND
port 614 nsew ground input
rlabel locali s 1121 226865 1340 227015 6 VGND
port 614 nsew ground input
rlabel locali s 298695 227015 298799 227123 6 VGND
port 614 nsew ground input
rlabel locali s 1121 227015 1225 227123 6 VGND
port 614 nsew ground input
rlabel locali s 298695 227661 298799 227769 6 VGND
port 614 nsew ground input
rlabel locali s 1121 227661 1225 227769 6 VGND
port 614 nsew ground input
rlabel locali s 298660 227769 298799 227919 6 VGND
port 614 nsew ground input
rlabel locali s 298660 227919 298816 227953 6 VGND
port 614 nsew ground input
rlabel locali s 298660 227953 298799 228103 6 VGND
port 614 nsew ground input
rlabel locali s 1121 227769 1340 227919 6 VGND
port 614 nsew ground input
rlabel locali s 1104 227919 1340 227953 6 VGND
port 614 nsew ground input
rlabel locali s 1121 227953 1340 228103 6 VGND
port 614 nsew ground input
rlabel locali s 298695 228103 298799 228211 6 VGND
port 614 nsew ground input
rlabel locali s 1121 228103 1225 228211 6 VGND
port 614 nsew ground input
rlabel locali s 298695 228749 298799 228857 6 VGND
port 614 nsew ground input
rlabel locali s 1121 228749 1225 228857 6 VGND
port 614 nsew ground input
rlabel locali s 298660 228857 298799 229007 6 VGND
port 614 nsew ground input
rlabel locali s 298660 229007 298816 229041 6 VGND
port 614 nsew ground input
rlabel locali s 298660 229041 298799 229191 6 VGND
port 614 nsew ground input
rlabel locali s 1121 228857 1340 229007 6 VGND
port 614 nsew ground input
rlabel locali s 1104 229007 1340 229041 6 VGND
port 614 nsew ground input
rlabel locali s 1121 229041 1340 229191 6 VGND
port 614 nsew ground input
rlabel locali s 298695 229191 298799 229299 6 VGND
port 614 nsew ground input
rlabel locali s 1121 229191 1225 229299 6 VGND
port 614 nsew ground input
rlabel locali s 298695 229837 298799 229945 6 VGND
port 614 nsew ground input
rlabel locali s 1121 229837 1225 229945 6 VGND
port 614 nsew ground input
rlabel locali s 298660 229945 298799 230095 6 VGND
port 614 nsew ground input
rlabel locali s 298660 230095 298816 230129 6 VGND
port 614 nsew ground input
rlabel locali s 298660 230129 298799 230279 6 VGND
port 614 nsew ground input
rlabel locali s 1121 229945 1340 230095 6 VGND
port 614 nsew ground input
rlabel locali s 1104 230095 1340 230129 6 VGND
port 614 nsew ground input
rlabel locali s 1121 230129 1340 230279 6 VGND
port 614 nsew ground input
rlabel locali s 298695 230279 298799 230387 6 VGND
port 614 nsew ground input
rlabel locali s 1121 230279 1225 230387 6 VGND
port 614 nsew ground input
rlabel locali s 298695 230925 298799 231033 6 VGND
port 614 nsew ground input
rlabel locali s 1121 230925 1225 231033 6 VGND
port 614 nsew ground input
rlabel locali s 298660 231033 298799 231183 6 VGND
port 614 nsew ground input
rlabel locali s 298660 231183 298816 231217 6 VGND
port 614 nsew ground input
rlabel locali s 298660 231217 298799 231367 6 VGND
port 614 nsew ground input
rlabel locali s 1121 231033 1340 231183 6 VGND
port 614 nsew ground input
rlabel locali s 1104 231183 1340 231217 6 VGND
port 614 nsew ground input
rlabel locali s 1121 231217 1340 231367 6 VGND
port 614 nsew ground input
rlabel locali s 298695 231367 298799 231475 6 VGND
port 614 nsew ground input
rlabel locali s 1121 231367 1225 231475 6 VGND
port 614 nsew ground input
rlabel locali s 298695 232013 298799 232121 6 VGND
port 614 nsew ground input
rlabel locali s 1121 232013 1225 232121 6 VGND
port 614 nsew ground input
rlabel locali s 298660 232121 298799 232271 6 VGND
port 614 nsew ground input
rlabel locali s 298660 232271 298816 232305 6 VGND
port 614 nsew ground input
rlabel locali s 298660 232305 298799 232455 6 VGND
port 614 nsew ground input
rlabel locali s 1121 232121 1340 232271 6 VGND
port 614 nsew ground input
rlabel locali s 1104 232271 1340 232305 6 VGND
port 614 nsew ground input
rlabel locali s 1121 232305 1340 232455 6 VGND
port 614 nsew ground input
rlabel locali s 298695 232455 298799 232563 6 VGND
port 614 nsew ground input
rlabel locali s 1121 232455 1225 232563 6 VGND
port 614 nsew ground input
rlabel locali s 298695 233101 298799 233209 6 VGND
port 614 nsew ground input
rlabel locali s 1121 233101 1225 233209 6 VGND
port 614 nsew ground input
rlabel locali s 298660 233209 298799 233359 6 VGND
port 614 nsew ground input
rlabel locali s 298660 233359 298816 233393 6 VGND
port 614 nsew ground input
rlabel locali s 298660 233393 298799 233543 6 VGND
port 614 nsew ground input
rlabel locali s 1121 233209 1340 233359 6 VGND
port 614 nsew ground input
rlabel locali s 1104 233359 1340 233393 6 VGND
port 614 nsew ground input
rlabel locali s 1121 233393 1340 233543 6 VGND
port 614 nsew ground input
rlabel locali s 298695 233543 298799 233651 6 VGND
port 614 nsew ground input
rlabel locali s 1121 233543 1225 233651 6 VGND
port 614 nsew ground input
rlabel locali s 298695 234189 298799 234297 6 VGND
port 614 nsew ground input
rlabel locali s 1121 234189 1225 234297 6 VGND
port 614 nsew ground input
rlabel locali s 298660 234297 298799 234447 6 VGND
port 614 nsew ground input
rlabel locali s 298660 234447 298816 234481 6 VGND
port 614 nsew ground input
rlabel locali s 298660 234481 298799 234631 6 VGND
port 614 nsew ground input
rlabel locali s 1121 234297 1340 234447 6 VGND
port 614 nsew ground input
rlabel locali s 1104 234447 1340 234481 6 VGND
port 614 nsew ground input
rlabel locali s 1121 234481 1340 234631 6 VGND
port 614 nsew ground input
rlabel locali s 298695 234631 298799 234739 6 VGND
port 614 nsew ground input
rlabel locali s 1121 234631 1225 234739 6 VGND
port 614 nsew ground input
rlabel locali s 298695 235277 298799 235385 6 VGND
port 614 nsew ground input
rlabel locali s 1121 235277 1225 235385 6 VGND
port 614 nsew ground input
rlabel locali s 298660 235385 298799 235535 6 VGND
port 614 nsew ground input
rlabel locali s 298660 235535 298816 235569 6 VGND
port 614 nsew ground input
rlabel locali s 298660 235569 298799 235719 6 VGND
port 614 nsew ground input
rlabel locali s 1121 235385 1340 235535 6 VGND
port 614 nsew ground input
rlabel locali s 1104 235535 1340 235569 6 VGND
port 614 nsew ground input
rlabel locali s 1121 235569 1340 235719 6 VGND
port 614 nsew ground input
rlabel locali s 298695 235719 298799 235827 6 VGND
port 614 nsew ground input
rlabel locali s 1121 235719 1225 235827 6 VGND
port 614 nsew ground input
rlabel locali s 298695 236365 298799 236473 6 VGND
port 614 nsew ground input
rlabel locali s 1121 236365 1225 236473 6 VGND
port 614 nsew ground input
rlabel locali s 298660 236473 298799 236623 6 VGND
port 614 nsew ground input
rlabel locali s 298660 236623 298816 236657 6 VGND
port 614 nsew ground input
rlabel locali s 298660 236657 298799 236807 6 VGND
port 614 nsew ground input
rlabel locali s 1121 236473 1340 236623 6 VGND
port 614 nsew ground input
rlabel locali s 1104 236623 1340 236657 6 VGND
port 614 nsew ground input
rlabel locali s 1121 236657 1340 236807 6 VGND
port 614 nsew ground input
rlabel locali s 298695 236807 298799 236915 6 VGND
port 614 nsew ground input
rlabel locali s 1121 236807 1225 236915 6 VGND
port 614 nsew ground input
rlabel locali s 298695 237453 298799 237561 6 VGND
port 614 nsew ground input
rlabel locali s 1121 237453 1225 237561 6 VGND
port 614 nsew ground input
rlabel locali s 298660 237561 298799 237711 6 VGND
port 614 nsew ground input
rlabel locali s 298660 237711 298816 237745 6 VGND
port 614 nsew ground input
rlabel locali s 298660 237745 298799 237895 6 VGND
port 614 nsew ground input
rlabel locali s 1121 237561 1340 237711 6 VGND
port 614 nsew ground input
rlabel locali s 1104 237711 1340 237745 6 VGND
port 614 nsew ground input
rlabel locali s 1121 237745 1340 237895 6 VGND
port 614 nsew ground input
rlabel locali s 298695 237895 298799 238003 6 VGND
port 614 nsew ground input
rlabel locali s 1121 237895 1225 238003 6 VGND
port 614 nsew ground input
rlabel locali s 298695 238541 298799 238649 6 VGND
port 614 nsew ground input
rlabel locali s 1121 238541 1225 238649 6 VGND
port 614 nsew ground input
rlabel locali s 298660 238649 298799 238799 6 VGND
port 614 nsew ground input
rlabel locali s 298660 238799 298816 238833 6 VGND
port 614 nsew ground input
rlabel locali s 298660 238833 298799 238983 6 VGND
port 614 nsew ground input
rlabel locali s 1121 238649 1340 238799 6 VGND
port 614 nsew ground input
rlabel locali s 1104 238799 1340 238833 6 VGND
port 614 nsew ground input
rlabel locali s 1121 238833 1340 238983 6 VGND
port 614 nsew ground input
rlabel locali s 298695 238983 298799 239091 6 VGND
port 614 nsew ground input
rlabel locali s 1121 238983 1225 239091 6 VGND
port 614 nsew ground input
rlabel locali s 298695 239629 298799 239737 6 VGND
port 614 nsew ground input
rlabel locali s 1121 239629 1225 239737 6 VGND
port 614 nsew ground input
rlabel locali s 298660 239737 298799 239887 6 VGND
port 614 nsew ground input
rlabel locali s 298660 239887 298816 239921 6 VGND
port 614 nsew ground input
rlabel locali s 298660 239921 298799 240071 6 VGND
port 614 nsew ground input
rlabel locali s 1121 239737 1340 239887 6 VGND
port 614 nsew ground input
rlabel locali s 1104 239887 1340 239921 6 VGND
port 614 nsew ground input
rlabel locali s 1121 239921 1340 240071 6 VGND
port 614 nsew ground input
rlabel locali s 298695 240071 298799 240179 6 VGND
port 614 nsew ground input
rlabel locali s 1121 240071 1225 240179 6 VGND
port 614 nsew ground input
rlabel locali s 298695 240717 298799 240825 6 VGND
port 614 nsew ground input
rlabel locali s 1121 240717 1225 240825 6 VGND
port 614 nsew ground input
rlabel locali s 298660 240825 298799 240975 6 VGND
port 614 nsew ground input
rlabel locali s 298660 240975 298816 241009 6 VGND
port 614 nsew ground input
rlabel locali s 298660 241009 298799 241159 6 VGND
port 614 nsew ground input
rlabel locali s 1121 240825 1340 240975 6 VGND
port 614 nsew ground input
rlabel locali s 1104 240975 1340 241009 6 VGND
port 614 nsew ground input
rlabel locali s 1121 241009 1340 241159 6 VGND
port 614 nsew ground input
rlabel locali s 298695 241159 298799 241267 6 VGND
port 614 nsew ground input
rlabel locali s 1121 241159 1225 241267 6 VGND
port 614 nsew ground input
rlabel locali s 298695 241805 298799 241913 6 VGND
port 614 nsew ground input
rlabel locali s 1121 241805 1225 241913 6 VGND
port 614 nsew ground input
rlabel locali s 298660 241913 298799 242063 6 VGND
port 614 nsew ground input
rlabel locali s 298660 242063 298816 242097 6 VGND
port 614 nsew ground input
rlabel locali s 298660 242097 298799 242247 6 VGND
port 614 nsew ground input
rlabel locali s 1121 241913 1340 242063 6 VGND
port 614 nsew ground input
rlabel locali s 1104 242063 1340 242097 6 VGND
port 614 nsew ground input
rlabel locali s 1121 242097 1340 242247 6 VGND
port 614 nsew ground input
rlabel locali s 298695 242247 298799 242355 6 VGND
port 614 nsew ground input
rlabel locali s 1121 242247 1225 242355 6 VGND
port 614 nsew ground input
rlabel locali s 298695 242893 298799 243001 6 VGND
port 614 nsew ground input
rlabel locali s 1121 242893 1225 243001 6 VGND
port 614 nsew ground input
rlabel locali s 298660 243001 298799 243151 6 VGND
port 614 nsew ground input
rlabel locali s 298660 243151 298816 243185 6 VGND
port 614 nsew ground input
rlabel locali s 298660 243185 298799 243335 6 VGND
port 614 nsew ground input
rlabel locali s 1121 243001 1340 243151 6 VGND
port 614 nsew ground input
rlabel locali s 1104 243151 1340 243185 6 VGND
port 614 nsew ground input
rlabel locali s 1121 243185 1340 243335 6 VGND
port 614 nsew ground input
rlabel locali s 298695 243335 298799 243443 6 VGND
port 614 nsew ground input
rlabel locali s 1121 243335 1225 243443 6 VGND
port 614 nsew ground input
rlabel locali s 298695 243981 298799 244089 6 VGND
port 614 nsew ground input
rlabel locali s 1121 243981 1225 244089 6 VGND
port 614 nsew ground input
rlabel locali s 298660 244089 298799 244239 6 VGND
port 614 nsew ground input
rlabel locali s 298660 244239 298816 244273 6 VGND
port 614 nsew ground input
rlabel locali s 298660 244273 298799 244423 6 VGND
port 614 nsew ground input
rlabel locali s 1121 244089 1340 244239 6 VGND
port 614 nsew ground input
rlabel locali s 1104 244239 1340 244273 6 VGND
port 614 nsew ground input
rlabel locali s 1121 244273 1340 244423 6 VGND
port 614 nsew ground input
rlabel locali s 298695 244423 298799 244531 6 VGND
port 614 nsew ground input
rlabel locali s 1121 244423 1225 244531 6 VGND
port 614 nsew ground input
rlabel locali s 298695 245069 298799 245177 6 VGND
port 614 nsew ground input
rlabel locali s 1121 245069 1225 245177 6 VGND
port 614 nsew ground input
rlabel locali s 298660 245177 298799 245327 6 VGND
port 614 nsew ground input
rlabel locali s 298660 245327 298816 245361 6 VGND
port 614 nsew ground input
rlabel locali s 298660 245361 298799 245511 6 VGND
port 614 nsew ground input
rlabel locali s 1121 245177 1340 245327 6 VGND
port 614 nsew ground input
rlabel locali s 1104 245327 1340 245361 6 VGND
port 614 nsew ground input
rlabel locali s 1121 245361 1340 245511 6 VGND
port 614 nsew ground input
rlabel locali s 298695 245511 298799 245619 6 VGND
port 614 nsew ground input
rlabel locali s 1121 245511 1225 245619 6 VGND
port 614 nsew ground input
rlabel locali s 298695 246157 298799 246265 6 VGND
port 614 nsew ground input
rlabel locali s 1121 246157 1225 246265 6 VGND
port 614 nsew ground input
rlabel locali s 298660 246265 298799 246415 6 VGND
port 614 nsew ground input
rlabel locali s 298660 246415 298816 246449 6 VGND
port 614 nsew ground input
rlabel locali s 298660 246449 298799 246599 6 VGND
port 614 nsew ground input
rlabel locali s 1121 246265 1340 246415 6 VGND
port 614 nsew ground input
rlabel locali s 1104 246415 1340 246449 6 VGND
port 614 nsew ground input
rlabel locali s 1121 246449 1340 246599 6 VGND
port 614 nsew ground input
rlabel locali s 298695 246599 298799 246707 6 VGND
port 614 nsew ground input
rlabel locali s 1121 246599 1225 246707 6 VGND
port 614 nsew ground input
rlabel locali s 298695 247245 298799 247353 6 VGND
port 614 nsew ground input
rlabel locali s 1121 247245 1225 247353 6 VGND
port 614 nsew ground input
rlabel locali s 298660 247353 298799 247503 6 VGND
port 614 nsew ground input
rlabel locali s 298660 247503 298816 247537 6 VGND
port 614 nsew ground input
rlabel locali s 298660 247537 298799 247687 6 VGND
port 614 nsew ground input
rlabel locali s 1121 247353 1340 247503 6 VGND
port 614 nsew ground input
rlabel locali s 1104 247503 1340 247537 6 VGND
port 614 nsew ground input
rlabel locali s 1121 247537 1340 247687 6 VGND
port 614 nsew ground input
rlabel locali s 298695 247687 298799 247795 6 VGND
port 614 nsew ground input
rlabel locali s 1121 247687 1225 247795 6 VGND
port 614 nsew ground input
rlabel locali s 298695 248333 298799 248441 6 VGND
port 614 nsew ground input
rlabel locali s 1121 248333 1225 248441 6 VGND
port 614 nsew ground input
rlabel locali s 298660 248441 298799 248591 6 VGND
port 614 nsew ground input
rlabel locali s 298660 248591 298816 248625 6 VGND
port 614 nsew ground input
rlabel locali s 298660 248625 298799 248775 6 VGND
port 614 nsew ground input
rlabel locali s 1121 248441 1340 248591 6 VGND
port 614 nsew ground input
rlabel locali s 1104 248591 1340 248625 6 VGND
port 614 nsew ground input
rlabel locali s 1121 248625 1340 248775 6 VGND
port 614 nsew ground input
rlabel locali s 298695 248775 298799 248883 6 VGND
port 614 nsew ground input
rlabel locali s 1121 248775 1225 248883 6 VGND
port 614 nsew ground input
rlabel locali s 298695 249421 298799 249529 6 VGND
port 614 nsew ground input
rlabel locali s 1121 249421 1225 249529 6 VGND
port 614 nsew ground input
rlabel locali s 298660 249529 298799 249679 6 VGND
port 614 nsew ground input
rlabel locali s 298660 249679 298816 249713 6 VGND
port 614 nsew ground input
rlabel locali s 298660 249713 298799 249863 6 VGND
port 614 nsew ground input
rlabel locali s 1121 249529 1340 249679 6 VGND
port 614 nsew ground input
rlabel locali s 1104 249679 1340 249713 6 VGND
port 614 nsew ground input
rlabel locali s 1121 249713 1340 249863 6 VGND
port 614 nsew ground input
rlabel locali s 298695 249863 298799 249971 6 VGND
port 614 nsew ground input
rlabel locali s 1121 249863 1225 249971 6 VGND
port 614 nsew ground input
rlabel locali s 298695 250509 298799 250617 6 VGND
port 614 nsew ground input
rlabel locali s 1121 250509 1225 250617 6 VGND
port 614 nsew ground input
rlabel locali s 298660 250617 298799 250767 6 VGND
port 614 nsew ground input
rlabel locali s 298660 250767 298816 250801 6 VGND
port 614 nsew ground input
rlabel locali s 298660 250801 298799 250951 6 VGND
port 614 nsew ground input
rlabel locali s 1121 250617 1340 250767 6 VGND
port 614 nsew ground input
rlabel locali s 1104 250767 1340 250801 6 VGND
port 614 nsew ground input
rlabel locali s 1121 250801 1340 250951 6 VGND
port 614 nsew ground input
rlabel locali s 298695 250951 298799 251059 6 VGND
port 614 nsew ground input
rlabel locali s 1121 250951 1225 251059 6 VGND
port 614 nsew ground input
rlabel locali s 298695 251597 298799 251705 6 VGND
port 614 nsew ground input
rlabel locali s 1121 251597 1225 251705 6 VGND
port 614 nsew ground input
rlabel locali s 298660 251705 298799 251855 6 VGND
port 614 nsew ground input
rlabel locali s 298660 251855 298816 251889 6 VGND
port 614 nsew ground input
rlabel locali s 298660 251889 298799 252039 6 VGND
port 614 nsew ground input
rlabel locali s 1121 251705 1340 251855 6 VGND
port 614 nsew ground input
rlabel locali s 1104 251855 1340 251889 6 VGND
port 614 nsew ground input
rlabel locali s 1121 251889 1340 252039 6 VGND
port 614 nsew ground input
rlabel locali s 298695 252039 298799 252147 6 VGND
port 614 nsew ground input
rlabel locali s 1121 252039 1225 252147 6 VGND
port 614 nsew ground input
rlabel locali s 298695 252685 298799 252793 6 VGND
port 614 nsew ground input
rlabel locali s 1121 252685 1225 252793 6 VGND
port 614 nsew ground input
rlabel locali s 298660 252793 298799 252943 6 VGND
port 614 nsew ground input
rlabel locali s 298660 252943 298816 252977 6 VGND
port 614 nsew ground input
rlabel locali s 298660 252977 298799 253127 6 VGND
port 614 nsew ground input
rlabel locali s 1121 252793 1340 252943 6 VGND
port 614 nsew ground input
rlabel locali s 1104 252943 1340 252977 6 VGND
port 614 nsew ground input
rlabel locali s 1121 252977 1340 253127 6 VGND
port 614 nsew ground input
rlabel locali s 298695 253127 298799 253235 6 VGND
port 614 nsew ground input
rlabel locali s 1121 253127 1225 253235 6 VGND
port 614 nsew ground input
rlabel locali s 298695 253773 298799 253881 6 VGND
port 614 nsew ground input
rlabel locali s 1121 253773 1225 253881 6 VGND
port 614 nsew ground input
rlabel locali s 298660 253881 298799 254031 6 VGND
port 614 nsew ground input
rlabel locali s 298660 254031 298816 254065 6 VGND
port 614 nsew ground input
rlabel locali s 298660 254065 298799 254215 6 VGND
port 614 nsew ground input
rlabel locali s 1121 253881 1340 254031 6 VGND
port 614 nsew ground input
rlabel locali s 1104 254031 1340 254065 6 VGND
port 614 nsew ground input
rlabel locali s 1121 254065 1340 254215 6 VGND
port 614 nsew ground input
rlabel locali s 298695 254215 298799 254323 6 VGND
port 614 nsew ground input
rlabel locali s 1121 254215 1225 254323 6 VGND
port 614 nsew ground input
rlabel locali s 298695 254861 298799 254969 6 VGND
port 614 nsew ground input
rlabel locali s 1121 254861 1225 254969 6 VGND
port 614 nsew ground input
rlabel locali s 298660 254969 298799 255119 6 VGND
port 614 nsew ground input
rlabel locali s 298660 255119 298816 255153 6 VGND
port 614 nsew ground input
rlabel locali s 298660 255153 298799 255303 6 VGND
port 614 nsew ground input
rlabel locali s 1121 254969 1340 255119 6 VGND
port 614 nsew ground input
rlabel locali s 1104 255119 1340 255153 6 VGND
port 614 nsew ground input
rlabel locali s 1121 255153 1340 255303 6 VGND
port 614 nsew ground input
rlabel locali s 298695 255303 298799 255411 6 VGND
port 614 nsew ground input
rlabel locali s 1121 255303 1225 255411 6 VGND
port 614 nsew ground input
rlabel locali s 298695 255949 298799 256057 6 VGND
port 614 nsew ground input
rlabel locali s 1121 255949 1225 256057 6 VGND
port 614 nsew ground input
rlabel locali s 298660 256057 298799 256207 6 VGND
port 614 nsew ground input
rlabel locali s 298660 256207 298816 256241 6 VGND
port 614 nsew ground input
rlabel locali s 298660 256241 298799 256391 6 VGND
port 614 nsew ground input
rlabel locali s 1121 256057 1340 256207 6 VGND
port 614 nsew ground input
rlabel locali s 1104 256207 1340 256241 6 VGND
port 614 nsew ground input
rlabel locali s 1121 256241 1340 256391 6 VGND
port 614 nsew ground input
rlabel locali s 298695 256391 298799 256499 6 VGND
port 614 nsew ground input
rlabel locali s 1121 256391 1225 256499 6 VGND
port 614 nsew ground input
rlabel locali s 298695 257037 298799 257145 6 VGND
port 614 nsew ground input
rlabel locali s 1121 257037 1225 257145 6 VGND
port 614 nsew ground input
rlabel locali s 298660 257145 298799 257295 6 VGND
port 614 nsew ground input
rlabel locali s 298660 257295 298816 257329 6 VGND
port 614 nsew ground input
rlabel locali s 298660 257329 298799 257479 6 VGND
port 614 nsew ground input
rlabel locali s 1121 257145 1340 257295 6 VGND
port 614 nsew ground input
rlabel locali s 1104 257295 1340 257329 6 VGND
port 614 nsew ground input
rlabel locali s 1121 257329 1340 257479 6 VGND
port 614 nsew ground input
rlabel locali s 298695 257479 298799 257587 6 VGND
port 614 nsew ground input
rlabel locali s 1121 257479 1225 257587 6 VGND
port 614 nsew ground input
rlabel locali s 298695 258125 298799 258233 6 VGND
port 614 nsew ground input
rlabel locali s 1121 258125 1225 258233 6 VGND
port 614 nsew ground input
rlabel locali s 298660 258233 298799 258383 6 VGND
port 614 nsew ground input
rlabel locali s 298660 258383 298816 258417 6 VGND
port 614 nsew ground input
rlabel locali s 298660 258417 298799 258567 6 VGND
port 614 nsew ground input
rlabel locali s 1121 258233 1340 258383 6 VGND
port 614 nsew ground input
rlabel locali s 1104 258383 1340 258417 6 VGND
port 614 nsew ground input
rlabel locali s 1121 258417 1340 258567 6 VGND
port 614 nsew ground input
rlabel locali s 298695 258567 298799 258675 6 VGND
port 614 nsew ground input
rlabel locali s 1121 258567 1225 258675 6 VGND
port 614 nsew ground input
rlabel locali s 298695 259213 298799 259321 6 VGND
port 614 nsew ground input
rlabel locali s 1121 259213 1225 259321 6 VGND
port 614 nsew ground input
rlabel locali s 298660 259321 298799 259471 6 VGND
port 614 nsew ground input
rlabel locali s 298660 259471 298816 259505 6 VGND
port 614 nsew ground input
rlabel locali s 298660 259505 298799 259655 6 VGND
port 614 nsew ground input
rlabel locali s 1121 259321 1340 259471 6 VGND
port 614 nsew ground input
rlabel locali s 1104 259471 1340 259505 6 VGND
port 614 nsew ground input
rlabel locali s 1121 259505 1340 259655 6 VGND
port 614 nsew ground input
rlabel locali s 298695 259655 298799 259763 6 VGND
port 614 nsew ground input
rlabel locali s 1121 259655 1225 259763 6 VGND
port 614 nsew ground input
rlabel locali s 298695 260301 298799 260409 6 VGND
port 614 nsew ground input
rlabel locali s 1121 260301 1225 260409 6 VGND
port 614 nsew ground input
rlabel locali s 298660 260409 298799 260559 6 VGND
port 614 nsew ground input
rlabel locali s 298660 260559 298816 260593 6 VGND
port 614 nsew ground input
rlabel locali s 298660 260593 298799 260743 6 VGND
port 614 nsew ground input
rlabel locali s 1121 260409 1340 260559 6 VGND
port 614 nsew ground input
rlabel locali s 1104 260559 1340 260593 6 VGND
port 614 nsew ground input
rlabel locali s 1121 260593 1340 260743 6 VGND
port 614 nsew ground input
rlabel locali s 298695 260743 298799 260851 6 VGND
port 614 nsew ground input
rlabel locali s 1121 260743 1225 260851 6 VGND
port 614 nsew ground input
rlabel locali s 298695 261389 298799 261497 6 VGND
port 614 nsew ground input
rlabel locali s 1121 261389 1225 261497 6 VGND
port 614 nsew ground input
rlabel locali s 298660 261497 298799 261647 6 VGND
port 614 nsew ground input
rlabel locali s 298660 261647 298816 261681 6 VGND
port 614 nsew ground input
rlabel locali s 298660 261681 298799 261831 6 VGND
port 614 nsew ground input
rlabel locali s 1121 261497 1340 261647 6 VGND
port 614 nsew ground input
rlabel locali s 1104 261647 1340 261681 6 VGND
port 614 nsew ground input
rlabel locali s 1121 261681 1340 261831 6 VGND
port 614 nsew ground input
rlabel locali s 298695 261831 298799 261939 6 VGND
port 614 nsew ground input
rlabel locali s 1121 261831 1225 261939 6 VGND
port 614 nsew ground input
rlabel locali s 298695 262477 298799 262585 6 VGND
port 614 nsew ground input
rlabel locali s 1121 262477 1225 262585 6 VGND
port 614 nsew ground input
rlabel locali s 298660 262585 298799 262735 6 VGND
port 614 nsew ground input
rlabel locali s 298660 262735 298816 262769 6 VGND
port 614 nsew ground input
rlabel locali s 298660 262769 298799 262919 6 VGND
port 614 nsew ground input
rlabel locali s 1121 262585 1340 262735 6 VGND
port 614 nsew ground input
rlabel locali s 1104 262735 1340 262769 6 VGND
port 614 nsew ground input
rlabel locali s 1121 262769 1340 262919 6 VGND
port 614 nsew ground input
rlabel locali s 298695 262919 298799 263027 6 VGND
port 614 nsew ground input
rlabel locali s 1121 262919 1225 263027 6 VGND
port 614 nsew ground input
rlabel locali s 298695 263565 298799 263673 6 VGND
port 614 nsew ground input
rlabel locali s 1121 263565 1225 263673 6 VGND
port 614 nsew ground input
rlabel locali s 298660 263673 298799 263823 6 VGND
port 614 nsew ground input
rlabel locali s 298660 263823 298816 263857 6 VGND
port 614 nsew ground input
rlabel locali s 298660 263857 298799 264007 6 VGND
port 614 nsew ground input
rlabel locali s 1121 263673 1340 263823 6 VGND
port 614 nsew ground input
rlabel locali s 1104 263823 1340 263857 6 VGND
port 614 nsew ground input
rlabel locali s 1121 263857 1340 264007 6 VGND
port 614 nsew ground input
rlabel locali s 298695 264007 298799 264115 6 VGND
port 614 nsew ground input
rlabel locali s 1121 264007 1225 264115 6 VGND
port 614 nsew ground input
rlabel locali s 298695 264653 298799 264761 6 VGND
port 614 nsew ground input
rlabel locali s 1121 264653 1225 264761 6 VGND
port 614 nsew ground input
rlabel locali s 298660 264761 298799 264911 6 VGND
port 614 nsew ground input
rlabel locali s 298660 264911 298816 264945 6 VGND
port 614 nsew ground input
rlabel locali s 298660 264945 298799 265095 6 VGND
port 614 nsew ground input
rlabel locali s 1121 264761 1340 264911 6 VGND
port 614 nsew ground input
rlabel locali s 1104 264911 1340 264945 6 VGND
port 614 nsew ground input
rlabel locali s 1121 264945 1340 265095 6 VGND
port 614 nsew ground input
rlabel locali s 298695 265095 298799 265203 6 VGND
port 614 nsew ground input
rlabel locali s 1121 265095 1225 265203 6 VGND
port 614 nsew ground input
rlabel locali s 298695 265741 298799 265849 6 VGND
port 614 nsew ground input
rlabel locali s 1121 265741 1225 265849 6 VGND
port 614 nsew ground input
rlabel locali s 298660 265849 298799 265999 6 VGND
port 614 nsew ground input
rlabel locali s 298660 265999 298816 266033 6 VGND
port 614 nsew ground input
rlabel locali s 298660 266033 298799 266183 6 VGND
port 614 nsew ground input
rlabel locali s 1121 265849 1340 265999 6 VGND
port 614 nsew ground input
rlabel locali s 1104 265999 1340 266033 6 VGND
port 614 nsew ground input
rlabel locali s 1121 266033 1340 266183 6 VGND
port 614 nsew ground input
rlabel locali s 298695 266183 298799 266291 6 VGND
port 614 nsew ground input
rlabel locali s 1121 266183 1225 266291 6 VGND
port 614 nsew ground input
rlabel locali s 298695 266829 298799 266937 6 VGND
port 614 nsew ground input
rlabel locali s 1121 266829 1225 266937 6 VGND
port 614 nsew ground input
rlabel locali s 298660 266937 298799 267087 6 VGND
port 614 nsew ground input
rlabel locali s 298660 267087 298816 267121 6 VGND
port 614 nsew ground input
rlabel locali s 298660 267121 298799 267271 6 VGND
port 614 nsew ground input
rlabel locali s 1121 266937 1340 267087 6 VGND
port 614 nsew ground input
rlabel locali s 1104 267087 1340 267121 6 VGND
port 614 nsew ground input
rlabel locali s 1121 267121 1340 267271 6 VGND
port 614 nsew ground input
rlabel locali s 298695 267271 298799 267379 6 VGND
port 614 nsew ground input
rlabel locali s 1121 267271 1225 267379 6 VGND
port 614 nsew ground input
rlabel locali s 298695 267917 298799 268025 6 VGND
port 614 nsew ground input
rlabel locali s 1121 267917 1225 268025 6 VGND
port 614 nsew ground input
rlabel locali s 298660 268025 298799 268175 6 VGND
port 614 nsew ground input
rlabel locali s 298660 268175 298816 268209 6 VGND
port 614 nsew ground input
rlabel locali s 298660 268209 298799 268359 6 VGND
port 614 nsew ground input
rlabel locali s 1121 268025 1340 268175 6 VGND
port 614 nsew ground input
rlabel locali s 1104 268175 1340 268209 6 VGND
port 614 nsew ground input
rlabel locali s 1121 268209 1340 268359 6 VGND
port 614 nsew ground input
rlabel locali s 298695 268359 298799 268467 6 VGND
port 614 nsew ground input
rlabel locali s 1121 268359 1225 268467 6 VGND
port 614 nsew ground input
rlabel locali s 298695 269005 298799 269113 6 VGND
port 614 nsew ground input
rlabel locali s 1121 269005 1225 269113 6 VGND
port 614 nsew ground input
rlabel locali s 298660 269113 298799 269263 6 VGND
port 614 nsew ground input
rlabel locali s 298660 269263 298816 269297 6 VGND
port 614 nsew ground input
rlabel locali s 298660 269297 298799 269447 6 VGND
port 614 nsew ground input
rlabel locali s 1121 269113 1340 269263 6 VGND
port 614 nsew ground input
rlabel locali s 1104 269263 1340 269297 6 VGND
port 614 nsew ground input
rlabel locali s 1121 269297 1340 269447 6 VGND
port 614 nsew ground input
rlabel locali s 298695 269447 298799 269555 6 VGND
port 614 nsew ground input
rlabel locali s 1121 269447 1225 269555 6 VGND
port 614 nsew ground input
rlabel locali s 298695 270093 298799 270201 6 VGND
port 614 nsew ground input
rlabel locali s 1121 270093 1225 270201 6 VGND
port 614 nsew ground input
rlabel locali s 298660 270201 298799 270351 6 VGND
port 614 nsew ground input
rlabel locali s 298660 270351 298816 270385 6 VGND
port 614 nsew ground input
rlabel locali s 298660 270385 298799 270535 6 VGND
port 614 nsew ground input
rlabel locali s 1121 270201 1340 270351 6 VGND
port 614 nsew ground input
rlabel locali s 1104 270351 1340 270385 6 VGND
port 614 nsew ground input
rlabel locali s 1121 270385 1340 270535 6 VGND
port 614 nsew ground input
rlabel locali s 298695 270535 298799 270643 6 VGND
port 614 nsew ground input
rlabel locali s 1121 270535 1225 270643 6 VGND
port 614 nsew ground input
rlabel locali s 298695 271181 298799 271289 6 VGND
port 614 nsew ground input
rlabel locali s 1121 271181 1225 271289 6 VGND
port 614 nsew ground input
rlabel locali s 298660 271289 298799 271439 6 VGND
port 614 nsew ground input
rlabel locali s 298660 271439 298816 271473 6 VGND
port 614 nsew ground input
rlabel locali s 298660 271473 298799 271623 6 VGND
port 614 nsew ground input
rlabel locali s 1121 271289 1340 271439 6 VGND
port 614 nsew ground input
rlabel locali s 1104 271439 1340 271473 6 VGND
port 614 nsew ground input
rlabel locali s 1121 271473 1340 271623 6 VGND
port 614 nsew ground input
rlabel locali s 298695 271623 298799 271731 6 VGND
port 614 nsew ground input
rlabel locali s 1121 271623 1225 271731 6 VGND
port 614 nsew ground input
rlabel locali s 298695 272269 298799 272377 6 VGND
port 614 nsew ground input
rlabel locali s 1121 272269 1225 272377 6 VGND
port 614 nsew ground input
rlabel locali s 298660 272377 298799 272527 6 VGND
port 614 nsew ground input
rlabel locali s 298660 272527 298816 272561 6 VGND
port 614 nsew ground input
rlabel locali s 298660 272561 298799 272711 6 VGND
port 614 nsew ground input
rlabel locali s 1121 272377 1340 272527 6 VGND
port 614 nsew ground input
rlabel locali s 1104 272527 1340 272561 6 VGND
port 614 nsew ground input
rlabel locali s 1121 272561 1340 272711 6 VGND
port 614 nsew ground input
rlabel locali s 298695 272711 298799 272819 6 VGND
port 614 nsew ground input
rlabel locali s 1121 272711 1225 272819 6 VGND
port 614 nsew ground input
rlabel locali s 298695 273357 298799 273465 6 VGND
port 614 nsew ground input
rlabel locali s 1121 273357 1225 273465 6 VGND
port 614 nsew ground input
rlabel locali s 298660 273465 298799 273615 6 VGND
port 614 nsew ground input
rlabel locali s 298660 273615 298816 273649 6 VGND
port 614 nsew ground input
rlabel locali s 298660 273649 298799 273799 6 VGND
port 614 nsew ground input
rlabel locali s 1121 273465 1340 273615 6 VGND
port 614 nsew ground input
rlabel locali s 1104 273615 1340 273649 6 VGND
port 614 nsew ground input
rlabel locali s 1121 273649 1340 273799 6 VGND
port 614 nsew ground input
rlabel locali s 298695 273799 298799 273907 6 VGND
port 614 nsew ground input
rlabel locali s 1121 273799 1225 273907 6 VGND
port 614 nsew ground input
rlabel locali s 298695 274445 298799 274553 6 VGND
port 614 nsew ground input
rlabel locali s 1121 274445 1225 274553 6 VGND
port 614 nsew ground input
rlabel locali s 298660 274553 298799 274703 6 VGND
port 614 nsew ground input
rlabel locali s 298660 274703 298816 274737 6 VGND
port 614 nsew ground input
rlabel locali s 298660 274737 298799 274887 6 VGND
port 614 nsew ground input
rlabel locali s 1121 274553 1340 274703 6 VGND
port 614 nsew ground input
rlabel locali s 1104 274703 1340 274737 6 VGND
port 614 nsew ground input
rlabel locali s 1121 274737 1340 274887 6 VGND
port 614 nsew ground input
rlabel locali s 298695 274887 298799 274995 6 VGND
port 614 nsew ground input
rlabel locali s 1121 274887 1225 274995 6 VGND
port 614 nsew ground input
rlabel locali s 298695 275533 298799 275641 6 VGND
port 614 nsew ground input
rlabel locali s 1121 275533 1225 275641 6 VGND
port 614 nsew ground input
rlabel locali s 298660 275641 298799 275791 6 VGND
port 614 nsew ground input
rlabel locali s 298660 275791 298816 275825 6 VGND
port 614 nsew ground input
rlabel locali s 298660 275825 298799 275975 6 VGND
port 614 nsew ground input
rlabel locali s 1121 275641 1340 275791 6 VGND
port 614 nsew ground input
rlabel locali s 1104 275791 1340 275825 6 VGND
port 614 nsew ground input
rlabel locali s 1121 275825 1340 275975 6 VGND
port 614 nsew ground input
rlabel locali s 298695 275975 298799 276083 6 VGND
port 614 nsew ground input
rlabel locali s 1121 275975 1225 276083 6 VGND
port 614 nsew ground input
rlabel locali s 298695 276621 298799 276729 6 VGND
port 614 nsew ground input
rlabel locali s 1121 276621 1225 276729 6 VGND
port 614 nsew ground input
rlabel locali s 298660 276729 298799 276879 6 VGND
port 614 nsew ground input
rlabel locali s 298660 276879 298816 276913 6 VGND
port 614 nsew ground input
rlabel locali s 298660 276913 298799 277063 6 VGND
port 614 nsew ground input
rlabel locali s 1121 276729 1340 276879 6 VGND
port 614 nsew ground input
rlabel locali s 1104 276879 1340 276913 6 VGND
port 614 nsew ground input
rlabel locali s 1121 276913 1340 277063 6 VGND
port 614 nsew ground input
rlabel locali s 298695 277063 298799 277171 6 VGND
port 614 nsew ground input
rlabel locali s 1121 277063 1225 277171 6 VGND
port 614 nsew ground input
rlabel locali s 298695 277709 298799 277817 6 VGND
port 614 nsew ground input
rlabel locali s 1121 277709 1225 277817 6 VGND
port 614 nsew ground input
rlabel locali s 298660 277817 298799 277967 6 VGND
port 614 nsew ground input
rlabel locali s 298660 277967 298816 278001 6 VGND
port 614 nsew ground input
rlabel locali s 298660 278001 298799 278151 6 VGND
port 614 nsew ground input
rlabel locali s 1121 277817 1340 277967 6 VGND
port 614 nsew ground input
rlabel locali s 1104 277967 1340 278001 6 VGND
port 614 nsew ground input
rlabel locali s 1121 278001 1340 278151 6 VGND
port 614 nsew ground input
rlabel locali s 298695 278151 298799 278259 6 VGND
port 614 nsew ground input
rlabel locali s 1121 278151 1225 278259 6 VGND
port 614 nsew ground input
rlabel locali s 298695 278797 298799 278905 6 VGND
port 614 nsew ground input
rlabel locali s 1121 278797 1225 278905 6 VGND
port 614 nsew ground input
rlabel locali s 298660 278905 298799 279055 6 VGND
port 614 nsew ground input
rlabel locali s 298660 279055 298816 279089 6 VGND
port 614 nsew ground input
rlabel locali s 298660 279089 298799 279239 6 VGND
port 614 nsew ground input
rlabel locali s 1121 278905 1340 279055 6 VGND
port 614 nsew ground input
rlabel locali s 1104 279055 1340 279089 6 VGND
port 614 nsew ground input
rlabel locali s 1121 279089 1340 279239 6 VGND
port 614 nsew ground input
rlabel locali s 298695 279239 298799 279347 6 VGND
port 614 nsew ground input
rlabel locali s 1121 279239 1225 279347 6 VGND
port 614 nsew ground input
rlabel locali s 298695 279885 298799 279993 6 VGND
port 614 nsew ground input
rlabel locali s 1121 279885 1225 279993 6 VGND
port 614 nsew ground input
rlabel locali s 298660 279993 298799 280143 6 VGND
port 614 nsew ground input
rlabel locali s 298660 280143 298816 280177 6 VGND
port 614 nsew ground input
rlabel locali s 298660 280177 298799 280327 6 VGND
port 614 nsew ground input
rlabel locali s 1121 279993 1340 280143 6 VGND
port 614 nsew ground input
rlabel locali s 1104 280143 1340 280177 6 VGND
port 614 nsew ground input
rlabel locali s 1121 280177 1340 280327 6 VGND
port 614 nsew ground input
rlabel locali s 298695 280327 298799 280435 6 VGND
port 614 nsew ground input
rlabel locali s 1121 280327 1225 280435 6 VGND
port 614 nsew ground input
rlabel locali s 298695 280973 298799 281081 6 VGND
port 614 nsew ground input
rlabel locali s 1121 280973 1225 281081 6 VGND
port 614 nsew ground input
rlabel locali s 298660 281081 298799 281231 6 VGND
port 614 nsew ground input
rlabel locali s 298660 281231 298816 281265 6 VGND
port 614 nsew ground input
rlabel locali s 298660 281265 298799 281415 6 VGND
port 614 nsew ground input
rlabel locali s 1121 281081 1340 281231 6 VGND
port 614 nsew ground input
rlabel locali s 1104 281231 1340 281265 6 VGND
port 614 nsew ground input
rlabel locali s 1121 281265 1340 281415 6 VGND
port 614 nsew ground input
rlabel locali s 298695 281415 298799 281523 6 VGND
port 614 nsew ground input
rlabel locali s 1121 281415 1225 281523 6 VGND
port 614 nsew ground input
rlabel locali s 298695 282061 298799 282169 6 VGND
port 614 nsew ground input
rlabel locali s 1121 282061 1225 282169 6 VGND
port 614 nsew ground input
rlabel locali s 298660 282169 298799 282319 6 VGND
port 614 nsew ground input
rlabel locali s 298660 282319 298816 282353 6 VGND
port 614 nsew ground input
rlabel locali s 298660 282353 298799 282503 6 VGND
port 614 nsew ground input
rlabel locali s 1121 282169 1340 282319 6 VGND
port 614 nsew ground input
rlabel locali s 1104 282319 1340 282353 6 VGND
port 614 nsew ground input
rlabel locali s 1121 282353 1340 282503 6 VGND
port 614 nsew ground input
rlabel locali s 298695 282503 298799 282611 6 VGND
port 614 nsew ground input
rlabel locali s 1121 282503 1225 282611 6 VGND
port 614 nsew ground input
rlabel locali s 298695 283149 298799 283257 6 VGND
port 614 nsew ground input
rlabel locali s 1121 283149 1225 283257 6 VGND
port 614 nsew ground input
rlabel locali s 298660 283257 298799 283407 6 VGND
port 614 nsew ground input
rlabel locali s 298660 283407 298816 283441 6 VGND
port 614 nsew ground input
rlabel locali s 298660 283441 298799 283591 6 VGND
port 614 nsew ground input
rlabel locali s 1121 283257 1340 283407 6 VGND
port 614 nsew ground input
rlabel locali s 1104 283407 1340 283441 6 VGND
port 614 nsew ground input
rlabel locali s 1121 283441 1340 283591 6 VGND
port 614 nsew ground input
rlabel locali s 298695 283591 298799 283699 6 VGND
port 614 nsew ground input
rlabel locali s 1121 283591 1225 283699 6 VGND
port 614 nsew ground input
rlabel locali s 298695 284237 298799 284345 6 VGND
port 614 nsew ground input
rlabel locali s 1121 284237 1225 284345 6 VGND
port 614 nsew ground input
rlabel locali s 298660 284345 298799 284495 6 VGND
port 614 nsew ground input
rlabel locali s 298660 284495 298816 284529 6 VGND
port 614 nsew ground input
rlabel locali s 298660 284529 298799 284679 6 VGND
port 614 nsew ground input
rlabel locali s 1121 284345 1340 284495 6 VGND
port 614 nsew ground input
rlabel locali s 1104 284495 1340 284529 6 VGND
port 614 nsew ground input
rlabel locali s 1121 284529 1340 284679 6 VGND
port 614 nsew ground input
rlabel locali s 298695 284679 298799 284787 6 VGND
port 614 nsew ground input
rlabel locali s 1121 284679 1225 284787 6 VGND
port 614 nsew ground input
rlabel locali s 298695 285325 298799 285433 6 VGND
port 614 nsew ground input
rlabel locali s 1121 285325 1225 285433 6 VGND
port 614 nsew ground input
rlabel locali s 298660 285433 298799 285583 6 VGND
port 614 nsew ground input
rlabel locali s 298660 285583 298816 285617 6 VGND
port 614 nsew ground input
rlabel locali s 298660 285617 298799 285767 6 VGND
port 614 nsew ground input
rlabel locali s 1121 285433 1340 285583 6 VGND
port 614 nsew ground input
rlabel locali s 1104 285583 1340 285617 6 VGND
port 614 nsew ground input
rlabel locali s 1121 285617 1340 285767 6 VGND
port 614 nsew ground input
rlabel locali s 298695 285767 298799 285875 6 VGND
port 614 nsew ground input
rlabel locali s 1121 285767 1225 285875 6 VGND
port 614 nsew ground input
rlabel locali s 298695 286413 298799 286521 6 VGND
port 614 nsew ground input
rlabel locali s 1121 286413 1225 286521 6 VGND
port 614 nsew ground input
rlabel locali s 298660 286521 298799 286671 6 VGND
port 614 nsew ground input
rlabel locali s 298660 286671 298816 286705 6 VGND
port 614 nsew ground input
rlabel locali s 298660 286705 298799 286855 6 VGND
port 614 nsew ground input
rlabel locali s 1121 286521 1340 286671 6 VGND
port 614 nsew ground input
rlabel locali s 1104 286671 1340 286705 6 VGND
port 614 nsew ground input
rlabel locali s 1121 286705 1340 286855 6 VGND
port 614 nsew ground input
rlabel locali s 298695 286855 298799 286963 6 VGND
port 614 nsew ground input
rlabel locali s 1121 286855 1225 286963 6 VGND
port 614 nsew ground input
rlabel locali s 298695 287501 298799 287609 6 VGND
port 614 nsew ground input
rlabel locali s 1121 287501 1225 287609 6 VGND
port 614 nsew ground input
rlabel locali s 298660 287609 298799 287759 6 VGND
port 614 nsew ground input
rlabel locali s 298660 287759 298816 287793 6 VGND
port 614 nsew ground input
rlabel locali s 298660 287793 298799 287943 6 VGND
port 614 nsew ground input
rlabel locali s 1121 287609 1340 287759 6 VGND
port 614 nsew ground input
rlabel locali s 1104 287759 1340 287793 6 VGND
port 614 nsew ground input
rlabel locali s 1121 287793 1340 287943 6 VGND
port 614 nsew ground input
rlabel locali s 298695 287943 298799 288051 6 VGND
port 614 nsew ground input
rlabel locali s 1121 287943 1225 288051 6 VGND
port 614 nsew ground input
rlabel locali s 298695 288589 298799 288697 6 VGND
port 614 nsew ground input
rlabel locali s 1121 288589 1225 288697 6 VGND
port 614 nsew ground input
rlabel locali s 298660 288697 298799 288847 6 VGND
port 614 nsew ground input
rlabel locali s 298660 288847 298816 288881 6 VGND
port 614 nsew ground input
rlabel locali s 298660 288881 298799 289031 6 VGND
port 614 nsew ground input
rlabel locali s 1121 288697 1340 288847 6 VGND
port 614 nsew ground input
rlabel locali s 1104 288847 1340 288881 6 VGND
port 614 nsew ground input
rlabel locali s 1121 288881 1340 289031 6 VGND
port 614 nsew ground input
rlabel locali s 298695 289031 298799 289139 6 VGND
port 614 nsew ground input
rlabel locali s 1121 289031 1225 289139 6 VGND
port 614 nsew ground input
rlabel locali s 298695 289677 298799 289785 6 VGND
port 614 nsew ground input
rlabel locali s 1121 289677 1225 289785 6 VGND
port 614 nsew ground input
rlabel locali s 298660 289785 298799 289935 6 VGND
port 614 nsew ground input
rlabel locali s 298660 289935 298816 289969 6 VGND
port 614 nsew ground input
rlabel locali s 298660 289969 298799 290119 6 VGND
port 614 nsew ground input
rlabel locali s 1121 289785 1340 289935 6 VGND
port 614 nsew ground input
rlabel locali s 1104 289935 1340 289969 6 VGND
port 614 nsew ground input
rlabel locali s 1121 289969 1340 290119 6 VGND
port 614 nsew ground input
rlabel locali s 298695 290119 298799 290227 6 VGND
port 614 nsew ground input
rlabel locali s 1121 290119 1225 290227 6 VGND
port 614 nsew ground input
rlabel locali s 298695 290765 298799 290873 6 VGND
port 614 nsew ground input
rlabel locali s 1121 290765 1225 290873 6 VGND
port 614 nsew ground input
rlabel locali s 298660 290873 298799 291023 6 VGND
port 614 nsew ground input
rlabel locali s 298660 291023 298816 291057 6 VGND
port 614 nsew ground input
rlabel locali s 298660 291057 298799 291207 6 VGND
port 614 nsew ground input
rlabel locali s 1121 290873 1340 291023 6 VGND
port 614 nsew ground input
rlabel locali s 1104 291023 1340 291057 6 VGND
port 614 nsew ground input
rlabel locali s 1121 291057 1340 291207 6 VGND
port 614 nsew ground input
rlabel locali s 298695 291207 298799 291315 6 VGND
port 614 nsew ground input
rlabel locali s 1121 291207 1225 291315 6 VGND
port 614 nsew ground input
rlabel locali s 298695 291853 298799 291961 6 VGND
port 614 nsew ground input
rlabel locali s 1121 291853 1225 291961 6 VGND
port 614 nsew ground input
rlabel locali s 298660 291961 298799 292111 6 VGND
port 614 nsew ground input
rlabel locali s 298660 292111 298816 292145 6 VGND
port 614 nsew ground input
rlabel locali s 298660 292145 298799 292295 6 VGND
port 614 nsew ground input
rlabel locali s 1121 291961 1340 292111 6 VGND
port 614 nsew ground input
rlabel locali s 1104 292111 1340 292145 6 VGND
port 614 nsew ground input
rlabel locali s 1121 292145 1340 292295 6 VGND
port 614 nsew ground input
rlabel locali s 298695 292295 298799 292403 6 VGND
port 614 nsew ground input
rlabel locali s 1121 292295 1225 292403 6 VGND
port 614 nsew ground input
rlabel locali s 298695 292941 298799 293049 6 VGND
port 614 nsew ground input
rlabel locali s 1121 292941 1225 293049 6 VGND
port 614 nsew ground input
rlabel locali s 298660 293049 298799 293199 6 VGND
port 614 nsew ground input
rlabel locali s 298660 293199 298816 293233 6 VGND
port 614 nsew ground input
rlabel locali s 298660 293233 298799 293383 6 VGND
port 614 nsew ground input
rlabel locali s 1121 293049 1340 293199 6 VGND
port 614 nsew ground input
rlabel locali s 1104 293199 1340 293233 6 VGND
port 614 nsew ground input
rlabel locali s 1121 293233 1340 293383 6 VGND
port 614 nsew ground input
rlabel locali s 298695 293383 298799 293491 6 VGND
port 614 nsew ground input
rlabel locali s 1121 293383 1225 293491 6 VGND
port 614 nsew ground input
rlabel locali s 298695 294029 298799 294137 6 VGND
port 614 nsew ground input
rlabel locali s 1121 294029 1225 294137 6 VGND
port 614 nsew ground input
rlabel locali s 298660 294137 298799 294287 6 VGND
port 614 nsew ground input
rlabel locali s 298660 294287 298816 294321 6 VGND
port 614 nsew ground input
rlabel locali s 298660 294321 298799 294471 6 VGND
port 614 nsew ground input
rlabel locali s 1121 294137 1340 294287 6 VGND
port 614 nsew ground input
rlabel locali s 1104 294287 1340 294321 6 VGND
port 614 nsew ground input
rlabel locali s 1121 294321 1340 294471 6 VGND
port 614 nsew ground input
rlabel locali s 298695 294471 298799 294579 6 VGND
port 614 nsew ground input
rlabel locali s 1121 294471 1225 294579 6 VGND
port 614 nsew ground input
rlabel locali s 298695 295117 298799 295225 6 VGND
port 614 nsew ground input
rlabel locali s 1121 295117 1225 295225 6 VGND
port 614 nsew ground input
rlabel locali s 298660 295225 298799 295375 6 VGND
port 614 nsew ground input
rlabel locali s 298660 295375 298816 295409 6 VGND
port 614 nsew ground input
rlabel locali s 298660 295409 298799 295559 6 VGND
port 614 nsew ground input
rlabel locali s 1121 295225 1340 295375 6 VGND
port 614 nsew ground input
rlabel locali s 1104 295375 1340 295409 6 VGND
port 614 nsew ground input
rlabel locali s 1121 295409 1340 295559 6 VGND
port 614 nsew ground input
rlabel locali s 298695 295559 298799 295667 6 VGND
port 614 nsew ground input
rlabel locali s 1121 295559 1225 295667 6 VGND
port 614 nsew ground input
rlabel locali s 298695 296205 298799 296313 6 VGND
port 614 nsew ground input
rlabel locali s 1121 296205 1225 296313 6 VGND
port 614 nsew ground input
rlabel locali s 298660 296313 298799 296463 6 VGND
port 614 nsew ground input
rlabel locali s 298660 296463 298816 296497 6 VGND
port 614 nsew ground input
rlabel locali s 298660 296497 298799 296647 6 VGND
port 614 nsew ground input
rlabel locali s 1121 296313 1340 296463 6 VGND
port 614 nsew ground input
rlabel locali s 1104 296463 1340 296497 6 VGND
port 614 nsew ground input
rlabel locali s 1121 296497 1340 296647 6 VGND
port 614 nsew ground input
rlabel locali s 298695 296647 298799 296755 6 VGND
port 614 nsew ground input
rlabel locali s 1121 296647 1225 296755 6 VGND
port 614 nsew ground input
rlabel locali s 298695 297293 298799 297401 6 VGND
port 614 nsew ground input
rlabel locali s 1121 297293 1225 297401 6 VGND
port 614 nsew ground input
rlabel locali s 298660 297401 298799 297551 6 VGND
port 614 nsew ground input
rlabel locali s 298660 297551 298816 297585 6 VGND
port 614 nsew ground input
rlabel locali s 1121 297401 1340 297551 6 VGND
port 614 nsew ground input
rlabel locali s 1104 297551 1340 297585 6 VGND
port 614 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 300000 300000
string LEFview TRUE
<< end >>
